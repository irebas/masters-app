<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Warmińsko-Mazurski Okręgowy Związek Pływacki" version="11.73385">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Olsztyn" name="Letnie Mistrzostwa Polski w pływaniu w kategoriach masters" course="LCM" deadline="2022-05-27" reservecount="2" startmethod="1" timing="AUTOMATIC" type="WMC" nation="POL">
      <AGEDATE value="2022-12-31" type="YEAR" />
      <POOL name="Aquasfera" lanemax="9" />
      <FACILITY city="Olsztyn" name="Aquasfera" nation="POL" />
      <POINTTABLE pointtableid="997" name="MASTERS FINA WR" version="2022" />
      <FEES>
        <FEE type="ATHLETE" value="100" />
      </FEES>
      <QUALIFY from="2020-05-01" until="2022-06-05" />
      <SESSIONS>
        <SESSION date="2022-06-10" daytime="14:00" endtime="20:36" name="PIĄTEK" number="1">
          <EVENTS>
            <EVENT eventid="1059" daytime="14:00" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1060" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3296" />
                    <RANKING order="2" place="2" resultid="4194" />
                    <RANKING order="3" place="3" resultid="3164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1061" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2520" />
                    <RANKING order="2" place="2" resultid="3260" />
                    <RANKING order="3" place="3" resultid="3393" />
                    <RANKING order="4" place="4" resultid="2127" />
                    <RANKING order="5" place="5" resultid="2288" />
                    <RANKING order="6" place="6" resultid="2790" />
                    <RANKING order="7" place="7" resultid="3488" />
                    <RANKING order="8" place="8" resultid="3402" />
                    <RANKING order="9" place="9" resultid="3154" />
                    <RANKING order="10" place="-1" resultid="2972" />
                    <RANKING order="11" place="-1" resultid="2617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3268" />
                    <RANKING order="2" place="2" resultid="3264" />
                    <RANKING order="3" place="3" resultid="2644" />
                    <RANKING order="4" place="4" resultid="4262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3497" />
                    <RANKING order="2" place="2" resultid="2544" />
                    <RANKING order="3" place="3" resultid="3287" />
                    <RANKING order="4" place="4" resultid="3742" />
                    <RANKING order="5" place="5" resultid="3110" />
                    <RANKING order="6" place="6" resultid="3848" />
                    <RANKING order="7" place="7" resultid="1940" />
                    <RANKING order="8" place="8" resultid="2065" />
                    <RANKING order="9" place="9" resultid="2825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3451" />
                    <RANKING order="2" place="2" resultid="3122" />
                    <RANKING order="3" place="3" resultid="2056" />
                    <RANKING order="4" place="4" resultid="2490" />
                    <RANKING order="5" place="5" resultid="2072" />
                    <RANKING order="6" place="6" resultid="2988" />
                    <RANKING order="7" place="7" resultid="1809" />
                    <RANKING order="8" place="8" resultid="2535" />
                    <RANKING order="9" place="9" resultid="2311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3675" />
                    <RANKING order="2" place="2" resultid="1826" />
                    <RANKING order="3" place="3" resultid="2204" />
                    <RANKING order="4" place="4" resultid="2297" />
                    <RANKING order="5" place="5" resultid="2321" />
                    <RANKING order="6" place="6" resultid="2333" />
                    <RANKING order="7" place="7" resultid="3762" />
                    <RANKING order="8" place="-1" resultid="2338" />
                    <RANKING order="9" place="-1" resultid="2761" />
                    <RANKING order="10" place="-1" resultid="3071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2327" />
                    <RANKING order="2" place="2" resultid="2316" />
                    <RANKING order="3" place="3" resultid="3838" />
                    <RANKING order="4" place="4" resultid="3811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2049" />
                    <RANKING order="2" place="2" resultid="2737" />
                    <RANKING order="3" place="3" resultid="1817" />
                    <RANKING order="4" place="-1" resultid="3324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3242" />
                    <RANKING order="2" place="2" resultid="2864" />
                    <RANKING order="3" place="3" resultid="2996" />
                    <RANKING order="4" place="4" resultid="3239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4074" />
                    <RANKING order="2" place="2" resultid="3689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1072" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1073" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1074" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4266" daytime="14:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4267" daytime="14:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4268" daytime="14:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4269" daytime="14:09" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4270" daytime="14:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4271" daytime="14:14" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4272" daytime="14:16" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="14:18" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1078" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2622" />
                    <RANKING order="2" place="2" resultid="4119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4141" />
                    <RANKING order="2" place="2" resultid="3484" />
                    <RANKING order="3" place="3" resultid="2216" />
                    <RANKING order="4" place="4" resultid="3410" />
                    <RANKING order="5" place="5" resultid="2272" />
                    <RANKING order="6" place="6" resultid="2835" />
                    <RANKING order="7" place="7" resultid="3563" />
                    <RANKING order="8" place="8" resultid="2840" />
                    <RANKING order="9" place="9" resultid="3384" />
                    <RANKING order="10" place="10" resultid="3250" />
                    <RANKING order="11" place="11" resultid="2939" />
                    <RANKING order="12" place="12" resultid="3590" />
                    <RANKING order="13" place="-1" resultid="3367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3180" />
                    <RANKING order="2" place="2" resultid="4182" />
                    <RANKING order="3" place="3" resultid="3987" />
                    <RANKING order="4" place="4" resultid="3159" />
                    <RANKING order="5" place="5" resultid="2772" />
                    <RANKING order="6" place="6" resultid="3966" />
                    <RANKING order="7" place="7" resultid="3778" />
                    <RANKING order="8" place="8" resultid="2236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2795" />
                    <RANKING order="2" place="2" resultid="2225" />
                    <RANKING order="3" place="3" resultid="3899" />
                    <RANKING order="4" place="4" resultid="3134" />
                    <RANKING order="5" place="5" resultid="3842" />
                    <RANKING order="6" place="6" resultid="3204" />
                    <RANKING order="7" place="7" resultid="4145" />
                    <RANKING order="8" place="8" resultid="2932" />
                    <RANKING order="9" place="9" resultid="3196" />
                    <RANKING order="10" place="10" resultid="2394" />
                    <RANKING order="11" place="11" resultid="2356" />
                    <RANKING order="12" place="-1" resultid="2245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3029" />
                    <RANKING order="2" place="2" resultid="2781" />
                    <RANKING order="3" place="3" resultid="2732" />
                    <RANKING order="4" place="4" resultid="4173" />
                    <RANKING order="5" place="5" resultid="4159" />
                    <RANKING order="6" place="6" resultid="2727" />
                    <RANKING order="7" place="7" resultid="2495" />
                    <RANKING order="8" place="8" resultid="2347" />
                    <RANKING order="9" place="9" resultid="3127" />
                    <RANKING order="10" place="10" resultid="1861" />
                    <RANKING order="11" place="11" resultid="2960" />
                    <RANKING order="12" place="12" resultid="2955" />
                    <RANKING order="13" place="13" resultid="4501" />
                    <RANKING order="14" place="14" resultid="4166" />
                    <RANKING order="15" place="15" resultid="4203" />
                    <RANKING order="16" place="16" resultid="2502" />
                    <RANKING order="17" place="17" resultid="3765" />
                    <RANKING order="18" place="18" resultid="2602" />
                    <RANKING order="19" place="19" resultid="3623" />
                    <RANKING order="20" place="20" resultid="2398" />
                    <RANKING order="21" place="21" resultid="3825" />
                    <RANKING order="22" place="22" resultid="3586" />
                    <RANKING order="23" place="23" resultid="3929" />
                    <RANKING order="24" place="-1" resultid="3140" />
                    <RANKING order="25" place="-1" resultid="3704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1845" />
                    <RANKING order="2" place="2" resultid="3001" />
                    <RANKING order="3" place="3" resultid="3347" />
                    <RANKING order="4" place="4" resultid="3216" />
                    <RANKING order="5" place="5" resultid="3515" />
                    <RANKING order="6" place="6" resultid="4229" />
                    <RANKING order="7" place="7" resultid="2220" />
                    <RANKING order="8" place="8" resultid="4151" />
                    <RANKING order="9" place="9" resultid="3333" />
                    <RANKING order="10" place="10" resultid="2650" />
                    <RANKING order="11" place="11" resultid="3506" />
                    <RANKING order="12" place="12" resultid="2387" />
                    <RANKING order="13" place="13" resultid="3478" />
                    <RANKING order="14" place="14" resultid="2498" />
                    <RANKING order="15" place="15" resultid="1853" />
                    <RANKING order="16" place="16" resultid="1838" />
                    <RANKING order="17" place="-1" resultid="3621" />
                    <RANKING order="18" place="-1" resultid="2926" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2095" />
                    <RANKING order="2" place="2" resultid="4211" />
                    <RANKING order="3" place="3" resultid="3095" />
                    <RANKING order="4" place="4" resultid="2209" />
                    <RANKING order="5" place="5" resultid="4041" />
                    <RANKING order="6" place="6" resultid="3904" />
                    <RANKING order="7" place="7" resultid="2891" />
                    <RANKING order="8" place="8" resultid="4196" />
                    <RANKING order="9" place="9" resultid="2251" />
                    <RANKING order="10" place="-1" resultid="1831" />
                    <RANKING order="11" place="-1" resultid="3719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2745" />
                    <RANKING order="2" place="2" resultid="2912" />
                    <RANKING order="3" place="3" resultid="2665" />
                    <RANKING order="4" place="4" resultid="4126" />
                    <RANKING order="5" place="5" resultid="3210" />
                    <RANKING order="6" place="6" resultid="3656" />
                    <RANKING order="7" place="7" resultid="3076" />
                    <RANKING order="8" place="8" resultid="2803" />
                    <RANKING order="9" place="9" resultid="3169" />
                    <RANKING order="10" place="10" resultid="3805" />
                    <RANKING order="11" place="11" resultid="1949" />
                    <RANKING order="12" place="-1" resultid="3772" />
                    <RANKING order="13" place="-1" resultid="3952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2903" />
                    <RANKING order="2" place="2" resultid="2086" />
                    <RANKING order="3" place="3" resultid="3306" />
                    <RANKING order="4" place="4" resultid="2820" />
                    <RANKING order="5" place="5" resultid="3978" />
                    <RANKING order="6" place="6" resultid="2380" />
                    <RANKING order="7" place="7" resultid="3636" />
                    <RANKING order="8" place="8" resultid="2656" />
                    <RANKING order="9" place="9" resultid="2030" />
                    <RANKING order="10" place="-1" resultid="2343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2921" />
                    <RANKING order="2" place="2" resultid="3752" />
                    <RANKING order="3" place="3" resultid="2371" />
                    <RANKING order="4" place="4" resultid="3759" />
                    <RANKING order="5" place="5" resultid="2480" />
                    <RANKING order="6" place="6" resultid="3008" />
                    <RANKING order="7" place="-1" resultid="2079" />
                    <RANKING order="8" place="-1" resultid="4253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3547" />
                    <RANKING order="2" place="1" resultid="4057" />
                    <RANKING order="3" place="3" resultid="2364" />
                    <RANKING order="4" place="4" resultid="3227" />
                    <RANKING order="5" place="5" resultid="3470" />
                    <RANKING order="6" place="6" resultid="3831" />
                    <RANKING order="7" place="7" resultid="4084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3641" />
                    <RANKING order="2" place="2" resultid="3084" />
                    <RANKING order="3" place="3" resultid="3724" />
                    <RANKING order="4" place="4" resultid="3574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4061" />
                    <RANKING order="2" place="2" resultid="3231" />
                    <RANKING order="3" place="3" resultid="3062" />
                    <RANKING order="4" place="4" resultid="3697" />
                    <RANKING order="5" place="-1" resultid="3568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1092" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4273" daytime="14:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4274" daytime="14:21" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4275" daytime="14:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4276" daytime="14:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4277" daytime="14:29" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4278" daytime="14:31" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4279" daytime="14:33" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4280" daytime="14:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4281" daytime="14:37" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4282" daytime="14:39" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4283" daytime="14:41" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4284" daytime="14:43" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4285" daytime="14:45" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4286" daytime="14:47" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1094" daytime="14:49" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1096" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2463" />
                    <RANKING order="2" place="2" resultid="3924" />
                    <RANKING order="3" place="3" resultid="3853" />
                    <RANKING order="4" place="4" resultid="3933" />
                    <RANKING order="5" place="-1" resultid="3297" />
                    <RANKING order="6" place="-1" resultid="2632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3394" />
                    <RANKING order="2" place="2" resultid="4103" />
                    <RANKING order="3" place="3" resultid="2404" />
                    <RANKING order="4" place="4" resultid="3489" />
                    <RANKING order="5" place="-1" resultid="2627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3498" />
                    <RANKING order="2" place="2" resultid="3288" />
                    <RANKING order="3" place="3" resultid="3743" />
                    <RANKING order="4" place="4" resultid="2545" />
                    <RANKING order="5" place="5" resultid="2039" />
                    <RANKING order="6" place="6" resultid="1941" />
                    <RANKING order="7" place="-1" resultid="3111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3452" />
                    <RANKING order="2" place="2" resultid="2057" />
                    <RANKING order="3" place="3" resultid="2073" />
                    <RANKING order="4" place="4" resultid="4220" />
                    <RANKING order="5" place="5" resultid="2989" />
                    <RANKING order="6" place="6" resultid="4001" />
                    <RANKING order="7" place="-1" resultid="2536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4010" />
                    <RANKING order="2" place="2" resultid="2869" />
                    <RANKING order="3" place="3" resultid="2409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2328" />
                    <RANKING order="2" place="2" resultid="1957" />
                    <RANKING order="3" place="3" resultid="3532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3325" />
                    <RANKING order="2" place="2" resultid="3184" />
                    <RANKING order="3" place="3" resultid="3612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2100" />
                    <RANKING order="2" place="2" resultid="2109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1107" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1108" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1109" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1110" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1111" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4287" daytime="14:49" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4288" daytime="14:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4289" daytime="15:01" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4290" daytime="15:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1112" daytime="15:11" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1113" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2722" />
                    <RANKING order="2" place="2" resultid="3433" />
                    <RANKING order="3" place="3" resultid="3940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2718" />
                    <RANKING order="2" place="2" resultid="1870" />
                    <RANKING order="3" place="3" resultid="3039" />
                    <RANKING order="4" place="4" resultid="3418" />
                    <RANKING order="5" place="5" resultid="3411" />
                    <RANKING order="6" place="-1" resultid="3251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3596" />
                    <RANKING order="2" place="2" resultid="3988" />
                    <RANKING order="3" place="3" resultid="4121" />
                    <RANKING order="4" place="-1" resultid="3791" />
                    <RANKING order="5" place="-1" resultid="3376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2933" />
                    <RANKING order="2" place="2" resultid="3524" />
                    <RANKING order="3" place="3" resultid="3135" />
                    <RANKING order="4" place="-1" resultid="3909" />
                    <RANKING order="5" place="-1" resultid="1892" />
                    <RANKING order="6" place="-1" resultid="2246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2782" />
                    <RANKING order="2" place="2" resultid="3277" />
                    <RANKING order="3" place="3" resultid="4174" />
                    <RANKING order="4" place="4" resultid="4160" />
                    <RANKING order="5" place="5" resultid="2676" />
                    <RANKING order="6" place="6" resultid="3540" />
                    <RANKING order="7" place="-1" resultid="1879" />
                    <RANKING order="8" place="-1" resultid="2348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3348" />
                    <RANKING order="2" place="2" resultid="3516" />
                    <RANKING order="3" place="3" resultid="4230" />
                    <RANKING order="4" place="4" resultid="2670" />
                    <RANKING order="5" place="5" resultid="2965" />
                    <RANKING order="6" place="6" resultid="3315" />
                    <RANKING order="7" place="-1" resultid="3782" />
                    <RANKING order="8" place="-1" resultid="2388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3089" />
                    <RANKING order="2" place="2" resultid="2607" />
                    <RANKING order="3" place="3" resultid="3905" />
                    <RANKING order="4" place="4" resultid="4197" />
                    <RANKING order="5" place="5" resultid="2858" />
                    <RANKING order="6" place="6" resultid="2892" />
                    <RANKING order="7" place="7" resultid="3973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2913" />
                    <RANKING order="2" place="2" resultid="3657" />
                    <RANKING order="3" place="3" resultid="3773" />
                    <RANKING order="4" place="4" resultid="2948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2904" />
                    <RANKING order="2" place="2" resultid="3307" />
                    <RANKING order="3" place="3" resultid="1886" />
                    <RANKING order="4" place="4" resultid="3881" />
                    <RANKING order="5" place="5" resultid="3980" />
                    <RANKING order="6" place="6" resultid="3637" />
                    <RANKING order="7" place="-1" resultid="2087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2700" />
                    <RANKING order="2" place="2" resultid="2372" />
                    <RANKING order="3" place="3" resultid="3888" />
                    <RANKING order="4" place="4" resultid="2879" />
                    <RANKING order="5" place="5" resultid="3680" />
                    <RANKING order="6" place="-1" resultid="2830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3914" />
                    <RANKING order="2" place="2" resultid="3013" />
                    <RANKING order="3" place="3" resultid="3339" />
                    <RANKING order="4" place="4" resultid="2365" />
                    <RANKING order="5" place="5" resultid="3460" />
                    <RANKING order="6" place="6" resultid="3832" />
                    <RANKING order="7" place="7" resultid="3955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1127" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1128" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4291" daytime="15:11" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4292" daytime="15:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4293" daytime="15:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4294" daytime="15:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4295" daytime="15:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4296" daytime="15:39" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4297" daytime="15:44" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1129" daytime="15:48" gender="X" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1145" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="1765" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1766" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3049" />
                    <RANKING order="2" place="2" resultid="5038" />
                    <RANKING order="3" place="3" resultid="1917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1767" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3144" />
                    <RANKING order="2" place="2" resultid="1918" />
                    <RANKING order="3" place="3" resultid="3190" />
                    <RANKING order="4" place="4" resultid="2445" />
                    <RANKING order="5" place="5" resultid="1979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1768" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2121" />
                    <RANKING order="2" place="2" resultid="2446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1769" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2447" />
                    <RANKING order="2" place="2" resultid="2900" />
                    <RANKING order="3" place="3" resultid="3583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1771" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4088" />
                    <RANKING order="2" place="2" resultid="3246" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4488" daytime="15:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4489" daytime="15:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1146" daytime="15:56" gender="F" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1147" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2464" />
                    <RANKING order="2" place="2" resultid="3165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4104" />
                    <RANKING order="2" place="2" resultid="2638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1149" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1150" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3651" />
                    <RANKING order="2" place="2" resultid="4221" />
                    <RANKING order="3" place="-1" resultid="3816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2258" />
                    <RANKING order="2" place="2" resultid="3629" />
                    <RANKING order="3" place="3" resultid="2410" />
                    <RANKING order="4" place="4" resultid="5039" />
                    <RANKING order="5" place="-1" resultid="2762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1958" />
                    <RANKING order="2" place="2" resultid="3533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4091" />
                    <RANKING order="2" place="2" resultid="4133" />
                    <RANKING order="3" place="3" resultid="3185" />
                    <RANKING order="4" place="4" resultid="4021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2710" />
                    <RANKING order="2" place="-1" resultid="3555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1158" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1160" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1161" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1162" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4300" daytime="15:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4301" daytime="16:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4302" daytime="16:30" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1163" daytime="16:52" gender="M" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1164" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1165" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2273" />
                    <RANKING order="2" place="2" resultid="3368" />
                    <RANKING order="3" place="3" resultid="3591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3989" />
                    <RANKING order="2" place="2" resultid="3779" />
                    <RANKING order="3" place="3" resultid="3377" />
                    <RANKING order="4" place="4" resultid="3968" />
                    <RANKING order="5" place="-1" resultid="3711" />
                    <RANKING order="6" place="-1" resultid="3792" />
                    <RANKING order="7" place="-1" resultid="2237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3900" />
                    <RANKING order="2" place="2" resultid="2226" />
                    <RANKING order="3" place="3" resultid="3525" />
                    <RANKING order="4" place="4" resultid="3867" />
                    <RANKING order="5" place="5" resultid="3175" />
                    <RANKING order="6" place="6" resultid="3582" />
                    <RANKING order="7" place="-1" resultid="3843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3278" />
                    <RANKING order="2" place="2" resultid="4167" />
                    <RANKING order="3" place="3" resultid="4204" />
                    <RANKING order="4" place="4" resultid="2603" />
                    <RANKING order="5" place="5" resultid="3541" />
                    <RANKING order="6" place="-1" resultid="1880" />
                    <RANKING order="7" place="-1" resultid="3705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1846" />
                    <RANKING order="2" place="2" resultid="3893" />
                    <RANKING order="3" place="3" resultid="1900" />
                    <RANKING order="4" place="4" resultid="3316" />
                    <RANKING order="5" place="5" resultid="3507" />
                    <RANKING order="6" place="6" resultid="2263" />
                    <RANKING order="7" place="7" resultid="3783" />
                    <RANKING order="8" place="8" resultid="2424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4212" />
                    <RANKING order="2" place="2" resultid="2210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4127" />
                    <RANKING order="2" place="2" resultid="2804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1887" />
                    <RANKING order="2" place="2" resultid="2657" />
                    <RANKING order="3" place="3" resultid="2031" />
                    <RANKING order="4" place="-1" resultid="2753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2880" />
                    <RANKING order="2" place="2" resultid="2481" />
                    <RANKING order="3" place="-1" resultid="4254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3548" />
                    <RANKING order="2" place="2" resultid="2418" />
                    <RANKING order="3" place="3" resultid="3461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1176" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1178" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4303" daytime="16:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4304" daytime="17:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4305" daytime="17:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4306" daytime="17:31" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4307" daytime="17:59" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1180" daytime="18:26" gender="F" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1181" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3934" />
                    <RANKING order="2" place="2" resultid="4099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="1183" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1184" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1185" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1186" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="1188" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3872" />
                    <RANKING order="2" place="2" resultid="3613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1191" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1193" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1194" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1195" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1196" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4308" daytime="18:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1197" daytime="19:06" gender="M" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1198" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2776" />
                    <RANKING order="2" place="2" resultid="1871" />
                    <RANKING order="3" place="3" resultid="3385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1862" />
                    <RANKING order="2" place="2" resultid="3717" />
                    <RANKING order="3" place="3" resultid="1908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4152" />
                    <RANKING order="2" place="2" resultid="3665" />
                    <RANKING order="3" place="3" resultid="2966" />
                    <RANKING order="4" place="4" resultid="4101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2859" />
                    <RANKING order="2" place="2" resultid="2608" />
                    <RANKING order="3" place="3" resultid="4042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3669" />
                    <RANKING order="2" place="-1" resultid="2344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3753" />
                    <RANKING order="2" place="2" resultid="3681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2873" />
                    <RANKING order="2" place="2" resultid="3471" />
                    <RANKING order="3" place="-1" resultid="3915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1211" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1212" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1213" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4309" daytime="19:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4310" daytime="19:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4311" daytime="20:01" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2022-06-11" daytime="09:00" endtime="16:18" name="SOBOTA" number="2">
          <EVENTS>
            <EVENT eventid="1215" daytime="09:00" gender="F" number="10" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1217" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2633" />
                    <RANKING order="2" place="2" resultid="3298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2521" />
                    <RANKING order="2" place="2" resultid="2973" />
                    <RANKING order="3" place="3" resultid="3395" />
                    <RANKING order="4" place="4" resultid="2472" />
                    <RANKING order="5" place="5" resultid="3272" />
                    <RANKING order="6" place="6" resultid="2618" />
                    <RANKING order="7" place="7" resultid="3403" />
                    <RANKING order="8" place="8" resultid="3155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3265" />
                    <RANKING order="2" place="2" resultid="2977" />
                    <RANKING order="3" place="3" resultid="4263" />
                    <RANKING order="4" place="4" resultid="2645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3289" />
                    <RANKING order="2" place="2" resultid="3499" />
                    <RANKING order="3" place="3" resultid="2546" />
                    <RANKING order="4" place="4" resultid="3744" />
                    <RANKING order="5" place="5" resultid="3112" />
                    <RANKING order="6" place="6" resultid="2066" />
                    <RANKING order="7" place="7" resultid="1942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2506" />
                    <RANKING order="2" place="2" resultid="2058" />
                    <RANKING order="3" place="3" resultid="3453" />
                    <RANKING order="4" place="4" resultid="4002" />
                    <RANKING order="5" place="5" resultid="1810" />
                    <RANKING order="6" place="6" resultid="2537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1827" />
                    <RANKING order="2" place="2" resultid="2259" />
                    <RANKING order="3" place="3" resultid="2812" />
                    <RANKING order="4" place="4" resultid="3677" />
                    <RANKING order="5" place="5" resultid="3763" />
                    <RANKING order="6" place="6" resultid="3630" />
                    <RANKING order="7" place="-1" resultid="2339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2329" />
                    <RANKING order="2" place="2" resultid="2317" />
                    <RANKING order="3" place="3" resultid="3534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2050" />
                    <RANKING order="2" place="2" resultid="2738" />
                    <RANKING order="3" place="3" resultid="4134" />
                    <RANKING order="4" place="4" resultid="3614" />
                    <RANKING order="5" place="5" resultid="3081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2305" />
                    <RANKING order="2" place="2" resultid="2111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2711" />
                    <RANKING order="2" place="2" resultid="3556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2865" />
                    <RANKING order="2" place="2" resultid="3240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4075" />
                    <RANKING order="2" place="2" resultid="3690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1230" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1231" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1232" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4312" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4313" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4314" daytime="09:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4315" daytime="09:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4316" daytime="09:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1267" daytime="09:11" gender="M" number="11" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1268" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3731" />
                    <RANKING order="2" place="-1" resultid="3941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3862" />
                    <RANKING order="2" place="2" resultid="3412" />
                    <RANKING order="3" place="3" resultid="3369" />
                    <RANKING order="4" place="4" resultid="3386" />
                    <RANKING order="5" place="-1" resultid="2836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1270" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4183" />
                    <RANKING order="2" place="2" resultid="3378" />
                    <RANKING order="3" place="3" resultid="2118" />
                    <RANKING order="4" place="4" resultid="3962" />
                    <RANKING order="5" place="5" resultid="2238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4242" />
                    <RANKING order="2" place="2" resultid="2357" />
                    <RANKING order="3" place="-1" resultid="2247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3030" />
                    <RANKING order="2" place="2" resultid="2783" />
                    <RANKING order="3" place="3" resultid="4175" />
                    <RANKING order="4" place="4" resultid="2728" />
                    <RANKING order="5" place="5" resultid="1863" />
                    <RANKING order="6" place="6" resultid="2677" />
                    <RANKING order="7" place="7" resultid="2956" />
                    <RANKING order="8" place="8" resultid="2399" />
                    <RANKING order="9" place="9" resultid="3624" />
                    <RANKING order="10" place="-1" resultid="2944" />
                    <RANKING order="11" place="-1" resultid="3105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3334" />
                    <RANKING order="2" place="2" resultid="2221" />
                    <RANKING order="3" place="3" resultid="4153" />
                    <RANKING order="4" place="4" resultid="3317" />
                    <RANKING order="5" place="5" resultid="4231" />
                    <RANKING order="6" place="6" resultid="1901" />
                    <RANKING order="7" place="7" resultid="2264" />
                    <RANKING order="8" place="8" resultid="3508" />
                    <RANKING order="9" place="9" resultid="3479" />
                    <RANKING order="10" place="10" resultid="3784" />
                    <RANKING order="11" place="11" resultid="2389" />
                    <RANKING order="12" place="12" resultid="1855" />
                    <RANKING order="13" place="-1" resultid="2927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3096" />
                    <RANKING order="2" place="2" resultid="4213" />
                    <RANKING order="3" place="3" resultid="4043" />
                    <RANKING order="4" place="4" resultid="2609" />
                    <RANKING order="5" place="5" resultid="2893" />
                    <RANKING order="6" place="6" resultid="2278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2914" />
                    <RANKING order="2" place="2" resultid="2746" />
                    <RANKING order="3" place="3" resultid="4128" />
                    <RANKING order="4" place="4" resultid="3359" />
                    <RANKING order="5" place="5" resultid="3806" />
                    <RANKING order="6" place="6" resultid="1966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3099" />
                    <RANKING order="2" place="2" resultid="2088" />
                    <RANKING order="3" place="3" resultid="2754" />
                    <RANKING order="4" place="4" resultid="2905" />
                    <RANKING order="5" place="5" resultid="2658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3760" />
                    <RANKING order="2" place="2" resultid="2373" />
                    <RANKING order="3" place="3" resultid="3683" />
                    <RANKING order="4" place="4" resultid="2482" />
                    <RANKING order="5" place="5" resultid="2881" />
                    <RANKING order="6" place="6" resultid="3009" />
                    <RANKING order="7" place="7" resultid="2080" />
                    <RANKING order="8" place="-1" resultid="4255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3916" />
                    <RANKING order="2" place="2" resultid="2874" />
                    <RANKING order="3" place="3" resultid="3340" />
                    <RANKING order="4" place="4" resultid="3462" />
                    <RANKING order="5" place="5" resultid="2431" />
                    <RANKING order="6" place="6" resultid="4085" />
                    <RANKING order="7" place="7" resultid="3833" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4052" />
                    <RANKING order="2" place="2" resultid="3085" />
                    <RANKING order="3" place="3" resultid="3575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3233" />
                    <RANKING order="2" place="2" resultid="3064" />
                    <RANKING order="3" place="3" resultid="3698" />
                    <RANKING order="4" place="-1" resultid="3569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1282" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1283" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4318" daytime="09:11" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4319" daytime="09:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4320" daytime="09:17" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4321" daytime="09:19" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4322" daytime="09:21" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4323" daytime="09:23" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4324" daytime="09:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4325" daytime="09:27" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1233" daytime="09:28" gender="F" number="12" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1234" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2465" />
                    <RANKING order="2" place="2" resultid="3925" />
                    <RANKING order="3" place="3" resultid="3855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2791" />
                    <RANKING order="2" place="2" resultid="2405" />
                    <RANKING order="3" place="3" resultid="3490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2978" />
                    <RANKING order="2" place="2" resultid="3046" />
                    <RANKING order="3" place="3" resultid="4016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2547" />
                    <RANKING order="2" place="2" resultid="2067" />
                    <RANKING order="3" place="-1" resultid="2826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4222" />
                    <RANKING order="2" place="2" resultid="3817" />
                    <RANKING order="3" place="3" resultid="2312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2870" />
                    <RANKING order="2" place="2" resultid="2298" />
                    <RANKING order="3" place="3" resultid="2411" />
                    <RANKING order="4" place="4" resultid="5040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3326" />
                    <RANKING order="2" place="2" resultid="1819" />
                    <RANKING order="3" place="3" resultid="3186" />
                    <RANKING order="4" place="-1" resultid="3019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1243" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1244" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2527" />
                    <RANKING order="2" place="2" resultid="4080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1247" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1249" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4326" daytime="09:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4327" daytime="09:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4328" daytime="09:44" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1250" daytime="09:48" gender="M" number="13" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1251" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3435" />
                    <RANKING order="2" place="-1" resultid="3942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2777" />
                    <RANKING order="2" place="2" resultid="3419" />
                    <RANKING order="3" place="3" resultid="3252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4122" />
                    <RANKING order="2" place="2" resultid="3713" />
                    <RANKING order="3" place="3" resultid="3597" />
                    <RANKING order="4" place="4" resultid="3963" />
                    <RANKING order="5" place="5" resultid="3793" />
                    <RANKING order="6" place="-1" resultid="2508" />
                    <RANKING order="7" place="-1" resultid="2850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2934" />
                    <RANKING order="2" place="2" resultid="3526" />
                    <RANKING order="3" place="3" resultid="3136" />
                    <RANKING order="4" place="4" resultid="2984" />
                    <RANKING order="5" place="5" resultid="1893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4161" />
                    <RANKING order="2" place="2" resultid="3279" />
                    <RANKING order="3" place="3" resultid="3443" />
                    <RANKING order="4" place="4" resultid="4205" />
                    <RANKING order="5" place="5" resultid="1910" />
                    <RANKING order="6" place="-1" resultid="1881" />
                    <RANKING order="7" place="-1" resultid="2349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2967" />
                    <RANKING order="2" place="2" resultid="3318" />
                    <RANKING order="3" place="3" resultid="1839" />
                    <RANKING order="4" place="4" resultid="2425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2292" />
                    <RANKING order="2" place="2" resultid="4198" />
                    <RANKING order="3" place="3" resultid="3707" />
                    <RANKING order="4" place="4" resultid="1832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2805" />
                    <RANKING order="2" place="2" resultid="2666" />
                    <RANKING order="3" place="3" resultid="2887" />
                    <RANKING order="4" place="4" resultid="1973" />
                    <RANKING order="5" place="-1" resultid="1950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2821" />
                    <RANKING order="2" place="2" resultid="2089" />
                    <RANKING order="3" place="3" resultid="1888" />
                    <RANKING order="4" place="4" resultid="2381" />
                    <RANKING order="5" place="5" resultid="3981" />
                    <RANKING order="6" place="6" resultid="2436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4094" />
                    <RANKING order="2" place="2" resultid="2701" />
                    <RANKING order="3" place="3" resultid="2374" />
                    <RANKING order="4" place="4" resultid="3889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3014" />
                    <RANKING order="2" place="2" resultid="3917" />
                    <RANKING order="3" place="3" resultid="2419" />
                    <RANKING order="4" place="4" resultid="3341" />
                    <RANKING order="5" place="5" resultid="3956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3643" />
                    <RANKING order="2" place="2" resultid="3576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4062" />
                    <RANKING order="2" place="2" resultid="3234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1265" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4329" daytime="09:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4330" daytime="09:57" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4331" daytime="10:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4332" daytime="10:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4333" daytime="10:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4334" daytime="10:20" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1284" daytime="10:24" gender="F" number="14" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1285" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3299" />
                    <RANKING order="2" place="2" resultid="3166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3261" />
                    <RANKING order="2" place="2" resultid="2128" />
                    <RANKING order="3" place="3" resultid="3396" />
                    <RANKING order="4" place="4" resultid="2289" />
                    <RANKING order="5" place="5" resultid="3491" />
                    <RANKING order="6" place="6" resultid="2619" />
                    <RANKING order="7" place="7" resultid="2628" />
                    <RANKING order="8" place="8" resultid="3156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3269" />
                    <RANKING order="2" place="2" resultid="3047" />
                    <RANKING order="3" place="3" resultid="2646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3500" />
                    <RANKING order="2" place="2" resultid="3290" />
                    <RANKING order="3" place="3" resultid="3113" />
                    <RANKING order="4" place="4" resultid="3849" />
                    <RANKING order="5" place="5" resultid="2041" />
                    <RANKING order="6" place="6" resultid="1943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3652" />
                    <RANKING order="2" place="2" resultid="3454" />
                    <RANKING order="3" place="3" resultid="3123" />
                    <RANKING order="4" place="4" resultid="2059" />
                    <RANKING order="5" place="5" resultid="2990" />
                    <RANKING order="6" place="6" resultid="2074" />
                    <RANKING order="7" place="7" resultid="4223" />
                    <RANKING order="8" place="8" resultid="3818" />
                    <RANKING order="9" place="9" resultid="3800" />
                    <RANKING order="10" place="10" resultid="1811" />
                    <RANKING order="11" place="11" resultid="2440" />
                    <RANKING order="12" place="12" resultid="2538" />
                    <RANKING order="13" place="-1" resultid="2491" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4006" />
                    <RANKING order="2" place="2" resultid="2205" />
                    <RANKING order="3" place="3" resultid="1828" />
                    <RANKING order="4" place="4" resultid="3631" />
                    <RANKING order="5" place="5" resultid="2322" />
                    <RANKING order="6" place="6" resultid="2334" />
                    <RANKING order="7" place="-1" resultid="3072" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2318" />
                    <RANKING order="2" place="2" resultid="1960" />
                    <RANKING order="3" place="3" resultid="3839" />
                    <RANKING order="4" place="4" resultid="3535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3873" />
                    <RANKING order="2" place="2" resultid="2051" />
                    <RANKING order="3" place="3" resultid="2739" />
                    <RANKING order="4" place="4" resultid="1820" />
                    <RANKING order="5" place="5" resultid="4135" />
                    <RANKING order="6" place="6" resultid="3615" />
                    <RANKING order="7" place="-1" resultid="3327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2306" />
                    <RANKING order="2" place="2" resultid="2102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2712" />
                    <RANKING order="2" place="2" resultid="3557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2866" />
                    <RANKING order="2" place="2" resultid="2528" />
                    <RANKING order="3" place="3" resultid="2998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4076" />
                    <RANKING order="2" place="2" resultid="3691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1298" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1299" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1300" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4335" daytime="10:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4336" daytime="10:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4337" daytime="10:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4338" daytime="10:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4339" daytime="10:39" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4340" daytime="10:41" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1301" daytime="10:43" gender="M" number="15" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1302" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2723" />
                    <RANKING order="2" place="2" resultid="3732" />
                    <RANKING order="3" place="-1" resultid="2623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1303" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4142" />
                    <RANKING order="2" place="2" resultid="2217" />
                    <RANKING order="3" place="3" resultid="3370" />
                    <RANKING order="4" place="4" resultid="1872" />
                    <RANKING order="5" place="5" resultid="3040" />
                    <RANKING order="6" place="6" resultid="4500" />
                    <RANKING order="7" place="7" resultid="3564" />
                    <RANKING order="8" place="8" resultid="3387" />
                    <RANKING order="9" place="9" resultid="3592" />
                    <RANKING order="10" place="10" resultid="2940" />
                    <RANKING order="11" place="11" resultid="3253" />
                    <RANKING order="12" place="-1" resultid="2837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3181" />
                    <RANKING order="2" place="2" resultid="3990" />
                    <RANKING order="3" place="3" resultid="2845" />
                    <RANKING order="4" place="4" resultid="4184" />
                    <RANKING order="5" place="5" resultid="3160" />
                    <RANKING order="6" place="6" resultid="2773" />
                    <RANKING order="7" place="7" resultid="3780" />
                    <RANKING order="8" place="8" resultid="2239" />
                    <RANKING order="9" place="9" resultid="3609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3603" />
                    <RANKING order="2" place="2" resultid="3118" />
                    <RANKING order="3" place="3" resultid="2797" />
                    <RANKING order="4" place="4" resultid="2227" />
                    <RANKING order="5" place="5" resultid="3901" />
                    <RANKING order="6" place="6" resultid="3024" />
                    <RANKING order="7" place="7" resultid="4146" />
                    <RANKING order="8" place="8" resultid="3844" />
                    <RANKING order="9" place="9" resultid="3205" />
                    <RANKING order="10" place="10" resultid="3176" />
                    <RANKING order="11" place="11" resultid="3197" />
                    <RANKING order="12" place="12" resultid="2395" />
                    <RANKING order="13" place="13" resultid="2358" />
                    <RANKING order="14" place="-1" resultid="2248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2784" />
                    <RANKING order="2" place="2" resultid="4176" />
                    <RANKING order="3" place="3" resultid="2496" />
                    <RANKING order="4" place="4" resultid="2733" />
                    <RANKING order="5" place="5" resultid="3128" />
                    <RANKING order="6" place="6" resultid="2350" />
                    <RANKING order="7" place="7" resultid="2961" />
                    <RANKING order="8" place="8" resultid="1864" />
                    <RANKING order="9" place="9" resultid="3447" />
                    <RANKING order="10" place="10" resultid="2503" />
                    <RANKING order="11" place="11" resultid="2604" />
                    <RANKING order="12" place="12" resultid="3625" />
                    <RANKING order="13" place="13" resultid="3826" />
                    <RANKING order="14" place="14" resultid="3930" />
                    <RANKING order="15" place="15" resultid="3587" />
                    <RANKING order="16" place="-1" resultid="3141" />
                    <RANKING order="17" place="-1" resultid="3201" />
                    <RANKING order="18" place="-1" resultid="3766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3349" />
                    <RANKING order="2" place="2" resultid="3002" />
                    <RANKING order="3" place="3" resultid="3517" />
                    <RANKING order="4" place="4" resultid="3217" />
                    <RANKING order="5" place="5" resultid="3894" />
                    <RANKING order="6" place="6" resultid="1902" />
                    <RANKING order="7" place="7" resultid="2651" />
                    <RANKING order="8" place="8" resultid="3480" />
                    <RANKING order="9" place="9" resultid="2390" />
                    <RANKING order="10" place="10" resultid="3785" />
                    <RANKING order="11" place="11" resultid="2499" />
                    <RANKING order="12" place="12" resultid="1840" />
                    <RANKING order="13" place="-1" resultid="1856" />
                    <RANKING order="14" place="-1" resultid="4232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3090" />
                    <RANKING order="2" place="2" resultid="2096" />
                    <RANKING order="3" place="3" resultid="4214" />
                    <RANKING order="4" place="4" resultid="2211" />
                    <RANKING order="5" place="5" resultid="3906" />
                    <RANKING order="6" place="6" resultid="2894" />
                    <RANKING order="7" place="7" resultid="1833" />
                    <RANKING order="8" place="8" resultid="3708" />
                    <RANKING order="9" place="-1" resultid="3720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2747" />
                    <RANKING order="2" place="2" resultid="2915" />
                    <RANKING order="3" place="3" resultid="3658" />
                    <RANKING order="4" place="4" resultid="3077" />
                    <RANKING order="5" place="5" resultid="3211" />
                    <RANKING order="6" place="6" resultid="3170" />
                    <RANKING order="7" place="7" resultid="3807" />
                    <RANKING order="8" place="8" resultid="1951" />
                    <RANKING order="9" place="9" resultid="4112" />
                    <RANKING order="10" place="10" resultid="1967" />
                    <RANKING order="11" place="-1" resultid="3774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2906" />
                    <RANKING order="2" place="2" resultid="2755" />
                    <RANKING order="3" place="3" resultid="3308" />
                    <RANKING order="4" place="4" resultid="2659" />
                    <RANKING order="5" place="5" resultid="3979" />
                    <RANKING order="6" place="6" resultid="3670" />
                    <RANKING order="7" place="7" resultid="2382" />
                    <RANKING order="8" place="8" resultid="2032" />
                    <RANKING order="9" place="-1" resultid="2345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2922" />
                    <RANKING order="2" place="2" resultid="3754" />
                    <RANKING order="3" place="3" resultid="2483" />
                    <RANKING order="4" place="4" resultid="3010" />
                    <RANKING order="5" place="5" resultid="2081" />
                    <RANKING order="6" place="-1" resultid="4256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3549" />
                    <RANKING order="2" place="2" resultid="2366" />
                    <RANKING order="3" place="3" resultid="4058" />
                    <RANKING order="4" place="4" resultid="3472" />
                    <RANKING order="5" place="5" resultid="3228" />
                    <RANKING order="6" place="-1" resultid="3834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3644" />
                    <RANKING order="2" place="2" resultid="3726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3065" />
                    <RANKING order="2" place="2" resultid="3699" />
                    <RANKING order="3" place="-1" resultid="3570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1316" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1317" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4341" daytime="10:43" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4342" daytime="10:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4343" daytime="10:49" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4344" daytime="10:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4345" daytime="10:57" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4346" daytime="10:59" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4347" daytime="11:01" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4348" daytime="11:04" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4349" daytime="11:06" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4350" daytime="11:08" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4351" daytime="11:10" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4352" daytime="11:12" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1335" daytime="11:14" gender="F" number="16" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1336" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2466" />
                    <RANKING order="2" place="2" resultid="2476" />
                    <RANKING order="3" place="3" resultid="3856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1337" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4105" />
                    <RANKING order="2" place="2" resultid="3404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1338" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1339" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3745" />
                    <RANKING order="2" place="2" resultid="2042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1340" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1341" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4013" />
                    <RANKING order="2" place="2" resultid="2813" />
                    <RANKING order="3" place="3" resultid="2412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1342" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="1343" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="1344" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2103" />
                    <RANKING order="2" place="2" resultid="2112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1346" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1347" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1348" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1349" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1350" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1351" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4353" daytime="11:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4354" daytime="11:19" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1352" daytime="11:24" gender="M" number="17" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1353" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1873" />
                    <RANKING order="2" place="2" resultid="2274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1355" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2509" />
                    <RANKING order="2" place="2" resultid="3794" />
                    <RANKING order="3" place="-1" resultid="2851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1356" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3868" />
                    <RANKING order="2" place="2" resultid="1894" />
                    <RANKING order="3" place="-1" resultid="3948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1357" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3280" />
                    <RANKING order="2" place="2" resultid="4168" />
                    <RANKING order="3" place="-1" resultid="3129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1358" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1847" />
                    <RANKING order="2" place="2" resultid="3666" />
                    <RANKING order="3" place="3" resultid="3335" />
                    <RANKING order="4" place="4" resultid="3509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1359" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4044" />
                    <RANKING order="2" place="2" resultid="2610" />
                    <RANKING order="3" place="3" resultid="1914" />
                    <RANKING order="4" place="4" resultid="2252" />
                    <RANKING order="5" place="5" resultid="3975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1360" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1974" />
                    <RANKING order="2" place="2" resultid="3360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1361" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3309" />
                    <RANKING order="2" place="2" resultid="3882" />
                    <RANKING order="3" place="3" resultid="2033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1362" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2702" />
                    <RANKING order="2" place="2" resultid="3682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1363" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3463" />
                    <RANKING order="2" place="2" resultid="3957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1364" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1365" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1366" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1367" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1368" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4355" daytime="11:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4356" daytime="11:31" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4357" daytime="11:35" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1369" daytime="11:39" gender="F" number="18" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1772" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="1773" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1774" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3050" />
                    <RANKING order="2" place="2" resultid="2448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1775" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4022" />
                    <RANKING order="2" place="2" resultid="1919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1776" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1777" agemax="279" agemin="240" calculate="TOTAL" />
                <AGEGROUP agegroupid="1778" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4490" daytime="11:39" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1386" daytime="11:43" gender="M" number="19" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1779" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="1780" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1781" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3051" />
                    <RANKING order="2" place="2" resultid="1920" />
                    <RANKING order="3" place="3" resultid="4247" />
                    <RANKING order="4" place="4" resultid="4190" />
                    <RANKING order="5" place="5" resultid="3191" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1782" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4189" />
                    <RANKING order="2" place="2" resultid="5044" />
                    <RANKING order="3" place="3" resultid="3828" />
                    <RANKING order="4" place="4" resultid="3052" />
                    <RANKING order="5" place="5" resultid="4237" />
                    <RANKING order="6" place="6" resultid="1921" />
                    <RANKING order="7" place="7" resultid="2450" />
                    <RANKING order="8" place="-1" resultid="3145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1783" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3354" />
                    <RANKING order="2" place="2" resultid="2451" />
                    <RANKING order="3" place="3" resultid="5045" />
                    <RANKING order="4" place="4" resultid="3053" />
                    <RANKING order="5" place="5" resultid="2122" />
                    <RANKING order="6" place="6" resultid="1922" />
                    <RANKING order="7" place="7" resultid="1980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1784" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1785" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2452" />
                    <RANKING order="2" place="2" resultid="4089" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4491" daytime="11:43" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4492" daytime="11:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4493" daytime="11:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2022-06-11" daytime="16:00" endtime="20:05" name="SOBOTA" number="3">
          <EVENTS>
            <EVENT eventid="1404" daytime="16:00" gender="F" number="20" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1408" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2467" />
                    <RANKING order="2" place="2" resultid="3926" />
                    <RANKING order="3" place="3" resultid="3300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1409" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2792" />
                    <RANKING order="2" place="2" resultid="3492" />
                    <RANKING order="3" place="3" resultid="2406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2979" />
                    <RANKING order="2" place="2" resultid="3048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2548" />
                    <RANKING order="2" place="2" resultid="3501" />
                    <RANKING order="3" place="3" resultid="2827" />
                    <RANKING order="4" place="4" resultid="2068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1412" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2492" />
                    <RANKING order="2" place="2" resultid="3819" />
                    <RANKING order="3" place="3" resultid="4003" />
                    <RANKING order="4" place="4" resultid="2539" />
                    <RANKING order="5" place="5" resultid="2313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3044" />
                    <RANKING order="2" place="2" resultid="2871" />
                    <RANKING order="3" place="3" resultid="2299" />
                    <RANKING order="4" place="4" resultid="5041" />
                    <RANKING order="5" place="5" resultid="2323" />
                    <RANKING order="6" place="6" resultid="2335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1961" />
                    <RANKING order="2" place="2" resultid="3812" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1415" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2052" />
                    <RANKING order="2" place="2" resultid="3328" />
                    <RANKING order="3" place="3" resultid="3187" />
                    <RANKING order="4" place="-1" resultid="3020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1417" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1418" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3243" />
                    <RANKING order="2" place="2" resultid="2529" />
                    <RANKING order="3" place="3" resultid="4081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1420" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1421" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1422" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1423" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4362" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4363" daytime="16:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4364" daytime="16:09" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4365" daytime="16:12" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1406" daytime="16:14" gender="M" number="21" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1424" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3485" />
                    <RANKING order="2" place="2" resultid="3420" />
                    <RANKING order="3" place="3" resultid="2841" />
                    <RANKING order="4" place="4" resultid="3254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3714" />
                    <RANKING order="2" place="2" resultid="4123" />
                    <RANKING order="3" place="3" resultid="3598" />
                    <RANKING order="4" place="4" resultid="2240" />
                    <RANKING order="5" place="-1" resultid="2852" />
                    <RANKING order="6" place="-1" resultid="3969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3527" />
                    <RANKING order="2" place="2" resultid="2985" />
                    <RANKING order="3" place="3" resultid="2935" />
                    <RANKING order="4" place="4" resultid="3137" />
                    <RANKING order="5" place="5" resultid="3910" />
                    <RANKING order="6" place="6" resultid="1895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4162" />
                    <RANKING order="2" place="2" resultid="2351" />
                    <RANKING order="3" place="3" resultid="4206" />
                    <RANKING order="4" place="4" resultid="1911" />
                    <RANKING order="5" place="5" resultid="3767" />
                    <RANKING order="6" place="6" resultid="2400" />
                    <RANKING order="7" place="-1" resultid="3444" />
                    <RANKING order="8" place="-1" resultid="1882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3003" />
                    <RANKING order="2" place="2" resultid="3518" />
                    <RANKING order="3" place="3" resultid="3350" />
                    <RANKING order="4" place="4" resultid="2265" />
                    <RANKING order="5" place="5" resultid="1841" />
                    <RANKING order="6" place="6" resultid="2426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2293" />
                    <RANKING order="2" place="2" resultid="4199" />
                    <RANKING order="3" place="3" resultid="1834" />
                    <RANKING order="4" place="4" resultid="3709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1431" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2667" />
                    <RANKING order="2" place="2" resultid="2806" />
                    <RANKING order="3" place="3" resultid="2888" />
                    <RANKING order="4" place="4" resultid="1952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1432" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2822" />
                    <RANKING order="2" place="2" resultid="3100" />
                    <RANKING order="3" place="3" resultid="3982" />
                    <RANKING order="4" place="4" resultid="2437" />
                    <RANKING order="5" place="5" resultid="2383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2703" />
                    <RANKING order="2" place="2" resultid="3890" />
                    <RANKING order="3" place="3" resultid="2375" />
                    <RANKING order="4" place="4" resultid="2082" />
                    <RANKING order="5" place="-1" resultid="2831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3015" />
                    <RANKING order="2" place="2" resultid="3918" />
                    <RANKING order="3" place="3" resultid="2420" />
                    <RANKING order="4" place="4" resultid="3342" />
                    <RANKING order="5" place="5" resultid="2432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1435" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3645" />
                    <RANKING order="2" place="2" resultid="3577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1436" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4063" />
                    <RANKING order="2" place="2" resultid="3235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1437" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1438" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1439" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4366" daytime="16:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4367" daytime="16:19" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4368" daytime="16:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4369" daytime="16:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4370" daytime="16:29" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4371" daytime="16:31" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1440" daytime="16:33" gender="F" number="22" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1441" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2635" />
                    <RANKING order="2" place="2" resultid="3301" />
                    <RANKING order="3" place="3" resultid="3927" />
                    <RANKING order="4" place="-1" resultid="3857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2522" />
                    <RANKING order="2" place="2" resultid="3262" />
                    <RANKING order="3" place="3" resultid="3397" />
                    <RANKING order="4" place="4" resultid="2129" />
                    <RANKING order="5" place="5" resultid="4106" />
                    <RANKING order="6" place="6" resultid="3405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3266" />
                    <RANKING order="2" place="2" resultid="3270" />
                    <RANKING order="3" place="3" resultid="2980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3455" />
                    <RANKING order="2" place="2" resultid="2060" />
                    <RANKING order="3" place="3" resultid="2075" />
                    <RANKING order="4" place="4" resultid="3820" />
                    <RANKING order="5" place="5" resultid="2991" />
                    <RANKING order="6" place="6" resultid="4224" />
                    <RANKING order="7" place="7" resultid="3801" />
                    <RANKING order="8" place="8" resultid="2441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2814" />
                    <RANKING order="2" place="2" resultid="4007" />
                    <RANKING order="3" place="3" resultid="3676" />
                    <RANKING order="4" place="-1" resultid="2340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2330" />
                    <RANKING order="2" place="2" resultid="3840" />
                    <RANKING order="3" place="3" resultid="3813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3329" />
                    <RANKING order="2" place="2" resultid="3616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2307" />
                    <RANKING order="2" place="2" resultid="2113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1451" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1452" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1453" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1454" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1455" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1456" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4372" daytime="16:33" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4373" daytime="16:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4374" daytime="16:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4375" daytime="16:39" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1457" daytime="16:41" gender="M" number="23" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1458" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3733" />
                    <RANKING order="2" place="2" resultid="2624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4143" />
                    <RANKING order="2" place="2" resultid="1874" />
                    <RANKING order="3" place="3" resultid="3371" />
                    <RANKING order="4" place="4" resultid="2218" />
                    <RANKING order="5" place="5" resultid="2838" />
                    <RANKING order="6" place="6" resultid="2283" />
                    <RANKING order="7" place="7" resultid="3565" />
                    <RANKING order="8" place="8" resultid="2842" />
                    <RANKING order="9" place="9" resultid="3388" />
                    <RANKING order="10" place="10" resultid="2941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1460" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3182" />
                    <RANKING order="2" place="2" resultid="4185" />
                    <RANKING order="3" place="3" resultid="3161" />
                    <RANKING order="4" place="4" resultid="2774" />
                    <RANKING order="5" place="5" resultid="3379" />
                    <RANKING order="6" place="6" resultid="3795" />
                    <RANKING order="7" place="-1" resultid="2853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1461" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3604" />
                    <RANKING order="2" place="2" resultid="3119" />
                    <RANKING order="3" place="3" resultid="2228" />
                    <RANKING order="4" place="4" resultid="2798" />
                    <RANKING order="5" place="5" resultid="4147" />
                    <RANKING order="6" place="6" resultid="3206" />
                    <RANKING order="7" place="7" resultid="3845" />
                    <RANKING order="8" place="8" resultid="3911" />
                    <RANKING order="9" place="9" resultid="1896" />
                    <RANKING order="10" place="10" resultid="4241" />
                    <RANKING order="11" place="11" resultid="3198" />
                    <RANKING order="12" place="12" resultid="2359" />
                    <RANKING order="13" place="-1" resultid="2249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1462" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2785" />
                    <RANKING order="2" place="2" resultid="2734" />
                    <RANKING order="3" place="3" resultid="2729" />
                    <RANKING order="4" place="4" resultid="3130" />
                    <RANKING order="5" place="5" resultid="2957" />
                    <RANKING order="6" place="6" resultid="3150" />
                    <RANKING order="7" place="7" resultid="3827" />
                    <RANKING order="8" place="8" resultid="3626" />
                    <RANKING order="9" place="-1" resultid="3031" />
                    <RANKING order="10" place="-1" resultid="3106" />
                    <RANKING order="11" place="-1" resultid="3142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1463" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1848" />
                    <RANKING order="2" place="2" resultid="3351" />
                    <RANKING order="3" place="3" resultid="4233" />
                    <RANKING order="4" place="4" resultid="2671" />
                    <RANKING order="5" place="5" resultid="2652" />
                    <RANKING order="6" place="6" resultid="2391" />
                    <RANKING order="7" place="-1" resultid="1857" />
                    <RANKING order="8" place="-1" resultid="2928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1464" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2097" />
                    <RANKING order="2" place="2" resultid="2611" />
                    <RANKING order="3" place="3" resultid="3907" />
                    <RANKING order="4" place="4" resultid="4045" />
                    <RANKING order="5" place="5" resultid="2212" />
                    <RANKING order="6" place="6" resultid="2253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2748" />
                    <RANKING order="2" place="2" resultid="2916" />
                    <RANKING order="3" place="3" resultid="3659" />
                    <RANKING order="4" place="4" resultid="3212" />
                    <RANKING order="5" place="5" resultid="3171" />
                    <RANKING order="6" place="6" resultid="1975" />
                    <RANKING order="7" place="7" resultid="2950" />
                    <RANKING order="8" place="-1" resultid="3953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1466" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2090" />
                    <RANKING order="2" place="2" resultid="2756" />
                    <RANKING order="3" place="3" resultid="3983" />
                    <RANKING order="4" place="4" resultid="2034" />
                    <RANKING order="5" place="5" resultid="3638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2376" />
                    <RANKING order="2" place="2" resultid="3684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1468" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3919" />
                    <RANKING order="2" place="2" resultid="4059" />
                    <RANKING order="3" place="3" resultid="3550" />
                    <RANKING order="4" place="4" resultid="3229" />
                    <RANKING order="5" place="5" resultid="4250" />
                    <RANKING order="6" place="-1" resultid="3473" />
                    <RANKING order="7" place="-1" resultid="3835" />
                    <RANKING order="8" place="-1" resultid="4086" />
                    <RANKING order="9" place="-1" resultid="2367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1469" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3646" />
                    <RANKING order="2" place="2" resultid="4053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1470" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1471" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1472" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1473" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4376" daytime="16:41" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4377" daytime="16:43" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4378" daytime="16:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4379" daytime="16:47" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4380" daytime="16:49" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4381" daytime="16:51" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4382" daytime="16:52" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4383" daytime="16:54" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4384" daytime="16:55" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1474" daytime="16:57" gender="F" number="24" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1475" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1476" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2523" />
                    <RANKING order="2" place="2" resultid="2974" />
                    <RANKING order="3" place="3" resultid="2620" />
                    <RANKING order="4" place="4" resultid="3157" />
                    <RANKING order="5" place="-1" resultid="2473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1477" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4264" />
                    <RANKING order="2" place="2" resultid="2647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1478" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3291" />
                    <RANKING order="2" place="2" resultid="3746" />
                    <RANKING order="3" place="3" resultid="3502" />
                    <RANKING order="4" place="4" resultid="2549" />
                    <RANKING order="5" place="5" resultid="2069" />
                    <RANKING order="6" place="6" resultid="1944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1479" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2061" />
                    <RANKING order="2" place="2" resultid="3456" />
                    <RANKING order="3" place="3" resultid="2540" />
                    <RANKING order="4" place="-1" resultid="1812" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1480" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4011" />
                    <RANKING order="2" place="2" resultid="1829" />
                    <RANKING order="3" place="3" resultid="2260" />
                    <RANKING order="4" place="-1" resultid="2300" />
                    <RANKING order="5" place="-1" resultid="2341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2319" />
                    <RANKING order="2" place="2" resultid="3536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2053" />
                    <RANKING order="2" place="2" resultid="2740" />
                    <RANKING order="3" place="3" resultid="4136" />
                    <RANKING order="4" place="4" resultid="3021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2104" />
                    <RANKING order="2" place="2" resultid="3222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1484" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2714" />
                    <RANKING order="2" place="2" resultid="3559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1485" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2867" />
                    <RANKING order="2" place="2" resultid="3244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1486" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4077" />
                    <RANKING order="2" place="2" resultid="3692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1487" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1488" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1489" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1490" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4385" daytime="16:57" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4386" daytime="17:01" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4387" daytime="17:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4388" daytime="17:10" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1491" daytime="17:13" gender="M" number="25" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1492" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2719" />
                    <RANKING order="2" place="2" resultid="3863" />
                    <RANKING order="3" place="3" resultid="3413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3380" />
                    <RANKING order="2" place="2" resultid="2241" />
                    <RANKING order="3" place="3" resultid="2119" />
                    <RANKING order="4" place="4" resultid="2510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1495" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1496" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3032" />
                    <RANKING order="2" place="2" resultid="2786" />
                    <RANKING order="3" place="3" resultid="4177" />
                    <RANKING order="4" place="4" resultid="2678" />
                    <RANKING order="5" place="5" resultid="3542" />
                    <RANKING order="6" place="6" resultid="2401" />
                    <RANKING order="7" place="-1" resultid="3107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1497" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3336" />
                    <RANKING order="2" place="2" resultid="4154" />
                    <RANKING order="3" place="3" resultid="2222" />
                    <RANKING order="4" place="4" resultid="4234" />
                    <RANKING order="5" place="5" resultid="2672" />
                    <RANKING order="6" place="6" resultid="1903" />
                    <RANKING order="7" place="7" resultid="2266" />
                    <RANKING order="8" place="8" resultid="3481" />
                    <RANKING order="9" place="9" resultid="3510" />
                    <RANKING order="10" place="10" resultid="3786" />
                    <RANKING order="11" place="-1" resultid="3319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1498" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4046" />
                    <RANKING order="2" place="2" resultid="3672" />
                    <RANKING order="3" place="3" resultid="2279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1499" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2917" />
                    <RANKING order="2" place="2" resultid="4129" />
                    <RANKING order="3" place="3" resultid="3660" />
                    <RANKING order="4" place="4" resultid="3808" />
                    <RANKING order="5" place="5" resultid="3361" />
                    <RANKING order="6" place="6" resultid="1968" />
                    <RANKING order="7" place="7" resultid="2443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1500" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2091" />
                    <RANKING order="2" place="2" resultid="3101" />
                    <RANKING order="3" place="3" resultid="3883" />
                    <RANKING order="4" place="4" resultid="2384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2923" />
                    <RANKING order="2" place="2" resultid="2882" />
                    <RANKING order="3" place="3" resultid="2484" />
                    <RANKING order="4" place="-1" resultid="3761" />
                    <RANKING order="5" place="-1" resultid="4257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1502" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3343" />
                    <RANKING order="2" place="2" resultid="2875" />
                    <RANKING order="3" place="3" resultid="3464" />
                    <RANKING order="4" place="4" resultid="2433" />
                    <RANKING order="5" place="-1" resultid="3836" />
                    <RANKING order="6" place="-1" resultid="4087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1503" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4054" />
                    <RANKING order="2" place="2" resultid="3086" />
                    <RANKING order="3" place="3" resultid="3578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1504" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3236" />
                    <RANKING order="2" place="2" resultid="3066" />
                    <RANKING order="3" place="3" resultid="3571" />
                    <RANKING order="4" place="4" resultid="3700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1505" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1506" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1507" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4389" daytime="17:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4390" daytime="17:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4391" daytime="17:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4392" daytime="17:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4393" daytime="17:28" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4394" daytime="17:30" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1508" daytime="17:33" gender="F" number="26" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1509" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2130" />
                    <RANKING order="2" place="2" resultid="3398" />
                    <RANKING order="3" place="3" resultid="3406" />
                    <RANKING order="4" place="4" resultid="3493" />
                    <RANKING order="5" place="5" resultid="2629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1511" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2648" />
                    <RANKING order="2" place="2" resultid="4017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1512" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3292" />
                    <RANKING order="2" place="2" resultid="3850" />
                    <RANKING order="3" place="3" resultid="3115" />
                    <RANKING order="4" place="4" resultid="3034" />
                    <RANKING order="5" place="5" resultid="1945" />
                    <RANKING order="6" place="-1" resultid="2043" />
                    <RANKING order="7" place="-1" resultid="4245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1513" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3653" />
                    <RANKING order="2" place="2" resultid="3124" />
                    <RANKING order="3" place="3" resultid="2076" />
                    <RANKING order="4" place="4" resultid="2992" />
                    <RANKING order="5" place="5" resultid="4225" />
                    <RANKING order="6" place="-1" resultid="1813" />
                    <RANKING order="7" place="-1" resultid="3802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1514" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4008" />
                    <RANKING order="2" place="2" resultid="3632" />
                    <RANKING order="3" place="3" resultid="2413" />
                    <RANKING order="4" place="4" resultid="5042" />
                    <RANKING order="5" place="-1" resultid="2206" />
                    <RANKING order="6" place="-1" resultid="3073" />
                    <RANKING order="7" place="-1" resultid="2324" />
                    <RANKING order="8" place="-1" resultid="4014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3874" />
                    <RANKING order="2" place="2" resultid="1821" />
                    <RANKING order="3" place="3" resultid="2741" />
                    <RANKING order="4" place="4" resultid="4137" />
                    <RANKING order="5" place="5" resultid="3617" />
                    <RANKING order="6" place="6" resultid="4019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2105" />
                    <RANKING order="2" place="2" resultid="3223" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1518" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1519" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1520" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1521" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1522" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1523" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1524" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4395" daytime="17:33" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4396" daytime="17:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4397" daytime="17:43" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4398" daytime="17:47" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1525" daytime="17:51" gender="M" number="27" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1526" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1527" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3372" />
                    <RANKING order="2" place="2" resultid="2275" />
                    <RANKING order="3" place="3" resultid="3041" />
                    <RANKING order="4" place="4" resultid="2284" />
                    <RANKING order="5" place="5" resultid="3389" />
                    <RANKING order="6" place="6" resultid="3593" />
                    <RANKING order="7" place="-1" resultid="2942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1528" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3991" />
                    <RANKING order="2" place="2" resultid="4186" />
                    <RANKING order="3" place="3" resultid="3781" />
                    <RANKING order="4" place="4" resultid="3610" />
                    <RANKING order="5" place="5" resultid="2846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1529" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3605" />
                    <RANKING order="2" place="2" resultid="2799" />
                    <RANKING order="3" place="3" resultid="2229" />
                    <RANKING order="4" place="4" resultid="4148" />
                    <RANKING order="5" place="5" resultid="3177" />
                    <RANKING order="6" place="6" resultid="2396" />
                    <RANKING order="7" place="7" resultid="2360" />
                    <RANKING order="8" place="-1" resultid="3199" />
                    <RANKING order="9" place="-1" resultid="3207" />
                    <RANKING order="10" place="-1" resultid="3528" />
                    <RANKING order="11" place="-1" resultid="3846" />
                    <RANKING order="12" place="-1" resultid="3902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1530" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3281" />
                    <RANKING order="2" place="2" resultid="1865" />
                    <RANKING order="3" place="3" resultid="2962" />
                    <RANKING order="4" place="4" resultid="4169" />
                    <RANKING order="5" place="5" resultid="2352" />
                    <RANKING order="6" place="6" resultid="3131" />
                    <RANKING order="7" place="7" resultid="4207" />
                    <RANKING order="8" place="8" resultid="3448" />
                    <RANKING order="9" place="9" resultid="2605" />
                    <RANKING order="10" place="10" resultid="3588" />
                    <RANKING order="11" place="-1" resultid="1883" />
                    <RANKING order="12" place="-1" resultid="2945" />
                    <RANKING order="13" place="-1" resultid="3202" />
                    <RANKING order="14" place="-1" resultid="3931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1531" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3218" />
                    <RANKING order="2" place="2" resultid="4155" />
                    <RANKING order="3" place="3" resultid="3519" />
                    <RANKING order="4" place="4" resultid="3895" />
                    <RANKING order="5" place="5" resultid="3004" />
                    <RANKING order="6" place="6" resultid="1904" />
                    <RANKING order="7" place="7" resultid="2653" />
                    <RANKING order="8" place="8" resultid="3511" />
                    <RANKING order="9" place="9" resultid="1858" />
                    <RANKING order="10" place="10" resultid="1842" />
                    <RANKING order="11" place="11" resultid="3787" />
                    <RANKING order="12" place="-1" resultid="2500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1532" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3091" />
                    <RANKING order="2" place="2" resultid="4215" />
                    <RANKING order="3" place="3" resultid="2213" />
                    <RANKING order="4" place="4" resultid="2860" />
                    <RANKING order="5" place="5" resultid="1915" />
                    <RANKING order="6" place="6" resultid="2896" />
                    <RANKING order="7" place="7" resultid="2254" />
                    <RANKING order="8" place="8" resultid="1835" />
                    <RANKING order="9" place="-1" resultid="3721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1533" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2749" />
                    <RANKING order="2" place="2" resultid="4130" />
                    <RANKING order="3" place="3" resultid="3078" />
                    <RANKING order="4" place="4" resultid="3213" />
                    <RANKING order="5" place="5" resultid="3775" />
                    <RANKING order="6" place="6" resultid="1953" />
                    <RANKING order="7" place="7" resultid="1969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1534" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2907" />
                    <RANKING order="2" place="2" resultid="2757" />
                    <RANKING order="3" place="3" resultid="3310" />
                    <RANKING order="4" place="4" resultid="2035" />
                    <RANKING order="5" place="-1" resultid="2660" />
                    <RANKING order="6" place="-1" resultid="4239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1535" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4095" />
                    <RANKING order="2" place="2" resultid="3755" />
                    <RANKING order="3" place="3" resultid="2485" />
                    <RANKING order="4" place="4" resultid="2083" />
                    <RANKING order="5" place="-1" resultid="4258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1536" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3551" />
                    <RANKING order="2" place="2" resultid="2368" />
                    <RANKING order="3" place="3" resultid="3474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1537" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1538" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3067" />
                    <RANKING order="2" place="2" resultid="3701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1539" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1540" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1541" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4399" daytime="17:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4400" daytime="17:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4401" daytime="18:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4402" daytime="18:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4403" daytime="18:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4404" daytime="18:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4405" daytime="18:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4406" daytime="18:28" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4407" daytime="18:32" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1542" daytime="18:35" gender="F" number="28" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1786" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="1787" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1788" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3054" />
                    <RANKING order="2" place="2" resultid="2453" />
                    <RANKING order="3" place="-1" resultid="1923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1789" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2123" />
                    <RANKING order="2" place="2" resultid="4024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1790" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1791" agemax="279" agemin="240" calculate="TOTAL" />
                <AGEGROUP agegroupid="1792" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4494" daytime="18:35" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1559" daytime="18:38" gender="M" number="29" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1793" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="1794" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1795" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3055" />
                    <RANKING order="2" place="2" resultid="4246" />
                    <RANKING order="3" place="3" resultid="3192" />
                    <RANKING order="4" place="4" resultid="3056" />
                    <RANKING order="5" place="-1" resultid="1924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1796" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4191" />
                    <RANKING order="2" place="2" resultid="5047" />
                    <RANKING order="3" place="3" resultid="2516" />
                    <RANKING order="4" place="4" resultid="4238" />
                    <RANKING order="5" place="5" resultid="1925" />
                    <RANKING order="6" place="6" resultid="2455" />
                    <RANKING order="7" place="-1" resultid="3829" />
                    <RANKING order="8" place="-1" resultid="3146" />
                    <RANKING order="9" place="-1" resultid="4023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1797" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3355" />
                    <RANKING order="2" place="2" resultid="3057" />
                    <RANKING order="3" place="3" resultid="5046" />
                    <RANKING order="4" place="4" resultid="2456" />
                    <RANKING order="5" place="5" resultid="1926" />
                    <RANKING order="6" place="-1" resultid="1981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1798" agemax="279" agemin="240" calculate="TOTAL" />
                <AGEGROUP agegroupid="1799" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2457" />
                    <RANKING order="2" place="2" resultid="4090" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4495" daytime="18:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4496" daytime="18:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4497" daytime="18:45" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1576" daytime="18:48" gender="F" number="30" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1577" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2468" />
                    <RANKING order="2" place="2" resultid="3935" />
                    <RANKING order="3" place="-1" resultid="3858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1578" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4107" />
                    <RANKING order="2" place="2" resultid="2407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1579" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1580" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3747" />
                    <RANKING order="2" place="2" resultid="2044" />
                    <RANKING order="3" place="3" resultid="3035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1581" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1582" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2815" />
                    <RANKING order="2" place="2" resultid="2414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="1584" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1586" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1587" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1588" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1589" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1590" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1591" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1592" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4412" daytime="18:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4413" daytime="18:56" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1593" daytime="19:04" gender="M" number="31" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1594" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3438" />
                    <RANKING order="2" place="-1" resultid="3944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1595" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2778" />
                    <RANKING order="2" place="2" resultid="1875" />
                    <RANKING order="3" place="3" resultid="3421" />
                    <RANKING order="4" place="4" resultid="3414" />
                    <RANKING order="5" place="-1" resultid="3255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1596" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3599" />
                    <RANKING order="2" place="2" resultid="4049" />
                    <RANKING order="3" place="3" resultid="3796" />
                    <RANKING order="4" place="-1" resultid="2511" />
                    <RANKING order="5" place="-1" resultid="2847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1597" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3282" />
                    <RANKING order="2" place="2" resultid="1866" />
                    <RANKING order="3" place="3" resultid="2679" />
                    <RANKING order="4" place="4" resultid="3543" />
                    <RANKING order="5" place="-1" resultid="4163" />
                    <RANKING order="6" place="-1" resultid="4178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1849" />
                    <RANKING order="2" place="2" resultid="3667" />
                    <RANKING order="3" place="-1" resultid="2968" />
                    <RANKING order="4" place="-1" resultid="2427" />
                    <RANKING order="5" place="-1" resultid="3320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2612" />
                    <RANKING order="2" place="2" resultid="4216" />
                    <RANKING order="3" place="3" resultid="3974" />
                    <RANKING order="4" place="-1" resultid="2861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2807" />
                    <RANKING order="2" place="2" resultid="3362" />
                    <RANKING order="3" place="3" resultid="1976" />
                    <RANKING order="4" place="4" resultid="2951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3311" />
                    <RANKING order="2" place="2" resultid="1889" />
                    <RANKING order="3" place="3" resultid="3671" />
                    <RANKING order="4" place="-1" resultid="2661" />
                    <RANKING order="5" place="-1" resultid="2908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2704" />
                    <RANKING order="2" place="2" resultid="3685" />
                    <RANKING order="3" place="-1" resultid="2883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3016" />
                    <RANKING order="2" place="2" resultid="3465" />
                    <RANKING order="3" place="3" resultid="3960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1606" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1607" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1608" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1609" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4414" daytime="19:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4415" daytime="19:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4416" daytime="19:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4417" daytime="19:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4418" daytime="19:40" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2022-06-12" daytime="09:00" name="NIEDZIELA" number="4">
          <EVENTS>
            <EVENT eventid="1611" daytime="09:00" gender="F" number="32" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1613" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2469" />
                    <RANKING order="2" place="2" resultid="2636" />
                    <RANKING order="3" place="3" resultid="3302" />
                    <RANKING order="4" place="-1" resultid="3859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1614" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4108" />
                    <RANKING order="2" place="2" resultid="3399" />
                    <RANKING order="3" place="3" resultid="3407" />
                    <RANKING order="4" place="-1" resultid="2524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1615" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1616" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3748" />
                    <RANKING order="2" place="2" resultid="3116" />
                    <RANKING order="3" place="3" resultid="2045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1617" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2077" />
                    <RANKING order="2" place="2" resultid="2993" />
                    <RANKING order="3" place="3" resultid="4004" />
                    <RANKING order="4" place="4" resultid="3803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4012" />
                    <RANKING order="2" place="2" resultid="2816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1620" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1621" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2308" />
                    <RANKING order="2" place="2" resultid="2106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1622" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1623" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1624" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1625" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1626" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1627" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1628" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4419" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4420" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4421" daytime="09:06" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1629" daytime="09:08" gender="M" number="33" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1630" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2724" />
                    <RANKING order="2" place="2" resultid="3735" />
                    <RANKING order="3" place="3" resultid="2625" />
                    <RANKING order="4" place="-1" resultid="3945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1631" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3373" />
                    <RANKING order="2" place="2" resultid="3042" />
                    <RANKING order="3" place="3" resultid="1876" />
                    <RANKING order="4" place="4" resultid="3566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1632" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2848" />
                    <RANKING order="2" place="2" resultid="4187" />
                    <RANKING order="3" place="3" resultid="3600" />
                    <RANKING order="4" place="4" resultid="3797" />
                    <RANKING order="5" place="-1" resultid="2854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3606" />
                    <RANKING order="2" place="2" resultid="3120" />
                    <RANKING order="3" place="3" resultid="2800" />
                    <RANKING order="4" place="4" resultid="4149" />
                    <RANKING order="5" place="5" resultid="1897" />
                    <RANKING order="6" place="6" resultid="2361" />
                    <RANKING order="7" place="-1" resultid="2230" />
                    <RANKING order="8" place="-1" resultid="3026" />
                    <RANKING order="9" place="-1" resultid="3949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2787" />
                    <RANKING order="2" place="2" resultid="3132" />
                    <RANKING order="3" place="3" resultid="4170" />
                    <RANKING order="4" place="4" resultid="3151" />
                    <RANKING order="5" place="-1" resultid="2735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1850" />
                    <RANKING order="2" place="2" resultid="3352" />
                    <RANKING order="3" place="3" resultid="4235" />
                    <RANKING order="4" place="4" resultid="2673" />
                    <RANKING order="5" place="5" resultid="2969" />
                    <RANKING order="6" place="6" resultid="2929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3092" />
                    <RANKING order="2" place="2" resultid="2613" />
                    <RANKING order="3" place="3" resultid="2255" />
                    <RANKING order="4" place="4" resultid="3976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2918" />
                    <RANKING order="2" place="2" resultid="3661" />
                    <RANKING order="3" place="3" resultid="1977" />
                    <RANKING order="4" place="-1" resultid="2952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1638" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3984" />
                    <RANKING order="2" place="2" resultid="2036" />
                    <RANKING order="3" place="-1" resultid="2092" />
                    <RANKING order="4" place="-1" resultid="2909" />
                    <RANKING order="5" place="-1" resultid="3885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1639" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2705" />
                    <RANKING order="2" place="2" resultid="3686" />
                    <RANKING order="3" place="3" resultid="2377" />
                    <RANKING order="4" place="4" resultid="2486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1640" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3921" />
                    <RANKING order="2" place="2" resultid="3466" />
                    <RANKING order="3" place="3" resultid="3959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1641" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1642" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1643" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1644" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1645" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4422" daytime="09:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4423" daytime="09:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4424" daytime="09:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4425" daytime="09:19" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4426" daytime="09:21" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4427" daytime="09:23" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1646" daytime="09:25" gender="F" number="34" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1647" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2477" />
                    <RANKING order="2" place="-1" resultid="3860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1648" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2474" />
                    <RANKING order="2" place="2" resultid="2630" />
                    <RANKING order="3" place="-1" resultid="2975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1649" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3293" />
                    <RANKING order="2" place="2" resultid="3749" />
                    <RANKING order="3" place="3" resultid="3503" />
                    <RANKING order="4" place="4" resultid="3851" />
                    <RANKING order="5" place="5" resultid="1946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2062" />
                    <RANKING order="2" place="2" resultid="4111" />
                    <RANKING order="3" place="3" resultid="1814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5037" />
                    <RANKING order="2" place="2" resultid="2817" />
                    <RANKING order="3" place="3" resultid="2261" />
                    <RANKING order="4" place="4" resultid="2415" />
                    <RANKING order="5" place="-1" resultid="2301" />
                    <RANKING order="6" place="-1" resultid="3074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1653" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1654" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4138" />
                    <RANKING order="2" place="2" resultid="1823" />
                    <RANKING order="3" place="-1" resultid="2742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1655" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3224" />
                    <RANKING order="2" place="2" resultid="2115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1656" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2715" />
                    <RANKING order="2" place="2" resultid="3560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1657" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1658" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4078" />
                    <RANKING order="2" place="2" resultid="3695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1659" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1660" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1661" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1662" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4428" daytime="09:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4429" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4430" daytime="09:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4431" daytime="09:55" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1663" daytime="10:00" gender="M" number="35" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1664" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3439" />
                    <RANKING order="2" place="-1" resultid="3946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1665" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2720" />
                    <RANKING order="2" place="2" resultid="2276" />
                    <RANKING order="3" place="3" resultid="3864" />
                    <RANKING order="4" place="4" resultid="1877" />
                    <RANKING order="5" place="5" resultid="3415" />
                    <RANKING order="6" place="-1" resultid="3256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1666" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3381" />
                    <RANKING order="2" place="2" resultid="3970" />
                    <RANKING order="3" place="3" resultid="2242" />
                    <RANKING order="4" place="-1" resultid="2512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1667" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1668" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2788" />
                    <RANKING order="2" place="2" resultid="4179" />
                    <RANKING order="3" place="3" resultid="1867" />
                    <RANKING order="4" place="3" resultid="2680" />
                    <RANKING order="5" place="5" resultid="3544" />
                    <RANKING order="6" place="-1" resultid="2946" />
                    <RANKING order="7" place="-1" resultid="3108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4156" />
                    <RANKING order="2" place="2" resultid="3337" />
                    <RANKING order="3" place="3" resultid="2674" />
                    <RANKING order="4" place="4" resultid="2223" />
                    <RANKING order="5" place="5" resultid="3321" />
                    <RANKING order="6" place="6" resultid="1905" />
                    <RANKING order="7" place="7" resultid="3482" />
                    <RANKING order="8" place="8" resultid="3512" />
                    <RANKING order="9" place="9" resultid="3788" />
                    <RANKING order="10" place="-1" resultid="3896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1670" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3097" />
                    <RANKING order="2" place="2" resultid="4217" />
                    <RANKING order="3" place="3" resultid="4047" />
                    <RANKING order="4" place="4" resultid="2897" />
                    <RANKING order="5" place="-1" resultid="2280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1671" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2919" />
                    <RANKING order="2" place="2" resultid="4131" />
                    <RANKING order="3" place="3" resultid="3809" />
                    <RANKING order="4" place="4" resultid="3363" />
                    <RANKING order="5" place="5" resultid="1970" />
                    <RANKING order="6" place="6" resultid="2444" />
                    <RANKING order="7" place="7" resultid="1978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1672" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2093" />
                    <RANKING order="2" place="2" resultid="3312" />
                    <RANKING order="3" place="3" resultid="2758" />
                    <RANKING order="4" place="4" resultid="2662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1673" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2924" />
                    <RANKING order="2" place="2" resultid="2884" />
                    <RANKING order="3" place="3" resultid="3687" />
                    <RANKING order="4" place="-1" resultid="4259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1674" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3344" />
                    <RANKING order="2" place="2" resultid="2421" />
                    <RANKING order="3" place="3" resultid="3467" />
                    <RANKING order="4" place="-1" resultid="2876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1675" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4055" />
                    <RANKING order="2" place="2" resultid="3579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1676" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3068" />
                    <RANKING order="2" place="2" resultid="3702" />
                    <RANKING order="3" place="-1" resultid="3572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1677" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1678" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1679" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4432" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4433" daytime="10:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4434" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4435" daytime="10:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4436" daytime="10:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4437" daytime="10:24" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1680" daytime="10:27" gender="F" number="36" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1681" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1682" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2793" />
                    <RANKING order="2" place="2" resultid="3494" />
                    <RANKING order="3" place="3" resultid="3400" />
                    <RANKING order="4" place="4" resultid="2131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1683" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1684" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2550" />
                    <RANKING order="2" place="2" resultid="3504" />
                    <RANKING order="3" place="3" resultid="3036" />
                    <RANKING order="4" place="4" resultid="2828" />
                    <RANKING order="5" place="5" resultid="2070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1685" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2493" />
                    <RANKING order="2" place="2" resultid="2063" />
                    <RANKING order="3" place="3" resultid="4226" />
                    <RANKING order="4" place="4" resultid="3125" />
                    <RANKING order="5" place="5" resultid="3821" />
                    <RANKING order="6" place="6" resultid="2541" />
                    <RANKING order="7" place="7" resultid="2314" />
                    <RANKING order="8" place="-1" resultid="3457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1686" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2302" />
                    <RANKING order="2" place="2" resultid="3633" />
                    <RANKING order="3" place="3" resultid="2207" />
                    <RANKING order="4" place="4" resultid="2325" />
                    <RANKING order="5" place="5" resultid="2336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1687" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1963" />
                    <RANKING order="2" place="2" resultid="3814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1688" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2054" />
                    <RANKING order="2" place="2" resultid="3188" />
                    <RANKING order="3" place="3" resultid="3331" />
                    <RANKING order="4" place="4" resultid="3082" />
                    <RANKING order="5" place="5" resultid="3618" />
                    <RANKING order="6" place="-1" resultid="3022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1689" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1690" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1691" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3245" />
                    <RANKING order="2" place="2" resultid="2532" />
                    <RANKING order="3" place="3" resultid="4082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1692" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4072" />
                    <RANKING order="2" place="2" resultid="3994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1693" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1694" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1695" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1696" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4438" daytime="10:27" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4439" daytime="10:31" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4440" daytime="10:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4441" daytime="10:36" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1697" daytime="10:37" gender="M" number="37" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1698" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1699" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3486" />
                    <RANKING order="2" place="2" resultid="3422" />
                    <RANKING order="3" place="3" resultid="2843" />
                    <RANKING order="4" place="4" resultid="3257" />
                    <RANKING order="5" place="5" resultid="3390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1700" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3715" />
                    <RANKING order="2" place="2" resultid="4124" />
                    <RANKING order="3" place="3" resultid="3601" />
                    <RANKING order="4" place="4" resultid="3162" />
                    <RANKING order="5" place="5" resultid="2120" />
                    <RANKING order="6" place="6" resultid="2243" />
                    <RANKING order="7" place="-1" resultid="2513" />
                    <RANKING order="8" place="-1" resultid="2855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1701" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2986" />
                    <RANKING order="2" place="2" resultid="3529" />
                    <RANKING order="3" place="3" resultid="2936" />
                    <RANKING order="4" place="4" resultid="3138" />
                    <RANKING order="5" place="5" resultid="3912" />
                    <RANKING order="6" place="6" resultid="3950" />
                    <RANKING order="7" place="7" resultid="1898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1702" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4164" />
                    <RANKING order="2" place="2" resultid="2353" />
                    <RANKING order="3" place="3" resultid="3283" />
                    <RANKING order="4" place="4" resultid="4180" />
                    <RANKING order="5" place="5" resultid="3768" />
                    <RANKING order="6" place="6" resultid="1912" />
                    <RANKING order="7" place="7" resultid="4208" />
                    <RANKING order="8" place="8" resultid="2958" />
                    <RANKING order="9" place="9" resultid="2402" />
                    <RANKING order="10" place="10" resultid="3627" />
                    <RANKING order="11" place="-1" resultid="1884" />
                    <RANKING order="12" place="-1" resultid="2730" />
                    <RANKING order="13" place="-1" resultid="3143" />
                    <RANKING order="14" place="-1" resultid="3445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1703" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3005" />
                    <RANKING order="2" place="2" resultid="3353" />
                    <RANKING order="3" place="3" resultid="3520" />
                    <RANKING order="4" place="4" resultid="4236" />
                    <RANKING order="5" place="5" resultid="3322" />
                    <RANKING order="6" place="6" resultid="2267" />
                    <RANKING order="7" place="7" resultid="2428" />
                    <RANKING order="8" place="8" resultid="2654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1704" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2294" />
                    <RANKING order="2" place="2" resultid="2098" />
                    <RANKING order="3" place="3" resultid="4200" />
                    <RANKING order="4" place="4" resultid="1836" />
                    <RANKING order="5" place="5" resultid="2281" />
                    <RANKING order="6" place="6" resultid="2256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1705" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2750" />
                    <RANKING order="2" place="2" resultid="2668" />
                    <RANKING order="3" place="3" resultid="2808" />
                    <RANKING order="4" place="4" resultid="3662" />
                    <RANKING order="5" place="5" resultid="2889" />
                    <RANKING order="6" place="6" resultid="1954" />
                    <RANKING order="7" place="-1" resultid="3172" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1706" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2823" />
                    <RANKING order="2" place="2" resultid="3102" />
                    <RANKING order="3" place="3" resultid="2438" />
                    <RANKING order="4" place="4" resultid="3985" />
                    <RANKING order="5" place="5" resultid="2385" />
                    <RANKING order="6" place="-1" resultid="3886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1707" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4096" />
                    <RANKING order="2" place="2" resultid="3891" />
                    <RANKING order="3" place="3" resultid="2706" />
                    <RANKING order="4" place="4" resultid="2378" />
                    <RANKING order="5" place="5" resultid="2084" />
                    <RANKING order="6" place="-1" resultid="2832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1708" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3017" />
                    <RANKING order="2" place="2" resultid="3922" />
                    <RANKING order="3" place="3" resultid="2422" />
                    <RANKING order="4" place="4" resultid="3345" />
                    <RANKING order="5" place="5" resultid="2434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1709" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3648" />
                    <RANKING order="2" place="2" resultid="3580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1710" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4065" />
                    <RANKING order="2" place="2" resultid="3237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1711" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1712" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1713" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4442" daytime="10:37" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4443" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4444" daytime="10:43" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4445" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4446" daytime="10:46" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4447" daytime="10:48" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4448" daytime="10:50" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4449" daytime="10:51" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1714" daytime="10:53" gender="X" number="38" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1800" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="1801" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1802" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3058" />
                    <RANKING order="2" place="2" resultid="1927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1803" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3147" />
                    <RANKING order="2" place="2" resultid="2458" />
                    <RANKING order="3" place="3" resultid="2517" />
                    <RANKING order="4" place="4" resultid="2124" />
                    <RANKING order="5" place="5" resultid="1928" />
                    <RANKING order="6" place="6" resultid="4248" />
                    <RANKING order="7" place="7" resultid="3193" />
                    <RANKING order="8" place="8" resultid="1982" />
                    <RANKING order="9" place="-1" resultid="3059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1804" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1805" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1806" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3247" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4498" daytime="10:53" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4499" daytime="10:56" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1731" daytime="11:00" gender="F" number="39" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1732" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2470" />
                    <RANKING order="2" place="2" resultid="3936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1733" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2132" />
                    <RANKING order="2" place="2" resultid="4109" />
                    <RANKING order="3" place="3" resultid="3408" />
                    <RANKING order="4" place="4" resultid="5105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1734" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1735" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3294" />
                    <RANKING order="2" place="2" resultid="4244" />
                    <RANKING order="3" place="3" resultid="2551" />
                    <RANKING order="4" place="4" resultid="2046" />
                    <RANKING order="5" place="5" resultid="3037" />
                    <RANKING order="6" place="6" resultid="1947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1736" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3654" />
                    <RANKING order="2" place="2" resultid="2994" />
                    <RANKING order="3" place="3" resultid="3822" />
                    <RANKING order="4" place="4" resultid="4227" />
                    <RANKING order="5" place="5" resultid="1815" />
                    <RANKING order="6" place="6" resultid="2542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1737" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3634" />
                    <RANKING order="2" place="2" resultid="2416" />
                    <RANKING order="3" place="3" resultid="5043" />
                    <RANKING order="4" place="-1" resultid="4009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1738" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1964" />
                    <RANKING order="2" place="2" resultid="3538" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1739" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3875" />
                    <RANKING order="2" place="2" resultid="1824" />
                    <RANKING order="3" place="3" resultid="4139" />
                    <RANKING order="4" place="4" resultid="3189" />
                    <RANKING order="5" place="5" resultid="4020" />
                    <RANKING order="6" place="-1" resultid="3619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1740" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2107" />
                    <RANKING order="2" place="2" resultid="3225" />
                    <RANKING order="3" place="3" resultid="2116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1741" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1742" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1743" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1744" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1745" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1746" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1747" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4452" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4453" daytime="11:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4454" daytime="11:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4455" daytime="11:28" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1748" daytime="11:35" gender="M" number="40" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1749" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1750" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2779" />
                    <RANKING order="2" place="2" resultid="2285" />
                    <RANKING order="3" place="3" resultid="3374" />
                    <RANKING order="4" place="4" resultid="3594" />
                    <RANKING order="5" place="5" resultid="3416" />
                    <RANKING order="6" place="6" resultid="3391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1751" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4188" />
                    <RANKING order="2" place="2" resultid="3971" />
                    <RANKING order="3" place="3" resultid="3382" />
                    <RANKING order="4" place="4" resultid="3798" />
                    <RANKING order="5" place="-1" resultid="3992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1752" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2801" />
                    <RANKING order="2" place="2" resultid="2231" />
                    <RANKING order="3" place="3" resultid="3027" />
                    <RANKING order="4" place="4" resultid="3870" />
                    <RANKING order="5" place="5" resultid="3530" />
                    <RANKING order="6" place="6" resultid="2515" />
                    <RANKING order="7" place="7" resultid="4240" />
                    <RANKING order="8" place="8" resultid="2362" />
                    <RANKING order="9" place="-1" resultid="2937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1753" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3284" />
                    <RANKING order="2" place="2" resultid="1868" />
                    <RANKING order="3" place="3" resultid="2963" />
                    <RANKING order="4" place="4" resultid="4171" />
                    <RANKING order="5" place="5" resultid="4209" />
                    <RANKING order="6" place="6" resultid="2681" />
                    <RANKING order="7" place="7" resultid="2504" />
                    <RANKING order="8" place="8" resultid="3545" />
                    <RANKING order="9" place="-1" resultid="2354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1754" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1851" />
                    <RANKING order="2" place="2" resultid="4157" />
                    <RANKING order="3" place="3" resultid="3219" />
                    <RANKING order="4" place="4" resultid="3897" />
                    <RANKING order="5" place="5" resultid="3521" />
                    <RANKING order="6" place="6" resultid="1906" />
                    <RANKING order="7" place="7" resultid="3006" />
                    <RANKING order="8" place="8" resultid="2930" />
                    <RANKING order="9" place="9" resultid="3789" />
                    <RANKING order="10" place="10" resultid="1843" />
                    <RANKING order="11" place="11" resultid="2429" />
                    <RANKING order="12" place="12" resultid="2392" />
                    <RANKING order="13" place="-1" resultid="1859" />
                    <RANKING order="14" place="-1" resultid="2970" />
                    <RANKING order="15" place="-1" resultid="3513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1755" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3093" />
                    <RANKING order="2" place="2" resultid="4218" />
                    <RANKING order="3" place="3" resultid="2214" />
                    <RANKING order="4" place="4" resultid="4048" />
                    <RANKING order="5" place="5" resultid="2614" />
                    <RANKING order="6" place="6" resultid="1916" />
                    <RANKING order="7" place="7" resultid="4201" />
                    <RANKING order="8" place="8" resultid="2898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1756" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3079" />
                    <RANKING order="2" place="2" resultid="2809" />
                    <RANKING order="3" place="3" resultid="3214" />
                    <RANKING order="4" place="4" resultid="3776" />
                    <RANKING order="5" place="5" resultid="2953" />
                    <RANKING order="6" place="6" resultid="1955" />
                    <RANKING order="7" place="7" resultid="1971" />
                    <RANKING order="8" place="-1" resultid="3364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1757" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3313" />
                    <RANKING order="2" place="2" resultid="1890" />
                    <RANKING order="3" place="3" resultid="2663" />
                    <RANKING order="4" place="-1" resultid="2037" />
                    <RANKING order="5" place="-1" resultid="2910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1758" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3756" />
                    <RANKING order="2" place="2" resultid="2487" />
                    <RANKING order="3" place="-1" resultid="2885" />
                    <RANKING order="4" place="-1" resultid="3011" />
                    <RANKING order="5" place="-1" resultid="4260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1759" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3552" />
                    <RANKING order="2" place="2" resultid="2369" />
                    <RANKING order="3" place="3" resultid="2877" />
                    <RANKING order="4" place="4" resultid="3475" />
                    <RANKING order="5" place="5" resultid="3958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1760" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1761" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1762" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1763" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1764" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4456" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4457" daytime="11:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4458" daytime="11:47" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4459" daytime="11:53" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4460" daytime="12:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4461" daytime="12:08" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4462" daytime="12:18" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4463" daytime="12:34" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="02211" nation="POL" region="11" clubid="2290" name="MUKS Gilus Gilowice">
          <ATHLETES>
            <ATHLETE firstname="Sławomir" lastname="Formas" birthdate="1969-11-05" gender="M" nation="POL" license="502211700187" swrid="4292540" athleteid="2291">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1250" points="803" reactiontime="+84" swimtime="00:02:38.85" resultid="2292" heatid="4329" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:55.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1406" points="812" reactiontime="+81" swimtime="00:01:11.16" resultid="2293" heatid="4366" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1697" points="804" reactiontime="+83" swimtime="00:00:32.43" resultid="2294" heatid="4443" lane="0" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02902" nation="POL" region="02" clubid="2600" name="Uks Czwórka Nakło">
          <ATHLETES>
            <ATHLETE firstname="Radosław" lastname="Staszkiewicz" birthdate="1968-04-21" gender="M" nation="POL" license="102902700326" swrid="5337392" athleteid="2606">
              <RESULTS>
                <RESULT eventid="1112" points="413" reactiontime="+119" swimtime="00:02:56.18" resultid="2607" heatid="4295" lane="9" entrytime="00:02:58.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:21.53" />
                    <SPLIT distance="150" swimtime="00:02:15.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1197" points="434" reactiontime="+125" swimtime="00:22:38.47" resultid="2608" heatid="4311" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:19.99" />
                    <SPLIT distance="150" swimtime="00:02:04.34" />
                    <SPLIT distance="200" swimtime="00:02:49.82" />
                    <SPLIT distance="250" swimtime="00:03:35.16" />
                    <SPLIT distance="300" swimtime="00:04:20.60" />
                    <SPLIT distance="350" swimtime="00:05:06.44" />
                    <SPLIT distance="400" swimtime="00:05:52.50" />
                    <SPLIT distance="450" swimtime="00:06:38.79" />
                    <SPLIT distance="500" swimtime="00:07:25.30" />
                    <SPLIT distance="550" swimtime="00:08:11.43" />
                    <SPLIT distance="600" swimtime="00:08:58.11" />
                    <SPLIT distance="650" swimtime="00:09:43.90" />
                    <SPLIT distance="700" swimtime="00:10:29.86" />
                    <SPLIT distance="750" swimtime="00:11:15.85" />
                    <SPLIT distance="800" swimtime="00:12:01.99" />
                    <SPLIT distance="850" swimtime="00:12:47.72" />
                    <SPLIT distance="900" swimtime="00:13:33.30" />
                    <SPLIT distance="950" swimtime="00:14:18.90" />
                    <SPLIT distance="1000" swimtime="00:15:04.49" />
                    <SPLIT distance="1050" swimtime="00:15:50.28" />
                    <SPLIT distance="1100" swimtime="00:16:36.39" />
                    <SPLIT distance="1150" swimtime="00:17:21.49" />
                    <SPLIT distance="1200" swimtime="00:18:07.24" />
                    <SPLIT distance="1250" swimtime="00:18:53.14" />
                    <SPLIT distance="1300" swimtime="00:19:39.52" />
                    <SPLIT distance="1350" swimtime="00:20:25.45" />
                    <SPLIT distance="1400" swimtime="00:21:10.92" />
                    <SPLIT distance="1450" swimtime="00:21:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="385" reactiontime="+94" swimtime="00:00:39.28" resultid="2609" heatid="4319" lane="6" />
                <RESULT eventid="1352" points="364" reactiontime="+115" swimtime="00:03:06.80" resultid="2610" heatid="4356" lane="7" entrytime="00:03:14.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:24.20" />
                    <SPLIT distance="150" swimtime="00:02:15.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="517" reactiontime="+99" swimtime="00:00:32.24" resultid="2611" heatid="4377" lane="5" />
                <RESULT eventid="1593" points="428" reactiontime="+114" swimtime="00:06:18.90" resultid="2612" heatid="4418" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:25.31" />
                    <SPLIT distance="150" swimtime="00:02:16.00" />
                    <SPLIT distance="200" swimtime="00:03:04.95" />
                    <SPLIT distance="250" swimtime="00:03:59.24" />
                    <SPLIT distance="300" swimtime="00:04:54.88" />
                    <SPLIT distance="350" swimtime="00:05:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="383" reactiontime="+125" swimtime="00:01:18.79" resultid="2613" heatid="4424" lane="6" entrytime="00:01:23.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="415" reactiontime="+105" swimtime="00:05:43.04" resultid="2614" heatid="4460" lane="4" entrytime="00:05:41.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:19.36" />
                    <SPLIT distance="150" swimtime="00:02:02.51" />
                    <SPLIT distance="200" swimtime="00:02:47.25" />
                    <SPLIT distance="250" swimtime="00:03:32.43" />
                    <SPLIT distance="300" swimtime="00:04:18.17" />
                    <SPLIT distance="350" swimtime="00:05:02.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Spychalski" birthdate="1980-09-05" gender="M" nation="POL" license="102902700357" swrid="5337379" athleteid="2601">
              <RESULTS>
                <RESULT eventid="1076" points="419" reactiontime="+80" swimtime="00:00:31.06" resultid="2602" heatid="4281" lane="9" entrytime="00:00:29.88" entrycourse="LCM" />
                <RESULT eventid="1163" points="424" reactiontime="+91" swimtime="00:11:26.56" resultid="2603" heatid="4307" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:58.83" />
                    <SPLIT distance="200" swimtime="00:02:42.16" />
                    <SPLIT distance="250" swimtime="00:03:25.58" />
                    <SPLIT distance="300" swimtime="00:04:09.85" />
                    <SPLIT distance="350" swimtime="00:04:54.74" />
                    <SPLIT distance="400" swimtime="00:05:38.47" />
                    <SPLIT distance="450" swimtime="00:06:22.16" />
                    <SPLIT distance="500" swimtime="00:07:06.14" />
                    <SPLIT distance="550" swimtime="00:07:50.78" />
                    <SPLIT distance="600" swimtime="00:08:34.71" />
                    <SPLIT distance="650" swimtime="00:09:19.17" />
                    <SPLIT distance="700" swimtime="00:10:03.68" />
                    <SPLIT distance="750" swimtime="00:10:46.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="408" reactiontime="+86" swimtime="00:01:09.03" resultid="2604" heatid="4352" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="385" reactiontime="+81" swimtime="00:02:36.23" resultid="2605" heatid="4400" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="150" swimtime="00:01:55.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3770" name="UŚKS Ostrołęka">
          <ATHLETES>
            <ATHLETE firstname="ADAM" lastname="JANCZEWSKI " birthdate="1990-01-01" gender="M" nation="POL" athleteid="3986">
              <RESULTS>
                <RESULT eventid="1076" points="665" reactiontime="+79" swimtime="00:00:25.35" resultid="3987" heatid="4286" lane="6" entrytime="00:00:25.00" />
                <RESULT eventid="1112" points="607" reactiontime="+87" swimtime="00:02:24.29" resultid="3988" heatid="4297" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                    <SPLIT distance="100" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:51.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="593" reactiontime="+88" swimtime="00:09:41.51" resultid="3989" heatid="4303" lane="7" entrytime="00:09:50.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:45.03" />
                    <SPLIT distance="200" swimtime="00:02:22.65" />
                    <SPLIT distance="250" swimtime="00:02:59.66" />
                    <SPLIT distance="300" swimtime="00:03:37.07" />
                    <SPLIT distance="350" swimtime="00:04:13.84" />
                    <SPLIT distance="400" swimtime="00:04:50.84" />
                    <SPLIT distance="450" swimtime="00:05:27.59" />
                    <SPLIT distance="500" swimtime="00:06:04.73" />
                    <SPLIT distance="550" swimtime="00:06:41.70" />
                    <SPLIT distance="600" swimtime="00:07:19.05" />
                    <SPLIT distance="650" swimtime="00:07:55.85" />
                    <SPLIT distance="700" swimtime="00:08:32.52" />
                    <SPLIT distance="750" swimtime="00:09:08.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="722" reactiontime="+89" swimtime="00:00:55.52" resultid="3990" heatid="4351" lane="5" entrytime="00:00:56.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="654" reactiontime="+90" swimtime="00:02:06.25" resultid="3991" heatid="4407" lane="2" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="100" swimtime="00:01:01.77" />
                    <SPLIT distance="150" swimtime="00:01:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="3992" heatid="4456" lane="0" entrytime="00:04:41.43" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="TOMASZ" lastname="AMBROZIAK" birthdate="1964-01-01" gender="M" nation="POL" athleteid="3771">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3772" heatid="4278" lane="1" entrytime="00:00:33.90" />
                <RESULT eventid="1112" points="247" reactiontime="+89" swimtime="00:03:44.34" resultid="3773" heatid="4293" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                    <SPLIT distance="100" swimtime="00:01:51.42" />
                    <SPLIT distance="150" swimtime="00:02:53.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" status="WDR" swimtime="00:00:00.00" resultid="3774" entrytime="00:01:30.00" />
                <RESULT eventid="1525" points="251" reactiontime="+89" swimtime="00:03:16.61" resultid="3775" heatid="4401" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:03:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="221" reactiontime="+82" swimtime="00:07:14.34" resultid="3776" heatid="4461" lane="6" entrytime="00:07:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:38.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4050" name="Weteran  Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW.JANA  4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE firstname="Daniel" lastname="Fecica" birthdate="1940-11-29" gender="M" nation="POL" license="102611700018" swrid="4102523" athleteid="4060">
              <RESULTS>
                <RESULT eventid="1076" points="418" swimtime="00:00:42.75" resultid="4061" heatid="4276" lane="8" entrytime="00:00:45.00" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1250" points="606" swimtime="00:04:05.40" resultid="4062" heatid="4331" lane="7" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.94" />
                    <SPLIT distance="100" swimtime="00:02:00.85" />
                    <SPLIT distance="150" swimtime="00:03:05.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="558" reactiontime="+85" swimtime="00:01:54.71" resultid="4063" heatid="4367" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="245" reactiontime="+106" swimtime="00:00:55.55" resultid="4064" heatid="4378" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1697" points="534" reactiontime="+112" swimtime="00:00:51.39" resultid="4065" heatid="4444" lane="9" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernard" lastname="Poloczek" birthdate="1947-02-25" gender="M" nation="POL" license="102611700032" swrid="4792004" athleteid="4051">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1267" points="426" reactiontime="+75" swimtime="00:00:45.77" resultid="4052" heatid="4321" lane="8" entrytime="00:00:45.58" />
                <RESULT eventid="1457" points="345" reactiontime="+85" swimtime="00:00:45.29" resultid="4053" heatid="4379" lane="8" entrytime="00:00:44.69" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1491" points="423" reactiontime="+78" swimtime="00:01:42.81" resultid="4054" heatid="4391" lane="8" entrytime="00:01:42.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="380" reactiontime="+81" swimtime="00:03:54.96" resultid="4055" heatid="4434" lane="8" entrytime="00:03:48.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.18" />
                    <SPLIT distance="100" swimtime="00:01:51.15" />
                    <SPLIT distance="150" swimtime="00:02:52.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Bosowski" birthdate="1948-05-22" gender="M" nation="POL" license="102611700014" swrid="4129761" athleteid="4083">
              <RESULTS>
                <RESULT eventid="1076" points="168" reactiontime="+110" swimtime="00:00:50.26" resultid="4084" heatid="4276" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1267" points="102" reactiontime="+117" swimtime="00:01:11.91" resultid="4085" heatid="4320" lane="8" entrytime="00:01:05.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="4086" heatid="4378" lane="1" entrytime="00:01:05.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="4087" heatid="4390" lane="6" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Renata" lastname="Bastek" birthdate="1943-12-02" gender="F" nation="POL" license="102611600023" swrid="4223066" athleteid="4073">
              <RESULTS>
                <RESULT eventid="1059" points="505" reactiontime="+84" swimtime="00:00:42.83" resultid="4074" heatid="4267" lane="3" />
                <RESULT eventid="1215" points="471" reactiontime="+74" swimtime="00:00:51.53" resultid="4075" heatid="4313" lane="2" />
                <RESULT eventid="1284" points="454" reactiontime="+86" swimtime="00:01:40.67" resultid="4076" heatid="4335" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="434" reactiontime="+80" swimtime="00:01:57.11" resultid="4077" heatid="4386" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="445" reactiontime="+74" swimtime="00:04:17.82" resultid="4078" heatid="4428" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.66" />
                    <SPLIT distance="100" swimtime="00:02:11.12" />
                    <SPLIT distance="150" swimtime="00:03:16.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Genowefa" lastname="Drużyńska" birthdate="1951-02-10" gender="F" nation="POL" license="102611600033" swrid="4655173" athleteid="4079">
              <RESULTS>
                <RESULT eventid="1233" points="223" reactiontime="+102" swimtime="00:05:45.32" resultid="4080" heatid="4327" lane="0" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.99" />
                    <SPLIT distance="100" swimtime="00:02:46.54" />
                    <SPLIT distance="150" swimtime="00:04:18.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="201" reactiontime="+98" swimtime="00:02:43.76" resultid="4081" heatid="4363" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="254" reactiontime="+105" swimtime="00:01:05.78" resultid="4082" heatid="4439" lane="2" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystyna" lastname="Fecica" birthdate="1943-03-12" gender="F" nation="POL" license="102611600019" swrid="4102524" athleteid="4066">
              <RESULTS>
                <RESULT eventid="1146" points="430" reactiontime="+137" swimtime="00:17:12.37" resultid="4067" heatid="4301" lane="6" entrytime="00:18:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.84" />
                    <SPLIT distance="100" swimtime="00:02:00.83" />
                    <SPLIT distance="150" swimtime="00:03:05.90" />
                    <SPLIT distance="200" swimtime="00:04:11.08" />
                    <SPLIT distance="250" swimtime="00:05:16.41" />
                    <SPLIT distance="300" swimtime="00:06:21.59" />
                    <SPLIT distance="350" swimtime="00:07:27.70" />
                    <SPLIT distance="400" swimtime="00:08:33.27" />
                    <SPLIT distance="450" swimtime="00:09:39.55" />
                    <SPLIT distance="500" swimtime="00:10:44.40" />
                    <SPLIT distance="550" swimtime="00:11:50.60" />
                    <SPLIT distance="600" swimtime="00:12:55.98" />
                    <SPLIT distance="650" swimtime="00:14:00.54" />
                    <SPLIT distance="700" swimtime="00:15:05.88" />
                    <SPLIT distance="750" swimtime="00:16:10.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="487" reactiontime="+113" swimtime="00:04:40.72" resultid="4068" heatid="4327" lane="1" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.39" />
                    <SPLIT distance="100" swimtime="00:02:11.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="530" reactiontime="+109" swimtime="00:02:02.10" resultid="4069" heatid="4363" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="356" reactiontime="+114" swimtime="00:00:54.93" resultid="4070" heatid="4373" lane="1" entrytime="00:00:56.00" />
                <RESULT eventid="1611" points="442" reactiontime="+113" swimtime="00:02:04.52" resultid="4071" heatid="4420" lane="0" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="489" reactiontime="+119" swimtime="00:00:55.77" resultid="4072" heatid="4439" lane="5" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiesław" lastname="Kornicki" birthdate="1949-01-28" gender="M" nation="POL" license="102611700015" swrid="4137183" athleteid="4056">
              <RESULTS>
                <RESULT eventid="1076" points="507" reactiontime="+90" swimtime="00:00:34.76" resultid="4057" heatid="4277" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1301" points="420" reactiontime="+93" swimtime="00:01:24.56" resultid="4058" heatid="4345" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="432" reactiontime="+88" swimtime="00:00:39.66" resultid="4059" heatid="4379" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1386" reactiontime="+71" swimtime="00:03:15.97" resultid="4089" heatid="4491" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.74" />
                    <SPLIT distance="100" swimtime="00:01:42.33" />
                    <SPLIT distance="150" swimtime="00:02:28.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4051" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4060" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4056" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="4083" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1559" reactiontime="+94" swimtime="00:02:49.14" resultid="4090" heatid="4495" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="100" swimtime="00:01:29.74" />
                    <SPLIT distance="150" swimtime="00:02:13.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4051" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="4083" number="2" />
                    <RELAYPOSITION athleteid="4060" number="3" reactiontime="+83" />
                    <RELAYPOSITION athleteid="4056" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" swimtime="00:02:58.60" resultid="4088" heatid="4488" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.33" />
                    <SPLIT distance="100" swimtime="00:01:34.57" />
                    <SPLIT distance="150" swimtime="00:02:19.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4066" number="1" />
                    <RELAYPOSITION athleteid="4073" number="2" />
                    <RELAYPOSITION athleteid="4060" number="3" />
                    <RELAYPOSITION athleteid="4056" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" clubid="4039" name="KS. Górnik Radlin">
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Kubica" birthdate="1972-02-22" gender="M" nation="POL" license="100211700343" swrid="5398297" athleteid="4040">
              <RESULTS>
                <RESULT eventid="1076" points="537" reactiontime="+82" swimtime="00:00:29.62" resultid="4041" heatid="4281" lane="2" entrytime="00:00:29.12" />
                <RESULT eventid="1197" points="422" reactiontime="+98" swimtime="00:22:51.08" resultid="4042" heatid="4310" lane="4" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:21.84" />
                    <SPLIT distance="150" swimtime="00:02:06.45" />
                    <SPLIT distance="200" swimtime="00:02:51.34" />
                    <SPLIT distance="250" swimtime="00:03:36.10" />
                    <SPLIT distance="300" swimtime="00:04:21.39" />
                    <SPLIT distance="350" swimtime="00:05:07.01" />
                    <SPLIT distance="400" swimtime="00:05:53.26" />
                    <SPLIT distance="450" swimtime="00:06:39.62" />
                    <SPLIT distance="500" swimtime="00:07:26.30" />
                    <SPLIT distance="550" swimtime="00:08:12.84" />
                    <SPLIT distance="600" swimtime="00:08:59.33" />
                    <SPLIT distance="650" swimtime="00:09:45.52" />
                    <SPLIT distance="700" swimtime="00:10:32.08" />
                    <SPLIT distance="750" swimtime="00:11:18.17" />
                    <SPLIT distance="800" swimtime="00:12:04.60" />
                    <SPLIT distance="850" swimtime="00:12:50.59" />
                    <SPLIT distance="900" swimtime="00:13:37.13" />
                    <SPLIT distance="950" swimtime="00:14:23.65" />
                    <SPLIT distance="1000" swimtime="00:15:10.05" />
                    <SPLIT distance="1050" swimtime="00:15:56.19" />
                    <SPLIT distance="1100" swimtime="00:16:42.87" />
                    <SPLIT distance="1150" swimtime="00:17:29.61" />
                    <SPLIT distance="1200" swimtime="00:18:16.00" />
                    <SPLIT distance="1250" swimtime="00:19:02.23" />
                    <SPLIT distance="1300" swimtime="00:19:48.49" />
                    <SPLIT distance="1350" swimtime="00:20:35.19" />
                    <SPLIT distance="1400" swimtime="00:21:21.24" />
                    <SPLIT distance="1450" swimtime="00:22:07.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="502" reactiontime="+84" swimtime="00:00:35.95" resultid="4043" heatid="4322" lane="3" entrytime="00:00:37.51" />
                <RESULT eventid="1352" points="388" reactiontime="+99" swimtime="00:03:02.78" resultid="4044" heatid="4356" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="150" swimtime="00:02:10.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="508" reactiontime="+80" swimtime="00:00:32.44" resultid="4045" heatid="4381" lane="0" entrytime="00:00:32.60" />
                <RESULT eventid="1491" points="455" reactiontime="+85" swimtime="00:01:20.05" resultid="4046" heatid="4392" lane="3" entrytime="00:01:20.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="438" reactiontime="+86" swimtime="00:02:57.12" resultid="4047" heatid="4435" lane="7" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:26.11" />
                    <SPLIT distance="150" swimtime="00:02:13.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="417" reactiontime="+97" swimtime="00:05:42.50" resultid="4048" heatid="4460" lane="5" entrytime="00:05:41.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:19.56" />
                    <SPLIT distance="150" swimtime="00:02:03.51" />
                    <SPLIT distance="200" swimtime="00:02:48.66" />
                    <SPLIT distance="250" swimtime="00:03:33.63" />
                    <SPLIT distance="300" swimtime="00:04:19.00" />
                    <SPLIT distance="350" swimtime="00:05:03.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05201" nation="POL" region="01" clubid="2028" name="KS JUST SWIM Jelenia Góra">
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Lipka" birthdate="1958-06-05" gender="M" nation="POL" license="505201700087" swrid="5435204" athleteid="2029">
              <RESULTS>
                <RESULT eventid="1076" points="311" reactiontime="+77" swimtime="00:00:37.22" resultid="2030" heatid="4274" lane="7" />
                <RESULT eventid="1163" points="313" reactiontime="+76" swimtime="00:13:59.32" resultid="2031" heatid="4305" lane="9" entrytime="00:13:40.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                    <SPLIT distance="100" swimtime="00:01:40.06" />
                    <SPLIT distance="150" swimtime="00:02:34.62" />
                    <SPLIT distance="200" swimtime="00:03:30.42" />
                    <SPLIT distance="250" swimtime="00:04:25.80" />
                    <SPLIT distance="300" swimtime="00:07:14.06" />
                    <SPLIT distance="350" swimtime="00:06:17.71" />
                    <SPLIT distance="400" swimtime="00:09:08.37" />
                    <SPLIT distance="450" swimtime="00:10:07.30" />
                    <SPLIT distance="500" swimtime="00:14:55.94" />
                    <SPLIT distance="550" swimtime="00:12:03.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="239" reactiontime="+71" swimtime="00:01:33.07" resultid="2032" heatid="4342" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="218" reactiontime="+106" swimtime="00:03:58.53" resultid="2033" heatid="4355" lane="5" entrytime="00:03:56.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.12" />
                    <SPLIT distance="100" swimtime="00:01:53.57" />
                    <SPLIT distance="150" swimtime="00:02:55.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="255" reactiontime="+89" swimtime="00:00:43.62" resultid="2034" heatid="4379" lane="2" entrytime="00:00:41.75" entrycourse="SCM" />
                <RESULT eventid="1525" points="259" reactiontime="+87" swimtime="00:03:20.34" resultid="2035" heatid="4402" lane="0" entrytime="00:03:10.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="241" reactiontime="+81" swimtime="00:01:39.57" resultid="2036" heatid="4424" lane="9" entrytime="00:01:42.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="2037" heatid="4461" lane="5" entrytime="00:06:40.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Lara" birthdate="1985-06-16" gender="F" nation="POL" license="505201600088" swrid="5435203" athleteid="2038">
              <RESULTS>
                <RESULT eventid="1094" points="263" reactiontime="+96" swimtime="00:03:40.69" resultid="2039" heatid="4288" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.27" />
                    <SPLIT distance="100" swimtime="00:01:55.83" />
                    <SPLIT distance="150" swimtime="00:02:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="368" reactiontime="+96" swimtime="00:12:45.68" resultid="2040" heatid="4300" lane="7" entrytime="00:12:23.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                    <SPLIT distance="100" swimtime="00:01:26.59" />
                    <SPLIT distance="150" swimtime="00:02:13.31" />
                    <SPLIT distance="200" swimtime="00:03:01.83" />
                    <SPLIT distance="250" swimtime="00:03:50.12" />
                    <SPLIT distance="300" swimtime="00:04:40.03" />
                    <SPLIT distance="350" swimtime="00:05:28.90" />
                    <SPLIT distance="400" swimtime="00:06:18.29" />
                    <SPLIT distance="450" swimtime="00:07:06.89" />
                    <SPLIT distance="500" swimtime="00:07:56.17" />
                    <SPLIT distance="550" swimtime="00:08:44.35" />
                    <SPLIT distance="600" swimtime="00:09:33.69" />
                    <SPLIT distance="650" swimtime="00:10:21.99" />
                    <SPLIT distance="700" swimtime="00:11:10.12" />
                    <SPLIT distance="750" swimtime="00:11:58.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="324" reactiontime="+92" swimtime="00:01:24.54" resultid="2041" heatid="4336" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1335" points="224" reactiontime="+102" swimtime="00:03:50.76" resultid="2042" heatid="4353" lane="5" entrytime="00:03:37.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.91" />
                    <SPLIT distance="100" swimtime="00:01:49.82" />
                    <SPLIT distance="150" swimtime="00:02:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="2043" heatid="4396" lane="8" />
                <RESULT eventid="1576" points="271" reactiontime="+95" swimtime="00:07:43.06" resultid="2044" heatid="4413" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.34" />
                    <SPLIT distance="100" swimtime="00:01:50.15" />
                    <SPLIT distance="150" swimtime="00:02:59.69" />
                    <SPLIT distance="200" swimtime="00:04:10.42" />
                    <SPLIT distance="250" swimtime="00:05:08.13" />
                    <SPLIT distance="300" swimtime="00:06:06.67" />
                    <SPLIT distance="350" swimtime="00:06:54.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="213" reactiontime="+97" swimtime="00:01:44.59" resultid="2045" heatid="4419" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="357" reactiontime="+97" swimtime="00:06:15.24" resultid="2046" heatid="4453" lane="3" entrytime="00:06:23.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:01:27.00" />
                    <SPLIT distance="150" swimtime="00:02:13.95" />
                    <SPLIT distance="200" swimtime="00:03:02.00" />
                    <SPLIT distance="250" swimtime="00:03:50.67" />
                    <SPLIT distance="300" swimtime="00:04:39.31" />
                    <SPLIT distance="350" swimtime="00:05:27.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="2525" name="UKP Unia Oświęcim">
          <ATHLETES>
            <ATHLETE firstname="Barbara" lastname="Lipniarska-Skubis" birthdate="1952-07-01" gender="F" nation="POL" license="501006600377" athleteid="2526">
              <RESULTS>
                <RESULT eventid="1233" points="326" reactiontime="+107" swimtime="00:05:03.96" resultid="2527" heatid="4326" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.65" />
                    <SPLIT distance="100" swimtime="00:02:26.39" />
                    <SPLIT distance="150" swimtime="00:03:46.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="160" swimtime="00:02:03.20" resultid="2528" heatid="4335" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="323" swimtime="00:02:19.80" resultid="2529" heatid="4362" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="196" swimtime="00:04:24.62" resultid="2530" heatid="4395" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.81" />
                    <SPLIT distance="100" swimtime="00:02:06.10" />
                    <SPLIT distance="150" swimtime="00:03:17.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="179" swimtime="00:05:00.40" resultid="2531" heatid="4428" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.39" />
                    <SPLIT distance="100" swimtime="00:02:25.98" />
                    <SPLIT distance="150" swimtime="00:03:44.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="280" swimtime="00:01:03.72" resultid="2532" heatid="4439" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4251" name="Masters Radom">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="ZIELEZIŃSKI" birthdate="1953-01-01" gender="M" nation="POL" athleteid="4252">
              <RESULTS>
                <RESULT eventid="1076" reactiontime="+108" status="WDR" swimtime="00:00:00.00" resultid="4253" heatid="4273" lane="5" />
                <RESULT eventid="1163" status="WDR" swimtime="00:00:00.00" resultid="4254" heatid="4307" lane="2" />
                <RESULT eventid="1267" status="WDR" swimtime="00:00:00.00" resultid="4255" heatid="4318" lane="1" />
                <RESULT eventid="1301" status="WDR" swimtime="00:00:00.00" resultid="4256" />
                <RESULT eventid="1491" status="WDR" swimtime="00:00:00.00" resultid="4257" heatid="4389" lane="2" />
                <RESULT eventid="1525" status="WDR" swimtime="00:00:00.00" resultid="4258" heatid="4400" lane="6" />
                <RESULT eventid="1663" status="WDR" swimtime="00:00:00.00" resultid="4259" heatid="4432" lane="5" />
                <RESULT eventid="1748" status="WDR" swimtime="00:00:00.00" resultid="4260" heatid="4462" lane="0" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TRPUL" nation="POL" clubid="3663" name="Uczniowski Klub Sportowy Trójka Puławy">
          <CONTACT name="Gogacz" phone="506694816" />
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Maciejczak" birthdate="1960-07-08" gender="M" nation="POL" athleteid="3668">
              <RESULTS>
                <RESULT eventid="1197" points="323" reactiontime="+110" swimtime="00:26:15.97" resultid="3669" heatid="4310" lane="7" entrytime="00:27:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                    <SPLIT distance="100" swimtime="00:01:30.74" />
                    <SPLIT distance="150" swimtime="00:02:22.68" />
                    <SPLIT distance="200" swimtime="00:03:16.21" />
                    <SPLIT distance="250" swimtime="00:04:10.25" />
                    <SPLIT distance="300" swimtime="00:05:04.25" />
                    <SPLIT distance="350" swimtime="00:05:58.31" />
                    <SPLIT distance="400" swimtime="00:06:52.97" />
                    <SPLIT distance="450" swimtime="00:07:47.07" />
                    <SPLIT distance="500" swimtime="00:08:41.71" />
                    <SPLIT distance="550" swimtime="00:09:36.27" />
                    <SPLIT distance="600" swimtime="00:10:31.41" />
                    <SPLIT distance="650" swimtime="00:11:25.42" />
                    <SPLIT distance="700" swimtime="00:14:10.83" />
                    <SPLIT distance="750" swimtime="00:13:15.55" />
                    <SPLIT distance="800" swimtime="00:16:01.55" />
                    <SPLIT distance="850" swimtime="00:15:06.18" />
                    <SPLIT distance="900" swimtime="00:17:52.90" />
                    <SPLIT distance="950" swimtime="00:16:56.57" />
                    <SPLIT distance="1000" swimtime="00:19:44.58" />
                    <SPLIT distance="1050" swimtime="00:18:49.41" />
                    <SPLIT distance="1100" swimtime="00:21:35.89" />
                    <SPLIT distance="1150" swimtime="00:20:39.81" />
                    <SPLIT distance="1200" swimtime="00:27:07.25" />
                    <SPLIT distance="1250" swimtime="00:22:31.48" />
                    <SPLIT distance="1350" swimtime="00:24:24.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="348" reactiontime="+97" swimtime="00:01:22.18" resultid="3670" heatid="4345" lane="8" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="203" reactiontime="+106" swimtime="00:08:44.06" resultid="3671" heatid="4416" lane="0" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.51" />
                    <SPLIT distance="100" swimtime="00:02:02.48" />
                    <SPLIT distance="150" swimtime="00:03:19.42" />
                    <SPLIT distance="200" swimtime="00:07:05.20" />
                    <SPLIT distance="250" swimtime="00:05:51.24" />
                    <SPLIT distance="300" swimtime="00:08:44.06" />
                    <SPLIT distance="350" swimtime="00:07:55.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" athleteid="3664">
              <RESULTS>
                <RESULT eventid="1197" points="536" reactiontime="+87" swimtime="00:20:29.59" resultid="3665" heatid="4311" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                    <SPLIT distance="100" swimtime="00:01:18.32" />
                    <SPLIT distance="150" swimtime="00:01:59.68" />
                    <SPLIT distance="200" swimtime="00:02:40.36" />
                    <SPLIT distance="250" swimtime="00:03:21.47" />
                    <SPLIT distance="300" swimtime="00:04:02.69" />
                    <SPLIT distance="350" swimtime="00:04:44.03" />
                    <SPLIT distance="400" swimtime="00:05:25.51" />
                    <SPLIT distance="450" swimtime="00:06:06.52" />
                    <SPLIT distance="500" swimtime="00:06:47.13" />
                    <SPLIT distance="550" swimtime="00:07:28.11" />
                    <SPLIT distance="600" swimtime="00:08:08.68" />
                    <SPLIT distance="650" swimtime="00:08:49.98" />
                    <SPLIT distance="700" swimtime="00:09:31.13" />
                    <SPLIT distance="750" swimtime="00:10:12.27" />
                    <SPLIT distance="800" swimtime="00:10:53.02" />
                    <SPLIT distance="850" swimtime="00:11:33.88" />
                    <SPLIT distance="900" swimtime="00:12:15.76" />
                    <SPLIT distance="950" swimtime="00:12:56.75" />
                    <SPLIT distance="1000" swimtime="00:13:37.52" />
                    <SPLIT distance="1050" swimtime="00:14:18.67" />
                    <SPLIT distance="1100" swimtime="00:14:59.88" />
                    <SPLIT distance="1150" swimtime="00:15:41.35" />
                    <SPLIT distance="1200" swimtime="00:16:22.64" />
                    <SPLIT distance="1250" swimtime="00:17:04.00" />
                    <SPLIT distance="1300" swimtime="00:17:45.18" />
                    <SPLIT distance="1350" swimtime="00:18:26.61" />
                    <SPLIT distance="1400" swimtime="00:19:08.88" />
                    <SPLIT distance="1450" swimtime="00:19:50.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="550" reactiontime="+92" swimtime="00:02:34.97" resultid="3666" heatid="4357" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:15.34" />
                    <SPLIT distance="150" swimtime="00:01:55.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="536" reactiontime="+96" swimtime="00:05:49.37" resultid="3667" heatid="4417" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                    <SPLIT distance="100" swimtime="00:01:16.39" />
                    <SPLIT distance="150" swimtime="00:02:06.94" />
                    <SPLIT distance="200" swimtime="00:02:54.98" />
                    <SPLIT distance="250" swimtime="00:03:42.65" />
                    <SPLIT distance="300" swimtime="00:04:31.36" />
                    <SPLIT distance="350" swimtime="00:05:10.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIKRA" nation="POL" clubid="3285" name="Stowarzyszenie Siemacha">
          <CONTACT email="pajka@poczta.onet.eu" name="Palmowska- Latuszek" phone="500044884" />
          <ATHLETES>
            <ATHLETE firstname="Paulina" lastname="Palmowska- Latuszek" birthdate="1985-08-01" gender="F" nation="POL" athleteid="3286">
              <RESULTS>
                <RESULT eventid="1059" points="570" reactiontime="+69" swimtime="00:00:31.33" resultid="3287" heatid="4267" lane="7" />
                <RESULT eventid="1094" points="522" reactiontime="+75" swimtime="00:02:55.69" resultid="3288" heatid="4290" lane="0" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:02:12.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="506" reactiontime="+67" swimtime="00:00:35.92" resultid="3289" heatid="4316" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1284" points="559" reactiontime="+73" swimtime="00:01:10.50" resultid="3290" heatid="4336" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="503" reactiontime="+65" swimtime="00:01:17.63" resultid="3291" heatid="4388" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="497" reactiontime="+67" swimtime="00:02:39.01" resultid="3292" heatid="4398" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:01:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="525" reactiontime="+61" swimtime="00:02:51.36" resultid="3293" heatid="4431" lane="5" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:20.80" />
                    <SPLIT distance="150" swimtime="00:02:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="473" reactiontime="+78" swimtime="00:05:41.62" resultid="3294" heatid="4452" lane="0" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:17.43" />
                    <SPLIT distance="150" swimtime="00:03:30.18" />
                    <SPLIT distance="200" swimtime="00:02:45.63" />
                    <SPLIT distance="300" swimtime="00:04:14.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ada" lastname="Malinowska" birthdate="1999-05-27" gender="F" nation="POL" athleteid="3295">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+77" swimtime="00:00:30.72" resultid="3296" heatid="4272" lane="0" entrytime="00:00:29.99" />
                <RESULT eventid="1094" status="DNS" swimtime="00:00:00.00" resultid="3297" heatid="4288" lane="7" />
                <RESULT eventid="1215" reactiontime="+87" swimtime="00:00:39.83" resultid="3298" heatid="4312" lane="9" />
                <RESULT eventid="1284" reactiontime="+76" swimtime="00:01:10.42" resultid="3299" heatid="4340" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" reactiontime="+66" swimtime="00:01:31.46" resultid="3300" heatid="4363" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" reactiontime="+76" swimtime="00:00:33.46" resultid="3301" heatid="4375" lane="9" entrytime="00:00:31.90" />
                <RESULT eventid="1611" reactiontime="+78" swimtime="00:01:18.69" resultid="3302" heatid="4421" lane="8" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" reactiontime="+77" swimtime="00:00:39.77" resultid="3303" heatid="4441" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03503" nation="POL" region="03" clubid="2234" name="MASTERS Lublin">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Dawidek" birthdate="1986-03-13" gender="M" nation="POL" license="103503700029" athleteid="2244">
              <RESULTS>
                <RESULT eventid="1076" status="WDR" swimtime="00:00:00.00" resultid="2245" heatid="4273" lane="2" />
                <RESULT eventid="1112" status="WDR" swimtime="00:00:00.00" resultid="2246" heatid="4291" lane="3" />
                <RESULT eventid="1267" status="WDR" swimtime="00:00:00.00" resultid="2247" heatid="4319" lane="2" />
                <RESULT eventid="1301" status="WDR" swimtime="00:00:00.00" resultid="2248" />
                <RESULT eventid="1457" status="WDR" swimtime="00:00:00.00" resultid="2249" heatid="4377" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Molenda" birthdate="1971-12-11" gender="M" nation="POL" license="103503700012" athleteid="2250">
              <RESULTS>
                <RESULT eventid="1076" points="315" reactiontime="+98" swimtime="00:00:35.38" resultid="2251" heatid="4275" lane="7" />
                <RESULT eventid="1352" points="167" reactiontime="+116" swimtime="00:04:02.29" resultid="2252" heatid="4355" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.10" />
                    <SPLIT distance="100" swimtime="00:02:02.16" />
                    <SPLIT distance="150" swimtime="00:03:03.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="286" reactiontime="+98" swimtime="00:00:39.30" resultid="2253" heatid="4377" lane="3" />
                <RESULT eventid="1525" points="279" reactiontime="+100" swimtime="00:03:01.44" resultid="2254" heatid="4401" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:24.79" />
                    <SPLIT distance="150" swimtime="00:02:14.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="162" reactiontime="+105" swimtime="00:01:44.90" resultid="2255" heatid="4422" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="255" reactiontime="+100" swimtime="00:00:47.59" resultid="2256" heatid="4443" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Wójcicki" birthdate="1975-04-28" gender="M" nation="POL" license="103503700001" swrid="5455050" athleteid="2262">
              <RESULTS>
                <RESULT eventid="1163" points="355" reactiontime="+94" swimtime="00:12:15.45" resultid="2263" heatid="4307" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:23.58" />
                    <SPLIT distance="150" swimtime="00:02:08.37" />
                    <SPLIT distance="200" swimtime="00:02:53.98" />
                    <SPLIT distance="250" swimtime="00:03:40.26" />
                    <SPLIT distance="300" swimtime="00:04:26.83" />
                    <SPLIT distance="350" swimtime="00:05:13.92" />
                    <SPLIT distance="400" swimtime="00:06:00.57" />
                    <SPLIT distance="450" swimtime="00:06:47.67" />
                    <SPLIT distance="500" swimtime="00:07:35.16" />
                    <SPLIT distance="550" swimtime="00:08:22.24" />
                    <SPLIT distance="600" swimtime="00:09:09.73" />
                    <SPLIT distance="650" swimtime="00:09:56.62" />
                    <SPLIT distance="700" swimtime="00:10:44.04" />
                    <SPLIT distance="750" swimtime="00:11:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="368" reactiontime="+80" swimtime="00:00:38.55" resultid="2264" heatid="4319" lane="0" />
                <RESULT eventid="1406" points="368" reactiontime="+87" swimtime="00:01:30.37" resultid="2265" heatid="4366" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="384" reactiontime="+78" swimtime="00:01:22.76" resultid="2266" heatid="4389" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="389" reactiontime="+78" swimtime="00:00:40.02" resultid="2267" heatid="4442" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Pietrzak" birthdate="1988-10-21" gender="M" nation="POL" license="103503700011" athleteid="2235">
              <RESULTS>
                <RESULT eventid="1076" points="434" reactiontime="+83" swimtime="00:00:29.23" resultid="2236" heatid="4274" lane="6" />
                <RESULT eventid="1163" status="WDR" swimtime="00:00:00.00" resultid="2237" heatid="4306" lane="0" />
                <RESULT eventid="1267" points="410" reactiontime="+90" swimtime="00:00:34.97" resultid="2238" heatid="4319" lane="8" />
                <RESULT eventid="1301" points="385" reactiontime="+83" swimtime="00:01:08.43" resultid="2239" heatid="4342" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="413" reactiontime="+73" swimtime="00:01:22.23" resultid="2240" heatid="4366" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="427" reactiontime="+79" swimtime="00:01:14.26" resultid="2241" heatid="4389" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="371" reactiontime="+78" swimtime="00:02:50.81" resultid="2242" heatid="4433" lane="0">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="385" reactiontime="+92" swimtime="00:00:38.42" resultid="2243" heatid="4443" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Wójcicka" birthdate="1975-05-28" gender="F" nation="POL" license="103503600002" athleteid="2257">
              <RESULTS>
                <RESULT eventid="1146" points="307" reactiontime="+153" swimtime="00:13:37.09" resultid="2258" heatid="4301" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:01:28.15" />
                    <SPLIT distance="150" swimtime="00:02:18.59" />
                    <SPLIT distance="200" swimtime="00:03:10.48" />
                    <SPLIT distance="250" swimtime="00:04:02.16" />
                    <SPLIT distance="300" swimtime="00:04:54.87" />
                    <SPLIT distance="350" swimtime="00:05:47.29" />
                    <SPLIT distance="400" swimtime="00:06:38.89" />
                    <SPLIT distance="450" swimtime="00:07:32.12" />
                    <SPLIT distance="500" swimtime="00:08:25.44" />
                    <SPLIT distance="550" swimtime="00:09:17.75" />
                    <SPLIT distance="600" swimtime="00:10:09.69" />
                    <SPLIT distance="650" swimtime="00:11:02.69" />
                    <SPLIT distance="700" swimtime="00:11:54.79" />
                    <SPLIT distance="750" swimtime="00:12:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="470" reactiontime="+91" swimtime="00:00:39.89" resultid="2259" heatid="4313" lane="7" />
                <RESULT eventid="1474" points="442" reactiontime="+102" swimtime="00:01:27.98" resultid="2260" heatid="4386" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="404" reactiontime="+103" swimtime="00:03:14.85" resultid="2261" heatid="4429" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                    <SPLIT distance="100" swimtime="00:01:33.57" />
                    <SPLIT distance="150" swimtime="00:02:25.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" clubid="3458" name="UKS ENERGETYK Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" name="Kondracki" phone="693852488" state="DOL" street="Maratońska" street2="2" zip="59-900" />
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Daszyński" birthdate="1948-11-29" gender="M" nation="POL" athleteid="3459">
              <RESULTS>
                <RESULT eventid="1112" points="224" reactiontime="+83" swimtime="00:04:28.43" resultid="3460" heatid="4292" lane="6" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.09" />
                    <SPLIT distance="100" swimtime="00:02:13.10" />
                    <SPLIT distance="150" swimtime="00:03:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="226" reactiontime="+91" swimtime="00:17:26.35" resultid="3461" heatid="4306" lane="6" entrytime="00:17:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.80" />
                    <SPLIT distance="100" swimtime="00:02:01.01" />
                    <SPLIT distance="150" swimtime="00:03:08.42" />
                    <SPLIT distance="200" swimtime="00:04:15.13" />
                    <SPLIT distance="250" swimtime="00:05:22.64" />
                    <SPLIT distance="300" swimtime="00:06:28.85" />
                    <SPLIT distance="350" swimtime="00:07:35.19" />
                    <SPLIT distance="400" swimtime="00:08:42.28" />
                    <SPLIT distance="450" swimtime="00:09:49.31" />
                    <SPLIT distance="500" swimtime="00:10:56.14" />
                    <SPLIT distance="550" swimtime="00:12:02.08" />
                    <SPLIT distance="600" swimtime="00:13:07.50" />
                    <SPLIT distance="650" swimtime="00:14:14.17" />
                    <SPLIT distance="700" swimtime="00:15:20.72" />
                    <SPLIT distance="750" swimtime="00:16:25.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="225" reactiontime="+94" swimtime="00:00:55.21" resultid="3462" heatid="4320" lane="6" entrytime="00:00:59.00" />
                <RESULT eventid="1352" points="127" reactiontime="+89" swimtime="00:05:32.43" resultid="3463" heatid="4355" lane="7" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.30" />
                    <SPLIT distance="100" swimtime="00:02:40.85" />
                    <SPLIT distance="150" swimtime="00:04:07.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="222" reactiontime="+100" swimtime="00:02:01.46" resultid="3464" heatid="4390" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="222" reactiontime="+94" swimtime="00:09:48.22" resultid="3465" heatid="4417" lane="4" entrytime="00:09:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.96" />
                    <SPLIT distance="100" swimtime="00:02:37.55" />
                    <SPLIT distance="150" swimtime="00:03:52.01" />
                    <SPLIT distance="200" swimtime="00:05:02.52" />
                    <SPLIT distance="250" swimtime="00:06:24.03" />
                    <SPLIT distance="300" swimtime="00:07:44.61" />
                    <SPLIT distance="350" swimtime="00:08:47.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="87" reactiontime="+93" swimtime="00:02:32.22" resultid="3466" heatid="4423" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="228" reactiontime="+100" swimtime="00:04:22.24" resultid="3467" heatid="4433" lane="4" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.57" />
                    <SPLIT distance="100" swimtime="00:02:12.09" />
                    <SPLIT distance="150" swimtime="00:03:20.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" clubid="3476" name="Uks Delfin Legionowo">
          <CONTACT city="LEGIONOWO" email="delfin-trener@wp.pl" internet="www.delfinlegionowo.pl" name="RAFAŁ PERL" phone="601 436 700" state="MAZ" street="KRÓLOWEJ JADWIGI 11" zip="05-120" />
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Żbikowska" birthdate="1996-01-01" gender="F" nation="POL" license="S01414100028" athleteid="3487">
              <RESULTS>
                <RESULT eventid="1059" points="574" reactiontime="+73" swimtime="00:00:30.58" resultid="3488" heatid="4271" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1094" points="504" reactiontime="+82" swimtime="00:02:56.77" resultid="3489" heatid="4290" lane="8" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:22.21" />
                    <SPLIT distance="150" swimtime="00:02:13.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="524" reactiontime="+84" swimtime="00:03:12.83" resultid="3490" heatid="4328" lane="2" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                    <SPLIT distance="100" swimtime="00:01:33.11" />
                    <SPLIT distance="150" swimtime="00:02:24.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="572" reactiontime="+81" swimtime="00:01:08.62" resultid="3491" heatid="4340" lane="0" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="596" reactiontime="+81" swimtime="00:01:23.85" resultid="3492" heatid="4365" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="505" reactiontime="+86" swimtime="00:02:36.44" resultid="3493" heatid="4398" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:14.66" />
                    <SPLIT distance="150" swimtime="00:01:57.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="613" reactiontime="+81" swimtime="00:00:37.20" resultid="3494" heatid="4441" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andzrej" lastname="Fajdasz" birthdate="1973-01-14" gender="M" nation="POL" license="101414700141" athleteid="3477">
              <RESULTS>
                <RESULT eventid="1076" points="408" reactiontime="+72" swimtime="00:00:31.74" resultid="3478" heatid="4279" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1267" points="349" reactiontime="+84" swimtime="00:00:39.24" resultid="3479" heatid="4322" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="1301" points="397" reactiontime="+80" swimtime="00:01:11.05" resultid="3480" heatid="4347" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="359" reactiontime="+87" swimtime="00:01:24.64" resultid="3481" heatid="4392" lane="7" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="339" reactiontime="+85" swimtime="00:03:08.65" resultid="3482" heatid="4435" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                    <SPLIT distance="100" swimtime="00:01:32.18" />
                    <SPLIT distance="150" swimtime="00:02:22.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Perl" birthdate="1996-06-07" gender="M" nation="POL" license="101414700068" athleteid="3483">
              <RESULTS>
                <RESULT eventid="1076" points="765" reactiontime="+67" swimtime="00:00:24.38" resultid="3484" heatid="4286" lane="4" entrytime="00:00:24.00" />
                <RESULT eventid="1406" points="680" reactiontime="+68" swimtime="00:01:08.69" resultid="3485" heatid="4371" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="727" reactiontime="+66" swimtime="00:00:30.26" resultid="3486" heatid="4449" lane="4" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2833" name="KU AZS Uniwersytetu Warszawskiego">
          <CONTACT name="Rębas Igor" phone="504784194" />
          <ATHLETES>
            <ATHLETE firstname="Rafał" lastname="Godlewski" birthdate="1996-01-01" gender="M" nation="POL" swrid="4285522" athleteid="2839">
              <RESULTS>
                <RESULT eventid="1076" points="539" reactiontime="+77" swimtime="00:00:27.40" resultid="2840" heatid="4282" lane="3" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1406" points="467" reactiontime="+79" swimtime="00:01:17.84" resultid="2841" heatid="4370" lane="5" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="398" reactiontime="+79" swimtime="00:00:32.24" resultid="2842" heatid="4382" lane="0" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1697" points="531" reactiontime="+77" swimtime="00:00:33.60" resultid="2843" heatid="4449" lane="1" entrytime="00:00:32.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rębas" birthdate="1989-01-01" gender="M" nation="POL" swrid="4251117" athleteid="2844">
              <RESULTS>
                <RESULT eventid="1301" points="708" reactiontime="+78" swimtime="00:00:55.88" resultid="2845" heatid="4350" lane="0" entrytime="00:01:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="231" reactiontime="+75" swimtime="00:02:58.68" resultid="2846" heatid="4400" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.20" />
                    <SPLIT distance="100" swimtime="00:00:56.34" />
                    <SPLIT distance="150" swimtime="00:02:08.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="2847" heatid="4418" lane="4" />
                <RESULT eventid="1629" points="688" reactiontime="+78" swimtime="00:01:00.77" resultid="2848" heatid="4426" lane="4" entrytime="00:01:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Kister" birthdate="1989-01-01" gender="M" nation="POL" swrid="4992691" athleteid="2849">
              <RESULTS>
                <RESULT eventid="1250" status="DNS" swimtime="00:00:00.00" resultid="2850" heatid="4333" lane="8" entrytime="00:02:59.00" entrycourse="LCM" />
                <RESULT eventid="1352" status="DNS" swimtime="00:00:00.00" resultid="2851" heatid="4357" lane="1" entrytime="00:02:44.00" entrycourse="LCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="2852" heatid="4370" lane="8" entrytime="00:01:18.50" entrycourse="LCM" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="2853" heatid="4382" lane="8" entrytime="00:00:29.90" entrycourse="LCM" />
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="2854" heatid="4425" lane="4" entrytime="00:01:09.90" entrycourse="LCM" />
                <RESULT eventid="1697" status="DNS" swimtime="00:00:00.00" resultid="2855" heatid="4447" lane="4" entrytime="00:00:34.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Micorek" birthdate="1993-01-01" gender="M" nation="POL" swrid="4086676" athleteid="2834">
              <RESULTS>
                <RESULT eventid="1076" points="617" reactiontime="+72" swimtime="00:00:26.20" resultid="2835" heatid="4284" lane="7" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="1267" status="DNS" swimtime="00:00:00.00" resultid="2836" heatid="4325" lane="6" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1301" reactiontime="+69" status="DNF" swimtime="00:00:00.00" resultid="2837" heatid="4341" lane="6" entrytime="00:00:54.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="635" reactiontime="+73" swimtime="00:00:27.58" resultid="2838" heatid="4383" lane="5" entrytime="00:00:28.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3673" name="3Waters">
          <ATHLETES>
            <ATHLETE firstname="Sonia" lastname="BORKOWSKA" birthdate="1975-01-01" gender="F" nation="POL" athleteid="3674">
              <RESULTS>
                <RESULT eventid="1059" points="542" reactiontime="+51" swimtime="00:00:32.61" resultid="3675" heatid="4270" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1440" points="375" reactiontime="+81" swimtime="00:00:39.38" resultid="3676" heatid="4373" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1215" points="370" reactiontime="+84" swimtime="00:00:43.22" resultid="3677" heatid="4315" lane="0" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01813" nation="POL" region="13" clubid="2518" name="SWIMLAND Olsztyn">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Wójtowicz" birthdate="1995-02-20" gender="F" nation="POL" license="101813600026" swrid="4265548" athleteid="2519">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1059" points="879" reactiontime="+64" swimtime="00:00:26.54" resultid="2520" heatid="4272" lane="4" entrytime="00:00:26.40" entrycourse="SCM" />
                <RESULT comment="Rekord Polski w kat.masters, Wynik lepszy od Rekordu Europy w kat. masters" eventid="1215" points="871" reactiontime="+65" swimtime="00:00:29.73" resultid="2521" heatid="4316" lane="4" entrytime="00:00:30.09" entrycourse="LCM" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1440" points="780" reactiontime="+54" swimtime="00:00:28.59" resultid="2522" heatid="4375" lane="4" entrytime="00:00:28.29" entrycourse="LCM" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1474" points="844" reactiontime="+69" swimtime="00:01:05.18" resultid="2523" heatid="4388" lane="4" entrytime="00:01:01.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="2524" heatid="4421" lane="4" entrytime="00:01:02.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02016" nation="POL" region="16" clubid="1983" name="Koszalińskie TKKF">
          <CONTACT email="roman.pieslak@gmail.com" name="Roman" phone="600227112" street="Pieślak" />
          <ATHLETES>
            <ATHLETE firstname="Izabela" lastname="Kijanka" birthdate="1982-08-02" gender="F" nation="POL" athleteid="4219">
              <RESULTS>
                <RESULT eventid="1094" points="430" reactiontime="+79" swimtime="00:03:12.19" resultid="4220" heatid="4289" lane="9" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:01:34.34" />
                    <SPLIT distance="150" swimtime="00:02:29.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="324" reactiontime="+95" swimtime="00:13:04.93" resultid="4221" heatid="4300" lane="0" entrytime="00:13:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:21.54" />
                    <SPLIT distance="100" swimtime="00:01:31.39" />
                    <SPLIT distance="150" swimtime="00:04:02.43" />
                    <SPLIT distance="200" swimtime="00:03:11.86" />
                    <SPLIT distance="250" swimtime="00:05:45.15" />
                    <SPLIT distance="300" swimtime="00:04:53.56" />
                    <SPLIT distance="350" swimtime="00:10:44.31" />
                    <SPLIT distance="400" swimtime="00:06:35.25" />
                    <SPLIT distance="500" swimtime="00:08:15.62" />
                    <SPLIT distance="600" swimtime="00:09:55.82" />
                    <SPLIT distance="700" swimtime="00:11:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="450" reactiontime="+91" swimtime="00:03:26.83" resultid="4222" heatid="4328" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                    <SPLIT distance="100" swimtime="00:01:37.78" />
                    <SPLIT distance="150" swimtime="00:02:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="402" reactiontime="+92" swimtime="00:01:18.67" resultid="4223" heatid="4339" lane="7" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="414" reactiontime="+84" swimtime="00:00:38.05" resultid="4224" heatid="4373" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1508" points="382" reactiontime="+85" swimtime="00:02:58.15" resultid="4225" heatid="4397" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:24.07" />
                    <SPLIT distance="150" swimtime="00:02:11.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="443" reactiontime="+87" swimtime="00:00:42.59" resultid="4226" heatid="4441" lane="9" entrytime="00:00:43.00" />
                <RESULT eventid="1731" points="306" reactiontime="+90" swimtime="00:06:30.25" resultid="4227" heatid="4453" lane="2" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                    <SPLIT distance="100" swimtime="00:01:30.14" />
                    <SPLIT distance="150" swimtime="00:02:18.97" />
                    <SPLIT distance="200" swimtime="00:03:08.84" />
                    <SPLIT distance="250" swimtime="00:03:58.98" />
                    <SPLIT distance="300" swimtime="00:04:49.84" />
                    <SPLIT distance="350" swimtime="00:05:41.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Pieślak" birthdate="1979-02-28" gender="M" nation="POL" athleteid="4202">
              <RESULTS>
                <RESULT eventid="1076" points="492" reactiontime="+75" swimtime="00:00:29.46" resultid="4203" heatid="4280" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1163" points="449" reactiontime="+76" swimtime="00:11:13.72" resultid="4204" heatid="4304" lane="2" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:53.22" />
                    <SPLIT distance="200" swimtime="00:02:33.68" />
                    <SPLIT distance="250" swimtime="00:03:14.52" />
                    <SPLIT distance="300" swimtime="00:03:55.86" />
                    <SPLIT distance="350" swimtime="00:04:37.43" />
                    <SPLIT distance="400" swimtime="00:05:19.82" />
                    <SPLIT distance="450" swimtime="00:06:02.61" />
                    <SPLIT distance="500" swimtime="00:06:46.29" />
                    <SPLIT distance="550" swimtime="00:07:30.18" />
                    <SPLIT distance="600" swimtime="00:08:14.26" />
                    <SPLIT distance="650" swimtime="00:08:58.60" />
                    <SPLIT distance="700" swimtime="00:09:43.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="456" reactiontime="+75" swimtime="00:02:59.98" resultid="4205" heatid="4332" lane="6" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="100" swimtime="00:01:25.69" />
                    <SPLIT distance="150" swimtime="00:02:12.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="467" reactiontime="+71" swimtime="00:01:22.00" resultid="4206" heatid="4369" lane="3" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="464" reactiontime="+71" swimtime="00:02:26.78" resultid="4207" heatid="4404" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:08.20" />
                    <SPLIT distance="150" swimtime="00:01:46.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="477" reactiontime="+74" swimtime="00:00:36.90" resultid="4208" heatid="4446" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1748" points="477" reactiontime="+77" swimtime="00:05:15.82" resultid="4209" heatid="4459" lane="3" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:14.91" />
                    <SPLIT distance="150" swimtime="00:01:54.58" />
                    <SPLIT distance="200" swimtime="00:02:35.39" />
                    <SPLIT distance="250" swimtime="00:03:16.56" />
                    <SPLIT distance="300" swimtime="00:03:57.29" />
                    <SPLIT distance="350" swimtime="00:04:37.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Mamrot" birthdate="1972-12-10" gender="M" nation="POL" athleteid="4195">
              <RESULTS>
                <RESULT eventid="1076" points="400" reactiontime="+83" swimtime="00:00:32.67" resultid="4196" heatid="4279" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1112" points="351" reactiontime="+84" swimtime="00:03:05.91" resultid="4197" heatid="4294" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="100" swimtime="00:01:27.65" />
                    <SPLIT distance="150" swimtime="00:02:21.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="349" reactiontime="+91" swimtime="00:03:29.70" resultid="4198" heatid="4332" lane="9" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.76" />
                    <SPLIT distance="100" swimtime="00:01:36.90" />
                    <SPLIT distance="150" swimtime="00:02:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="365" reactiontime="+85" swimtime="00:01:32.95" resultid="4199" heatid="4369" lane="0" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="396" reactiontime="+82" swimtime="00:00:41.07" resultid="4200" heatid="4445" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1748" points="339" reactiontime="+81" swimtime="00:06:06.87" resultid="4201" heatid="4460" lane="7" entrytime="00:06:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                    <SPLIT distance="100" swimtime="00:01:24.82" />
                    <SPLIT distance="150" swimtime="00:02:11.78" />
                    <SPLIT distance="200" swimtime="00:02:59.30" />
                    <SPLIT distance="250" swimtime="00:03:47.97" />
                    <SPLIT distance="300" swimtime="00:04:36.17" />
                    <SPLIT distance="350" swimtime="00:05:23.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Winiarczyk" birthdate="1972-01-23" gender="M" nation="POL" athleteid="4210">
              <RESULTS>
                <RESULT eventid="1076" points="608" reactiontime="+77" swimtime="00:00:28.42" resultid="4211" heatid="4280" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1163" points="553" reactiontime="+70" swimtime="00:10:51.83" resultid="4212" heatid="4304" lane="6" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="150" swimtime="00:01:53.35" />
                    <SPLIT distance="200" swimtime="00:02:34.03" />
                    <SPLIT distance="250" swimtime="00:03:14.76" />
                    <SPLIT distance="300" swimtime="00:03:55.90" />
                    <SPLIT distance="350" swimtime="00:04:37.93" />
                    <SPLIT distance="400" swimtime="00:05:19.76" />
                    <SPLIT distance="450" swimtime="00:06:01.96" />
                    <SPLIT distance="500" swimtime="00:06:44.29" />
                    <SPLIT distance="550" swimtime="00:07:26.36" />
                    <SPLIT distance="600" swimtime="00:08:09.23" />
                    <SPLIT distance="650" swimtime="00:08:52.29" />
                    <SPLIT distance="700" swimtime="00:09:33.75" />
                    <SPLIT distance="750" swimtime="00:10:15.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="509" reactiontime="+74" swimtime="00:00:35.79" resultid="4213" heatid="4322" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1301" points="628" reactiontime="+64" swimtime="00:01:03.23" resultid="4214" heatid="4347" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="579" reactiontime="+64" swimtime="00:02:22.32" resultid="4215" heatid="4405" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:09.37" />
                    <SPLIT distance="150" swimtime="00:01:47.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="418" reactiontime="+72" swimtime="00:06:22.02" resultid="4216" heatid="4415" lane="8" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:01:27.56" />
                    <SPLIT distance="150" swimtime="00:02:20.29" />
                    <SPLIT distance="200" swimtime="00:03:10.40" />
                    <SPLIT distance="250" swimtime="00:04:03.00" />
                    <SPLIT distance="300" swimtime="00:04:57.32" />
                    <SPLIT distance="350" swimtime="00:05:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="454" reactiontime="+62" swimtime="00:02:55.04" resultid="4217" heatid="4435" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:25.72" />
                    <SPLIT distance="150" swimtime="00:02:12.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="553" reactiontime="+66" swimtime="00:05:11.74" resultid="4218" heatid="4459" lane="5" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:13.25" />
                    <SPLIT distance="150" swimtime="00:01:53.48" />
                    <SPLIT distance="200" swimtime="00:02:34.48" />
                    <SPLIT distance="250" swimtime="00:03:15.38" />
                    <SPLIT distance="300" swimtime="00:03:56.21" />
                    <SPLIT distance="350" swimtime="00:04:36.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kielar" birthdate="1974-01-21" gender="M" nation="POL" athleteid="4228">
              <RESULTS>
                <RESULT eventid="1076" points="590" reactiontime="+88" swimtime="00:00:28.08" resultid="4229" heatid="4283" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="1112" points="552" reactiontime="+93" swimtime="00:02:38.58" resultid="4230" heatid="4295" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:14.04" />
                    <SPLIT distance="150" swimtime="00:02:02.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="498" reactiontime="+78" swimtime="00:00:34.85" resultid="4231" heatid="4324" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="4232" heatid="4349" lane="8" entrytime="00:01:03.00" />
                <RESULT eventid="1457" points="667" reactiontime="+99" swimtime="00:00:28.89" resultid="4233" heatid="4383" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1491" points="507" reactiontime="+79" swimtime="00:01:15.43" resultid="4234" heatid="4393" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="631" reactiontime="+79" swimtime="00:01:06.27" resultid="4235" heatid="4425" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="529" reactiontime="+84" swimtime="00:00:36.13" resultid="4236" heatid="4445" lane="3" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1386" points="494" swimtime="00:02:13.41" resultid="4237" heatid="4493" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:12.40" />
                    <SPLIT distance="150" swimtime="00:01:41.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4210" number="1" />
                    <RELAYPOSITION athleteid="4202" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4228" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4195" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1559" points="531" reactiontime="+85" swimtime="00:01:57.22" resultid="4238" heatid="4497" lane="8" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                    <SPLIT distance="100" swimtime="00:00:59.62" />
                    <SPLIT distance="150" swimtime="00:01:29.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4228" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="4195" number="2" />
                    <RELAYPOSITION athleteid="4202" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4210" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="2270" name="MKS ,,Astoria&apos;&apos; Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Bartosz" lastname="Ciężki" birthdate="1994-09-30" gender="M" nation="POL" license="102202700137" swrid="4289450" athleteid="2271">
              <RESULTS>
                <RESULT eventid="1076" points="626" reactiontime="+77" swimtime="00:00:26.07" resultid="2272" heatid="4286" lane="8" entrytime="00:00:25.89" entrycourse="LCM" />
                <RESULT eventid="1163" points="596" reactiontime="+88" swimtime="00:09:59.73" resultid="2273" heatid="4306" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="100" swimtime="00:01:02.97" />
                    <SPLIT distance="150" swimtime="00:01:38.25" />
                    <SPLIT distance="200" swimtime="00:02:14.59" />
                    <SPLIT distance="250" swimtime="00:02:51.83" />
                    <SPLIT distance="300" swimtime="00:03:30.05" />
                    <SPLIT distance="350" swimtime="00:04:07.94" />
                    <SPLIT distance="400" swimtime="00:04:46.64" />
                    <SPLIT distance="450" swimtime="00:05:25.50" />
                    <SPLIT distance="500" swimtime="00:06:05.06" />
                    <SPLIT distance="550" swimtime="00:06:44.46" />
                    <SPLIT distance="600" swimtime="00:07:24.60" />
                    <SPLIT distance="650" swimtime="00:08:04.72" />
                    <SPLIT distance="700" swimtime="00:08:44.84" />
                    <SPLIT distance="750" swimtime="00:09:23.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="430" reactiontime="+87" swimtime="00:02:40.29" resultid="2274" heatid="4357" lane="2" entrytime="00:02:33.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="150" swimtime="00:01:52.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="643" reactiontime="+82" swimtime="00:02:08.31" resultid="2275" heatid="4407" lane="6" entrytime="00:02:03.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                    <SPLIT distance="100" swimtime="00:00:59.55" />
                    <SPLIT distance="150" swimtime="00:01:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="537" reactiontime="+72" swimtime="00:02:31.00" resultid="2276" heatid="4432" lane="3" entrytime="00:02:35.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:52.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Krasicki" birthdate="1995-02-17" gender="M" nation="POL" license="102202700140" swrid="4169744" athleteid="2282">
              <RESULTS>
                <RESULT eventid="1457" points="603" reactiontime="+74" swimtime="00:00:28.06" resultid="2283" heatid="4377" lane="1" />
                <RESULT eventid="1525" points="623" reactiontime="+71" swimtime="00:02:09.67" resultid="2284" heatid="4406" lane="3" entrytime="00:02:10.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                    <SPLIT distance="100" swimtime="00:01:01.73" />
                    <SPLIT distance="150" swimtime="00:01:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="616" reactiontime="+75" swimtime="00:04:43.19" resultid="2285" heatid="4463" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="100" swimtime="00:01:04.44" />
                    <SPLIT distance="150" swimtime="00:01:39.80" />
                    <SPLIT distance="200" swimtime="00:02:16.51" />
                    <SPLIT distance="250" swimtime="00:02:53.37" />
                    <SPLIT distance="300" swimtime="00:03:30.87" />
                    <SPLIT distance="350" swimtime="00:04:07.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" license="102202700126" swrid="5471726" athleteid="2277">
              <RESULTS>
                <RESULT eventid="1267" points="164" reactiontime="+96" swimtime="00:00:52.19" resultid="2278" heatid="4320" lane="5" entrytime="00:00:53.09" entrycourse="SCM" />
                <RESULT eventid="1491" points="141" reactiontime="+92" swimtime="00:01:58.27" resultid="2279" heatid="4390" lane="4" entrytime="00:01:55.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" status="DNS" swimtime="00:00:00.00" resultid="2280" heatid="4433" lane="9" />
                <RESULT eventid="1697" points="273" reactiontime="+80" swimtime="00:00:46.50" resultid="2281" heatid="4443" lane="4" entrytime="00:00:52.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="AUS" clubid="5115" name="Tomatoes Swim Club">
          <ATHLETES>
            <ATHLETE firstname="MACIEJ" lastname="SLUGOCKI" birthdate="1952-01-01" gender="M" nation="AUS" athleteid="3913">
              <RESULTS>
                <RESULT eventid="1112" points="657" reactiontime="+87" swimtime="00:03:07.40" resultid="3914" heatid="4294" lane="7" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                    <SPLIT distance="100" swimtime="00:01:30.57" />
                    <SPLIT distance="150" swimtime="00:02:24.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1197" reactiontime="+92" status="DNF" swimtime="00:00:00.00" resultid="3915" heatid="4310" lane="5" entrytime="00:22:35.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                    <SPLIT distance="150" swimtime="00:02:08.03" />
                    <SPLIT distance="200" swimtime="00:02:51.12" />
                    <SPLIT distance="250" swimtime="00:03:34.60" />
                    <SPLIT distance="300" swimtime="00:04:17.52" />
                    <SPLIT distance="350" swimtime="00:05:00.28" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1267" points="551" reactiontime="+105" swimtime="00:00:40.97" resultid="3916" heatid="4321" lane="3" entrytime="00:00:41.80" />
                <RESULT eventid="1250" points="605" reactiontime="+100" swimtime="00:03:38.53" resultid="3917" heatid="4331" lane="3" entrytime="00:03:48.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.16" />
                    <SPLIT distance="100" swimtime="00:01:48.64" />
                    <SPLIT distance="150" swimtime="00:02:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="635" reactiontime="+86" swimtime="00:01:35.40" resultid="3918" heatid="4368" lane="7" entrytime="00:01:39.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="503" reactiontime="+91" swimtime="00:00:37.70" resultid="3919" heatid="4379" lane="7" entrytime="00:00:43.63" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1491" points="486" reactiontime="+100" status="EXH" swimtime="00:01:33.47" resultid="3920" heatid="4391" lane="2" entrytime="00:01:36.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1629" points="387" reactiontime="+96" swimtime="00:01:32.48" resultid="3921" heatid="4423" lane="3" entrytime="00:01:48.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="623" reactiontime="+95" swimtime="00:00:42.40" resultid="3922" heatid="4444" lane="1" entrytime="00:00:48.73" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3740" name="Swim Club Masters Ślęza">
          <ATHLETES>
            <ATHLETE firstname="JOANNA" lastname="CHOJCAN" birthdate="1986-01-01" gender="F" nation="POL" athleteid="3741">
              <RESULTS>
                <RESULT eventid="1059" points="522" reactiontime="+79" swimtime="00:00:32.27" resultid="3742" heatid="4271" lane="8" entrytime="00:00:32.50" />
                <RESULT eventid="1094" points="508" reactiontime="+78" swimtime="00:02:57.35" resultid="3743" heatid="4289" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:15.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="470" reactiontime="+68" swimtime="00:00:36.83" resultid="3744" heatid="4315" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1335" points="366" reactiontime="+80" swimtime="00:03:15.99" resultid="3745" heatid="4354" lane="1" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:25.61" />
                    <SPLIT distance="150" swimtime="00:02:17.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="466" reactiontime="+70" swimtime="00:01:19.63" resultid="3746" heatid="4388" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1576" points="498" reactiontime="+74" swimtime="00:06:17.91" resultid="3747" heatid="4412" lane="7" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:13.44" />
                    <SPLIT distance="200" swimtime="00:03:00.41" />
                    <SPLIT distance="250" swimtime="00:03:54.26" />
                    <SPLIT distance="300" swimtime="00:04:48.92" />
                    <SPLIT distance="350" swimtime="00:05:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="473" reactiontime="+78" swimtime="00:01:20.16" resultid="3748" heatid="4420" lane="5" entrytime="00:01:27.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="488" reactiontime="+83" swimtime="00:02:55.52" resultid="3749" heatid="4431" lane="1" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:23.92" />
                    <SPLIT distance="150" swimtime="00:02:10.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="14814" nation="POL" region="14" clubid="2478" name="Stowarzyszenie Pływackie Legia Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Bogdan" lastname="Dubiński" birthdate="1953-05-05" gender="M" nation="POL" license="514814700003" swrid="4992696" athleteid="2479">
              <RESULTS>
                <RESULT eventid="1076" points="408" reactiontime="+86" swimtime="00:00:35.35" resultid="2480" heatid="4277" lane="6" entrytime="00:00:36.58" entrycourse="LCM" />
                <RESULT eventid="1163" points="357" reactiontime="+85" swimtime="00:14:21.36" resultid="2481" heatid="4306" lane="5" entrytime="00:15:37.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                    <SPLIT distance="100" swimtime="00:01:32.18" />
                    <SPLIT distance="150" swimtime="00:02:25.37" />
                    <SPLIT distance="200" swimtime="00:03:19.27" />
                    <SPLIT distance="250" swimtime="00:04:15.07" />
                    <SPLIT distance="300" swimtime="00:05:09.38" />
                    <SPLIT distance="350" swimtime="00:06:05.52" />
                    <SPLIT distance="400" swimtime="00:07:02.39" />
                    <SPLIT distance="450" swimtime="00:07:59.14" />
                    <SPLIT distance="500" swimtime="00:08:54.89" />
                    <SPLIT distance="550" swimtime="00:09:50.21" />
                    <SPLIT distance="600" swimtime="00:10:45.65" />
                    <SPLIT distance="650" swimtime="00:11:40.57" />
                    <SPLIT distance="700" swimtime="00:12:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="365" reactiontime="+98" swimtime="00:00:43.31" resultid="2482" heatid="4321" lane="2" entrytime="00:00:43.68" entrycourse="LCM" />
                <RESULT eventid="1301" points="383" reactiontime="+94" swimtime="00:01:21.90" resultid="2483" heatid="4341" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="350" reactiontime="+92" swimtime="00:01:39.01" resultid="2484" heatid="4389" lane="6" />
                <RESULT eventid="1525" points="325" reactiontime="+94" swimtime="00:03:08.21" resultid="2485" heatid="4401" lane="5" entrytime="00:03:25.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                    <SPLIT distance="100" swimtime="00:01:30.40" />
                    <SPLIT distance="150" swimtime="00:02:21.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="187" reactiontime="+92" swimtime="00:01:55.12" resultid="2486" heatid="4422" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="311" reactiontime="+97" swimtime="00:06:50.08" resultid="2487" heatid="4461" lane="7" entrytime="00:07:25.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                    <SPLIT distance="100" swimtime="00:01:33.43" />
                    <SPLIT distance="150" swimtime="00:02:27.33" />
                    <SPLIT distance="200" swimtime="00:03:21.37" />
                    <SPLIT distance="250" swimtime="00:04:15.27" />
                    <SPLIT distance="350" swimtime="00:06:02.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3304" name="Motyl Master">
          <CONTACT city="Stalowa Wola" email="elzbietalorkowska@gmail.com" name="Chmielewski Andrzej" phone="15-84473-38" state="POD" street="Hutnicza 165" zip="37-450" />
          <ATHLETES>
            <ATHLETE firstname="Arkadiusz" lastname="Berwecki" birthdate="1973-01-14" gender="M" nation="POL" athleteid="3346">
              <RESULTS>
                <RESULT eventid="1076" points="643" reactiontime="+71" swimtime="00:00:27.29" resultid="3347" heatid="4285" lane="7" entrytime="00:00:26.49" />
                <RESULT eventid="1112" points="698" reactiontime="+80" swimtime="00:02:26.62" resultid="3348" heatid="4297" lane="8" entrytime="00:02:24.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="100" swimtime="00:01:09.05" />
                    <SPLIT distance="150" swimtime="00:01:50.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="713" reactiontime="+77" swimtime="00:00:58.48" resultid="3349" heatid="4351" lane="8" entrytime="00:00:58.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="600" reactiontime="+82" swimtime="00:01:16.78" resultid="3350" heatid="4371" lane="9" entrytime="00:01:14.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="698" reactiontime="+71" swimtime="00:00:28.46" resultid="3351" heatid="4383" lane="4" entrytime="00:00:27.99" />
                <RESULT eventid="1629" points="738" reactiontime="+78" swimtime="00:01:02.92" resultid="3352" heatid="4427" lane="8" entrytime="00:01:01.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="613" reactiontime="+78" swimtime="00:00:34.39" resultid="3353" heatid="4448" lane="7" entrytime="00:00:33.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Pawłowski" birthdate="1977-06-26" gender="M" nation="POL" athleteid="3314">
              <RESULTS>
                <RESULT eventid="1112" points="430" reactiontime="+86" swimtime="00:02:52.37" resultid="3315" heatid="4294" lane="3" entrytime="00:03:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:02:11.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="394" reactiontime="+83" swimtime="00:11:50.13" resultid="3316" heatid="4305" lane="3" entrytime="00:12:05.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                    <SPLIT distance="150" swimtime="00:02:02.41" />
                    <SPLIT distance="200" swimtime="00:02:46.60" />
                    <SPLIT distance="250" swimtime="00:03:30.96" />
                    <SPLIT distance="300" swimtime="00:04:16.08" />
                    <SPLIT distance="350" swimtime="00:05:00.47" />
                    <SPLIT distance="400" swimtime="00:05:46.24" />
                    <SPLIT distance="450" swimtime="00:06:31.53" />
                    <SPLIT distance="500" swimtime="00:07:17.45" />
                    <SPLIT distance="550" swimtime="00:08:02.82" />
                    <SPLIT distance="600" swimtime="00:08:48.39" />
                    <SPLIT distance="650" swimtime="00:09:33.64" />
                    <SPLIT distance="700" swimtime="00:10:19.21" />
                    <SPLIT distance="750" swimtime="00:11:04.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="519" reactiontime="+73" swimtime="00:00:34.36" resultid="3317" heatid="4322" lane="4" entrytime="00:00:36.80" />
                <RESULT eventid="1250" points="366" reactiontime="+86" swimtime="00:03:14.86" resultid="3318" heatid="4332" lane="2" entrytime="00:03:08.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:33.72" />
                    <SPLIT distance="150" swimtime="00:02:24.89" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O3" eventid="1491" reactiontime="+79" status="DSQ" swimtime="00:01:16.68" resultid="3319" heatid="4393" lane="9" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="3320" heatid="4415" lane="7" entrytime="00:06:12.70" />
                <RESULT eventid="1663" points="404" reactiontime="+97" swimtime="00:02:58.03" resultid="3321" heatid="4436" lane="8" entrytime="00:02:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:24.67" />
                    <SPLIT distance="150" swimtime="00:02:11.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="413" reactiontime="+82" swimtime="00:00:39.24" resultid="3322" heatid="4446" lane="4" entrytime="00:00:36.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Jarzyna" birthdate="1949-08-09" gender="M" nation="POL" athleteid="3338">
              <RESULTS>
                <RESULT eventid="1112" points="356" reactiontime="+91" swimtime="00:03:49.97" resultid="3339" heatid="4293" lane="0" entrytime="00:03:55.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.77" />
                    <SPLIT distance="100" swimtime="00:01:53.17" />
                    <SPLIT distance="150" swimtime="00:03:02.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="366" reactiontime="+100" swimtime="00:00:46.95" resultid="3340" heatid="4320" lane="3" entrytime="00:00:58.80" />
                <RESULT eventid="1250" points="427" reactiontime="+113" swimtime="00:04:05.46" resultid="3341" heatid="4331" lane="8" entrytime="00:04:01.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.68" />
                    <SPLIT distance="100" swimtime="00:01:57.70" />
                    <SPLIT distance="150" swimtime="00:03:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="402" reactiontime="+115" swimtime="00:01:51.10" resultid="3342" heatid="4367" lane="3" entrytime="00:01:59.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="358" reactiontime="+87" swimtime="00:01:43.50" resultid="3343" heatid="4390" lane="5" entrytime="00:01:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="359" reactiontime="+108" swimtime="00:03:45.46" resultid="3344" heatid="4434" lane="9" entrytime="00:03:58.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.37" />
                    <SPLIT distance="100" swimtime="00:01:52.67" />
                    <SPLIT distance="150" swimtime="00:02:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="426" reactiontime="+98" swimtime="00:00:48.12" resultid="3345" heatid="4443" lane="3" entrytime="00:00:59.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Baran" birthdate="1975-03-19" gender="M" nation="POL" athleteid="3332">
              <RESULTS>
                <RESULT eventid="1076" points="558" reactiontime="+89" swimtime="00:00:28.60" resultid="3333" heatid="4284" lane="9" entrytime="00:00:27.20" />
                <RESULT eventid="1267" points="683" reactiontime="+82" swimtime="00:00:31.36" resultid="3334" heatid="4324" lane="2" entrytime="00:00:32.10" />
                <RESULT eventid="1352" points="379" reactiontime="+93" swimtime="00:02:55.35" resultid="3335" heatid="4356" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                    <SPLIT distance="100" swimtime="00:01:24.91" />
                    <SPLIT distance="150" swimtime="00:02:13.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="644" reactiontime="+81" swimtime="00:01:09.62" resultid="3336" heatid="4394" lane="2" entrytime="00:01:08.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="567" reactiontime="+80" swimtime="00:02:38.91" resultid="3337" heatid="4436" lane="5" entrytime="00:02:38.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:15.99" />
                    <SPLIT distance="150" swimtime="00:01:58.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Lorkowski" birthdate="1960-02-27" gender="M" nation="POL" athleteid="3305">
              <RESULTS>
                <RESULT eventid="1076" points="505" reactiontime="+80" swimtime="00:00:31.68" resultid="3306" heatid="4278" lane="3" entrytime="00:00:32.80" />
                <RESULT eventid="1112" points="489" reactiontime="+85" swimtime="00:03:00.26" resultid="3307" heatid="4294" lane="2" entrytime="00:03:06.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:24.08" />
                    <SPLIT distance="150" swimtime="00:02:19.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="531" reactiontime="+94" swimtime="00:01:11.38" resultid="3308" heatid="4346" lane="2" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="331" reactiontime="+88" swimtime="00:03:27.57" resultid="3309" heatid="4356" lane="8" entrytime="00:03:35.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:32.80" />
                    <SPLIT distance="150" swimtime="00:02:28.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="481" reactiontime="+95" swimtime="00:02:43.01" resultid="3310" heatid="4403" lane="8" entrytime="00:02:45.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:01:18.73" />
                    <SPLIT distance="150" swimtime="00:02:01.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="479" reactiontime="+99" swimtime="00:06:33.82" resultid="3311" heatid="4415" lane="9" entrytime="00:06:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:01:32.44" />
                    <SPLIT distance="150" swimtime="00:02:23.26" />
                    <SPLIT distance="200" swimtime="00:03:12.88" />
                    <SPLIT distance="250" swimtime="00:04:10.27" />
                    <SPLIT distance="300" swimtime="00:05:07.89" />
                    <SPLIT distance="350" swimtime="00:05:52.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="489" reactiontime="+100" swimtime="00:03:05.48" resultid="3312" heatid="4434" lane="5" entrytime="00:03:15.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                    <SPLIT distance="100" swimtime="00:01:30.39" />
                    <SPLIT distance="150" swimtime="00:02:19.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="479" reactiontime="+90" swimtime="00:05:53.81" resultid="3313" heatid="4460" lane="6" entrytime="00:05:59.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:21.95" />
                    <SPLIT distance="150" swimtime="00:02:06.55" />
                    <SPLIT distance="200" swimtime="00:02:52.80" />
                    <SPLIT distance="250" swimtime="00:03:39.05" />
                    <SPLIT distance="300" swimtime="00:04:25.92" />
                    <SPLIT distance="350" swimtime="00:05:11.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Petecka" birthdate="1967-04-17" gender="F" nation="POL" athleteid="3323">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="3324" heatid="4269" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1094" points="440" reactiontime="+87" swimtime="00:03:19.14" resultid="3325" heatid="4289" lane="8" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:37.70" />
                    <SPLIT distance="150" swimtime="00:02:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="513" reactiontime="+85" swimtime="00:03:43.44" resultid="3326" heatid="4327" lane="6" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.37" />
                    <SPLIT distance="100" swimtime="00:01:49.00" />
                    <SPLIT distance="150" swimtime="00:02:47.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" status="DNS" swimtime="00:00:00.00" resultid="3327" heatid="4338" lane="0" entrytime="00:01:23.00" />
                <RESULT eventid="1404" points="416" reactiontime="+90" swimtime="00:01:47.05" resultid="3328" heatid="4364" lane="7" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="387" reactiontime="+92" swimtime="00:00:41.89" resultid="3329" heatid="4373" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1611" points="340" reactiontime="+87" swimtime="00:01:39.55" resultid="3330" heatid="4420" lane="1" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="395" reactiontime="+81" swimtime="00:00:48.99" resultid="3331" heatid="4440" lane="1" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1386" points="621" reactiontime="+87" swimtime="00:02:09.91" resultid="3354" heatid="4493" lane="9" entrytime="00:02:12.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:38.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3332" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3314" number="2" />
                    <RELAYPOSITION athleteid="3346" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3305" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" points="584" reactiontime="+90" swimtime="00:01:57.54" resultid="3355" heatid="4496" lane="3" entrytime="00:02:01.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:01.24" />
                    <SPLIT distance="150" swimtime="00:01:30.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3332" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="3305" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="3314" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="3346" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02805" nation="POL" region="05" clubid="2295" name="MUKS Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ANDRZEJA 14" zip="95-100" />
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Sypniewski" birthdate="1957-02-01" gender="M" nation="POL" license="102805700035" swrid="5373999" athleteid="2370">
              <RESULTS>
                <RESULT eventid="1076" points="481" reactiontime="+70" swimtime="00:00:33.45" resultid="2371" heatid="4274" lane="1" />
                <RESULT eventid="1112" points="350" reactiontime="+68" swimtime="00:03:26.03" resultid="2372" heatid="4291" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                    <SPLIT distance="100" swimtime="00:01:35.19" />
                    <SPLIT distance="150" swimtime="00:02:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="432" reactiontime="+72" swimtime="00:00:40.93" resultid="2373" heatid="4318" lane="2" />
                <RESULT eventid="1250" points="377" reactiontime="+72" swimtime="00:03:43.59" resultid="2374" heatid="4329" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.90" />
                    <SPLIT distance="100" swimtime="00:01:45.42" />
                    <SPLIT distance="150" swimtime="00:02:45.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="402" reactiontime="+76" swimtime="00:01:41.27" resultid="2375" heatid="4366" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="414" reactiontime="+79" swimtime="00:00:38.08" resultid="2376" heatid="4378" lane="8" />
                <RESULT eventid="1629" points="221" reactiontime="+79" swimtime="00:01:48.95" resultid="2377" heatid="4423" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="454" reactiontime="+78" swimtime="00:00:43.32" resultid="2378" heatid="4442" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Gajda" birthdate="1978-02-23" gender="M" nation="POL" license="502805700059" swrid="5272788" athleteid="2397">
              <RESULTS>
                <RESULT eventid="1076" points="367" reactiontime="+97" swimtime="00:00:32.47" resultid="2398" heatid="4280" lane="8" entrytime="00:00:30.94" entrycourse="LCM" />
                <RESULT eventid="1267" points="416" reactiontime="+78" swimtime="00:00:36.34" resultid="2399" heatid="4323" lane="9" entrytime="00:00:36.72" entrycourse="LCM" />
                <RESULT eventid="1406" points="285" reactiontime="+89" swimtime="00:01:36.59" resultid="2400" heatid="4368" lane="5" entrytime="00:01:34.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="314" reactiontime="+80" swimtime="00:01:26.03" resultid="2401" heatid="4392" lane="8" entrytime="00:01:24.08" entrycourse="LCM" />
                <RESULT eventid="1697" points="343" reactiontime="+89" swimtime="00:00:41.19" resultid="2402" heatid="4445" lane="6" entrytime="00:00:39.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Waldemar" lastname="Jagiełło" birthdate="1979-03-01" gender="M" nation="POL" license="502805700042" swrid="4541616" athleteid="2346">
              <RESULTS>
                <RESULT eventid="1076" points="632" reactiontime="+84" swimtime="00:00:27.09" resultid="2347" heatid="4275" lane="8" />
                <RESULT eventid="1112" status="DNS" swimtime="00:00:00.00" resultid="2348" heatid="4291" lane="2" />
                <RESULT eventid="1250" status="DNS" swimtime="00:00:00.00" resultid="2349" heatid="4330" lane="0" />
                <RESULT eventid="1301" points="576" reactiontime="+81" swimtime="00:01:01.54" resultid="2350" heatid="4342" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="602" reactiontime="+79" swimtime="00:01:15.33" resultid="2351" heatid="4366" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="481" reactiontime="+86" swimtime="00:02:25.01" resultid="2352" heatid="4401" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="150" swimtime="00:01:48.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="661" reactiontime="+79" swimtime="00:00:33.11" resultid="2353" heatid="4442" lane="3" />
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="2354" heatid="4463" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" swrid="4992745" athleteid="2326">
              <RESULTS>
                <RESULT eventid="1059" points="677" reactiontime="+80" swimtime="00:00:30.85" resultid="2327" heatid="4266" lane="3" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1094" points="703" reactiontime="+79" swimtime="00:02:49.88" resultid="2328" heatid="4287" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:02:49.88" />
                    <SPLIT distance="150" swimtime="00:02:09.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="618" reactiontime="+89" swimtime="00:00:37.09" resultid="2329" heatid="4312" lane="3" />
                <RESULT eventid="1440" points="749" reactiontime="+83" swimtime="00:00:32.83" resultid="2330" heatid="4374" lane="4" entrytime="00:00:32.06" entrycourse="LCM" />
                <RESULT eventid="1611" points="773" reactiontime="+71" swimtime="00:01:13.89" resultid="2331" heatid="4421" lane="7" entrytime="00:01:12.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-01-05" gender="F" nation="POL" license="502805600055" swrid="4655158" athleteid="2296">
              <RESULTS>
                <RESULT eventid="1059" points="287" reactiontime="+69" swimtime="00:00:40.32" resultid="2297" heatid="4267" lane="4" />
                <RESULT eventid="1233" points="389" reactiontime="+76" swimtime="00:03:44.37" resultid="2298" heatid="4327" lane="2" entrytime="00:03:47.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.64" />
                    <SPLIT distance="100" swimtime="00:01:50.25" />
                    <SPLIT distance="150" swimtime="00:02:48.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="363" reactiontime="+76" swimtime="00:01:43.02" resultid="2299" heatid="4364" lane="1" entrytime="00:01:46.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="2300" heatid="4385" lane="3" />
                <RESULT eventid="1646" status="DNS" swimtime="00:00:00.00" resultid="2301" heatid="4429" lane="3" />
                <RESULT eventid="1680" points="363" reactiontime="+76" swimtime="00:00:47.06" resultid="2302" heatid="4440" lane="2" entrytime="00:00:47.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Morozowski" birthdate="1973-05-09" gender="M" nation="POL" license="102805700051" swrid="5416829" athleteid="2423">
              <RESULTS>
                <RESULT eventid="1163" points="269" reactiontime="+107" swimtime="00:13:26.61" resultid="2424" heatid="4307" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:24.37" />
                    <SPLIT distance="150" swimtime="00:02:13.25" />
                    <SPLIT distance="200" swimtime="00:03:04.48" />
                    <SPLIT distance="250" swimtime="00:03:55.42" />
                    <SPLIT distance="300" swimtime="00:04:47.91" />
                    <SPLIT distance="350" swimtime="00:05:40.16" />
                    <SPLIT distance="400" swimtime="00:06:33.18" />
                    <SPLIT distance="450" swimtime="00:07:25.23" />
                    <SPLIT distance="500" swimtime="00:08:17.52" />
                    <SPLIT distance="550" swimtime="00:09:09.51" />
                    <SPLIT distance="600" swimtime="00:10:01.50" />
                    <SPLIT distance="650" swimtime="00:10:53.82" />
                    <SPLIT distance="700" swimtime="00:11:46.11" />
                    <SPLIT distance="750" swimtime="00:12:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="307" reactiontime="+96" swimtime="00:03:26.78" resultid="2425" heatid="4330" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                    <SPLIT distance="100" swimtime="00:01:36.94" />
                    <SPLIT distance="150" swimtime="00:02:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="305" reactiontime="+91" swimtime="00:01:36.18" resultid="2426" heatid="4366" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="2427" heatid="4417" lane="6" />
                <RESULT eventid="1697" points="380" reactiontime="+100" swimtime="00:00:40.33" resultid="2428" heatid="4442" lane="1" />
                <RESULT eventid="1748" points="279" reactiontime="+106" swimtime="00:06:24.02" resultid="2429" heatid="4463" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:26.02" />
                    <SPLIT distance="150" swimtime="00:02:15.15" />
                    <SPLIT distance="200" swimtime="00:03:05.36" />
                    <SPLIT distance="250" swimtime="00:03:55.42" />
                    <SPLIT distance="300" swimtime="00:04:46.61" />
                    <SPLIT distance="350" swimtime="00:05:36.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" swrid="4754660" athleteid="2303">
              <RESULTS>
                <RESULT eventid="1059" points="567" reactiontime="+86" swimtime="00:00:34.92" resultid="2304" heatid="4270" lane="6" entrytime="00:00:34.31" entrycourse="LCM" />
                <RESULT eventid="1215" points="515" reactiontime="+75" swimtime="00:00:42.23" resultid="2305" heatid="4312" lane="4" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1284" points="551" reactiontime="+91" swimtime="00:01:17.88" resultid="2306" heatid="4338" lane="4" entrytime="00:01:19.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="627" reactiontime="+88" swimtime="00:00:36.34" resultid="2307" heatid="4374" lane="3" entrytime="00:00:36.30" entrycourse="LCM" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1611" points="512" reactiontime="+102" swimtime="00:01:30.10" resultid="2308" heatid="4420" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="558" reactiontime="+101" swimtime="00:00:45.56" resultid="2309" heatid="4439" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Węgrzycka" birthdate="1977-01-26" gender="F" nation="POL" license="502805600056" swrid="5464095" athleteid="2320">
              <RESULTS>
                <RESULT eventid="1059" points="233" reactiontime="+98" swimtime="00:00:43.22" resultid="2321" heatid="4269" lane="8" entrytime="00:00:43.22" entrycourse="LCM" />
                <RESULT eventid="1284" points="177" reactiontime="+95" swimtime="00:01:42.26" resultid="2322" heatid="4337" lane="6" entrytime="00:01:39.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="206" reactiontime="+97" swimtime="00:02:04.53" resultid="2323" heatid="4363" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" reactiontime="+92" status="DNF" swimtime="00:00:00.00" resultid="2324" heatid="4396" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="223" reactiontime="+96" swimtime="00:00:55.31" resultid="2325" heatid="4439" lane="4" entrytime="00:00:53.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="502805600152" swrid="5464091" athleteid="2408">
              <RESULTS>
                <RESULT eventid="1094" points="265" reactiontime="+112" swimtime="00:03:49.85" resultid="2409" heatid="4288" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.27" />
                    <SPLIT distance="100" swimtime="00:01:57.78" />
                    <SPLIT distance="150" swimtime="00:02:59.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="235" reactiontime="+161" swimtime="00:14:53.59" resultid="2410" heatid="4301" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                    <SPLIT distance="100" swimtime="00:01:41.16" />
                    <SPLIT distance="150" swimtime="00:02:37.24" />
                    <SPLIT distance="200" swimtime="00:03:33.88" />
                    <SPLIT distance="250" swimtime="00:04:30.70" />
                    <SPLIT distance="300" swimtime="00:05:27.93" />
                    <SPLIT distance="350" swimtime="00:06:23.64" />
                    <SPLIT distance="400" swimtime="00:07:21.28" />
                    <SPLIT distance="450" swimtime="00:08:18.19" />
                    <SPLIT distance="500" swimtime="00:09:14.74" />
                    <SPLIT distance="550" swimtime="00:10:11.80" />
                    <SPLIT distance="600" swimtime="00:11:08.20" />
                    <SPLIT distance="650" swimtime="00:12:05.54" />
                    <SPLIT distance="700" swimtime="00:13:02.87" />
                    <SPLIT distance="750" swimtime="00:14:01.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="325" reactiontime="+105" swimtime="00:03:58.03" resultid="2411" heatid="4326" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.17" />
                    <SPLIT distance="100" swimtime="00:01:55.99" />
                    <SPLIT distance="150" swimtime="00:02:57.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1335" points="225" reactiontime="+108" swimtime="00:03:57.24" resultid="2412" heatid="4353" lane="3" entrytime="00:04:17.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.13" />
                    <SPLIT distance="150" swimtime="00:02:58.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="277" reactiontime="+106" swimtime="00:03:19.47" resultid="2413" heatid="4396" lane="6" entrytime="00:03:42.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                    <SPLIT distance="100" swimtime="00:01:36.66" />
                    <SPLIT distance="150" swimtime="00:02:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1576" points="259" reactiontime="+94" swimtime="00:08:12.07" resultid="2414" heatid="4413" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.79" />
                    <SPLIT distance="100" swimtime="00:04:16.98" />
                    <SPLIT distance="150" swimtime="00:03:07.69" />
                    <SPLIT distance="200" swimtime="00:06:26.71" />
                    <SPLIT distance="250" swimtime="00:05:22.21" />
                    <SPLIT distance="300" swimtime="00:08:12.07" />
                    <SPLIT distance="350" swimtime="00:07:20.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="150" reactiontime="+136" swimtime="00:04:31.14" resultid="2415" heatid="4429" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.17" />
                    <SPLIT distance="100" swimtime="00:02:15.88" />
                    <SPLIT distance="150" swimtime="00:03:24.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="267" reactiontime="+107" swimtime="00:07:02.23" resultid="2416" heatid="4454" lane="3" entrytime="00:07:44.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                    <SPLIT distance="100" swimtime="00:01:38.04" />
                    <SPLIT distance="150" swimtime="00:02:32.90" />
                    <SPLIT distance="200" swimtime="00:03:26.90" />
                    <SPLIT distance="250" swimtime="00:04:22.25" />
                    <SPLIT distance="300" swimtime="00:05:17.44" />
                    <SPLIT distance="350" swimtime="00:06:12.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Kaczmarek" birthdate="1976-11-27" gender="F" nation="POL" license="502805600149" athleteid="2332">
              <RESULTS>
                <RESULT eventid="1059" points="109" swimtime="00:00:55.70" resultid="2333" heatid="4267" lane="5" />
                <RESULT eventid="1284" points="78" swimtime="00:02:14.29" resultid="2334" heatid="4335" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="129" reactiontime="+60" swimtime="00:02:25.39" resultid="2335" heatid="4362" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="134" swimtime="00:01:05.62" resultid="2336" heatid="4438" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Bednarek" birthdate="1951-03-24" gender="M" nation="POL" license="502805700052" swrid="5464087" athleteid="2363">
              <RESULTS>
                <RESULT eventid="1076" points="460" reactiontime="+101" swimtime="00:00:35.90" resultid="2364" heatid="4277" lane="2" entrytime="00:00:36.84" entrycourse="LCM" />
                <RESULT eventid="1112" points="345" reactiontime="+104" swimtime="00:03:52.23" resultid="2365" heatid="4292" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.86" />
                    <SPLIT distance="100" swimtime="00:01:54.02" />
                    <SPLIT distance="150" swimtime="00:03:02.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="447" reactiontime="+104" swimtime="00:01:22.84" resultid="2366" heatid="4342" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" status="WDR" swimtime="00:00:00.00" resultid="2367" />
                <RESULT eventid="1525" points="431" reactiontime="+108" swimtime="00:03:09.71" resultid="2368" heatid="4399" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                    <SPLIT distance="100" swimtime="00:01:29.04" />
                    <SPLIT distance="150" swimtime="00:02:19.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="395" reactiontime="+109" swimtime="00:06:53.65" resultid="2369" heatid="4462" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                    <SPLIT distance="100" swimtime="00:01:35.43" />
                    <SPLIT distance="150" swimtime="00:02:28.75" />
                    <SPLIT distance="200" swimtime="00:03:23.23" />
                    <SPLIT distance="250" swimtime="00:04:16.48" />
                    <SPLIT distance="300" swimtime="00:05:10.54" />
                    <SPLIT distance="350" swimtime="00:06:03.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Lis - Piwowarski" birthdate="1984-05-29" gender="M" nation="POL" license="502805700146" swrid="5506632" athleteid="2355">
              <RESULTS>
                <RESULT eventid="1076" points="226" reactiontime="+81" swimtime="00:00:37.38" resultid="2356" heatid="4274" lane="0" />
                <RESULT eventid="1267" points="123" reactiontime="+65" swimtime="00:00:53.12" resultid="2357" heatid="4318" lane="7" />
                <RESULT eventid="1301" points="152" reactiontime="+79" swimtime="00:01:35.10" resultid="2358" heatid="4343" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="107" reactiontime="+84" swimtime="00:00:50.85" resultid="2359" heatid="4377" lane="7" />
                <RESULT eventid="1525" points="110" reactiontime="+82" swimtime="00:03:55.69" resultid="2360" heatid="4399" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                    <SPLIT distance="100" swimtime="00:01:46.77" />
                    <SPLIT distance="150" swimtime="00:02:51.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="67" reactiontime="+80" swimtime="00:02:12.13" resultid="2361" heatid="4422" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="105" reactiontime="+82" swimtime="00:08:41.12" resultid="2362" heatid="4463" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.91" />
                    <SPLIT distance="100" swimtime="00:01:54.30" />
                    <SPLIT distance="150" swimtime="00:02:59.00" />
                    <SPLIT distance="200" swimtime="00:04:06.92" />
                    <SPLIT distance="250" swimtime="00:05:16.75" />
                    <SPLIT distance="300" swimtime="00:06:26.57" />
                    <SPLIT distance="350" swimtime="00:07:36.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Piekarski" birthdate="1986-04-22" gender="M" nation="POL" license="502805700144" athleteid="2393">
              <RESULTS>
                <RESULT eventid="1076" points="235" reactiontime="+93" swimtime="00:00:36.89" resultid="2394" heatid="4274" lane="3" />
                <RESULT eventid="1301" points="186" reactiontime="+101" swimtime="00:01:28.89" resultid="2395" heatid="4342" lane="8" />
                <RESULT eventid="1525" points="128" reactiontime="+122" swimtime="00:03:43.86" resultid="2396" heatid="4401" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.18" />
                    <SPLIT distance="100" swimtime="00:01:45.58" />
                    <SPLIT distance="150" swimtime="00:02:46.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dagmara" lastname="Luzniakowska" birthdate="1980-04-29" gender="F" nation="POL" license="102805600154" athleteid="2439">
              <RESULTS>
                <RESULT eventid="1284" points="287" reactiontime="+90" swimtime="00:01:28.01" resultid="2440" heatid="4336" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="180" reactiontime="+97" swimtime="00:00:50.23" resultid="2441" heatid="4372" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Dziedziczak" birthdate="1977-02-04" gender="M" nation="POL" license="502805700153" athleteid="2386">
              <RESULTS>
                <RESULT eventid="1076" points="412" reactiontime="+82" swimtime="00:00:31.64" resultid="2387" heatid="4274" lane="8" />
                <RESULT eventid="1112" status="DNS" swimtime="00:00:00.00" resultid="2388" heatid="4291" lane="5" />
                <RESULT eventid="1267" points="294" reactiontime="+93" swimtime="00:00:41.56" resultid="2389" heatid="4319" lane="9" />
                <RESULT eventid="1301" points="356" reactiontime="+85" swimtime="00:01:13.69" resultid="2390" heatid="4343" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="362" reactiontime="+77" swimtime="00:00:35.40" resultid="2391" heatid="4376" lane="4" />
                <RESULT eventid="1748" points="246" reactiontime="+84" swimtime="00:06:40.89" resultid="2392" heatid="4463" lane="0">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.66" />
                    <SPLIT distance="200" swimtime="00:03:08.19" />
                    <SPLIT distance="300" swimtime="00:04:57.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daria" lastname="Fajkowska" birthdate="1973-03-18" gender="F" nation="POL" license="502805600044" swrid="4992744" athleteid="2337">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="2338" heatid="4267" lane="6" />
                <RESULT eventid="1215" status="DNS" swimtime="00:00:00.00" resultid="2339" heatid="4313" lane="6" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="2340" heatid="4372" lane="2" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="2341" heatid="4386" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tadeusz" lastname="Obiedziński" birthdate="1959-05-12" gender="M" nation="POL" license="502805700040" swrid="4992722" athleteid="2435">
              <RESULTS>
                <RESULT eventid="1250" points="308" reactiontime="+95" swimtime="00:03:57.24" resultid="2436" heatid="4330" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.27" />
                    <SPLIT distance="100" swimtime="00:01:51.25" />
                    <SPLIT distance="150" swimtime="00:02:56.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="338" reactiontime="+91" swimtime="00:01:42.97" resultid="2437" heatid="4366" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="467" reactiontime="+95" swimtime="00:00:42.27" resultid="2438" heatid="4442" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-26" gender="F" nation="POL" license="502805600123" swrid="5464096" athleteid="2310">
              <RESULTS>
                <RESULT eventid="1059" points="159" reactiontime="+125" swimtime="00:00:48.78" resultid="2311" heatid="4268" lane="6" entrytime="00:01:02.85" entrycourse="LCM" />
                <RESULT eventid="1233" points="140" reactiontime="+121" swimtime="00:05:05.00" resultid="2312" heatid="4326" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.40" />
                    <SPLIT distance="100" swimtime="00:02:25.91" />
                    <SPLIT distance="150" swimtime="00:03:47.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="135" reactiontime="+121" swimtime="00:02:21.66" resultid="2313" heatid="4363" lane="3" entrytime="00:02:19.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="145" reactiontime="+116" swimtime="00:01:01.87" resultid="2314" heatid="4438" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Jasiński" birthdate="1960-07-23" gender="M" nation="POL" license="502805700027" swrid="5374015" athleteid="2379">
              <RESULTS>
                <RESULT eventid="1076" points="381" reactiontime="+91" swimtime="00:00:34.79" resultid="2380" heatid="4274" lane="4" />
                <RESULT eventid="1250" points="338" reactiontime="+94" swimtime="00:03:49.86" resultid="2381" heatid="4330" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.70" />
                    <SPLIT distance="100" swimtime="00:01:48.26" />
                    <SPLIT distance="150" swimtime="00:02:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="325" reactiontime="+95" swimtime="00:01:24.07" resultid="2382" heatid="4343" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="333" reactiontime="+78" swimtime="00:01:43.47" resultid="2383" heatid="4366" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="231" reactiontime="+106" swimtime="00:01:47.73" resultid="2384" heatid="4389" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="292" reactiontime="+59" swimtime="00:00:49.42" resultid="2385" heatid="4442" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Dziarek" birthdate="1959-02-19" gender="M" nation="POL" license="502805700029" swrid="4841500" athleteid="2342">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2343" heatid="4278" lane="7" entrytime="00:00:33.56" entrycourse="LCM" />
                <RESULT eventid="1197" status="DNS" swimtime="00:00:00.00" resultid="2344" heatid="4311" lane="5" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="2345" heatid="4345" lane="4" entrytime="00:01:16.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Sikorski" birthdate="1951-05-03" gender="M" nation="POL" license="502805700036" athleteid="2430">
              <RESULTS>
                <RESULT eventid="1267" points="189" reactiontime="+86" swimtime="00:00:58.56" resultid="2431" heatid="4318" lane="5" />
                <RESULT eventid="1406" points="231" reactiontime="+189" swimtime="00:02:13.53" resultid="2432" heatid="4366" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="160" reactiontime="+81" swimtime="00:02:15.31" resultid="2433" heatid="4389" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="289" reactiontime="+104" swimtime="00:00:54.76" resultid="2434" heatid="4442" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Matczak" birthdate="1989-08-12" gender="M" nation="POL" license="502805700" swrid="4071609" athleteid="4120">
              <RESULTS>
                <RESULT eventid="1112" points="605" reactiontime="+72" swimtime="00:02:24.48" resultid="4121" heatid="4296" lane="6" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:09.50" />
                    <SPLIT distance="150" swimtime="00:01:50.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="725" reactiontime="+69" swimtime="00:02:33.68" resultid="4122" heatid="4334" lane="5" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:53.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="657" reactiontime="+76" swimtime="00:01:10.44" resultid="4123" heatid="4371" lane="3" entrytime="00:01:07.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="665" reactiontime="+71" swimtime="00:00:32.02" resultid="4124" heatid="4449" lane="3" entrytime="00:00:30.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Niedźwiedź" birthdate="1963-07-18" gender="M" nation="POL" license="502805700023" swrid="4754661" athleteid="2442">
              <RESULTS>
                <RESULT eventid="1491" points="176" reactiontime="+92" swimtime="00:01:53.33" resultid="2443" heatid="4389" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="181" reactiontime="+91" swimtime="00:04:09.14" resultid="2444" heatid="4433" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.29" />
                    <SPLIT distance="100" swimtime="00:02:02.43" />
                    <SPLIT distance="150" swimtime="00:03:06.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Rembowska-Świeboda" birthdate="1968-06-27" gender="F" nation="POL" license="102805600031" swrid="5439505" athleteid="2315">
              <RESULTS>
                <RESULT eventid="1059" points="490" reactiontime="+72" swimtime="00:00:34.37" resultid="2316" heatid="4268" lane="7" />
                <RESULT eventid="1215" points="524" reactiontime="+86" swimtime="00:00:39.18" resultid="2317" heatid="4313" lane="0" />
                <RESULT eventid="1284" points="461" reactiontime="+77" swimtime="00:01:18.21" resultid="2318" heatid="4335" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="506" reactiontime="+81" swimtime="00:01:25.51" resultid="2319" heatid="4385" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Bartniak" birthdate="1997-11-06" gender="F" nation="POL" license="502805600156" swrid="4287745" athleteid="2403">
              <RESULTS>
                <RESULT eventid="1094" points="614" reactiontime="+81" swimtime="00:02:45.51" resultid="2404" heatid="4287" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:18.59" />
                    <SPLIT distance="150" swimtime="00:02:05.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="585" reactiontime="+79" swimtime="00:03:05.85" resultid="2405" heatid="4326" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                    <SPLIT distance="100" swimtime="00:01:30.38" />
                    <SPLIT distance="150" swimtime="00:02:18.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="570" reactiontime="+78" swimtime="00:01:25.12" resultid="2406" heatid="4363" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1576" points="588" reactiontime="+83" swimtime="00:06:01.40" resultid="2407" heatid="4413" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:26.13" />
                    <SPLIT distance="150" swimtime="00:02:13.37" />
                    <SPLIT distance="200" swimtime="00:02:58.54" />
                    <SPLIT distance="250" swimtime="00:03:47.69" />
                    <SPLIT distance="300" swimtime="00:04:38.04" />
                    <SPLIT distance="350" swimtime="00:05:20.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Wiczel" birthdate="1948-01-22" gender="M" nation="POL" license="502805700021" swrid="4876444" athleteid="2417">
              <RESULTS>
                <RESULT eventid="1163" points="263" reactiontime="+121" swimtime="00:16:35.72" resultid="2418" heatid="4307" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.72" />
                    <SPLIT distance="100" swimtime="00:01:56.85" />
                    <SPLIT distance="150" swimtime="00:03:01.09" />
                    <SPLIT distance="200" swimtime="00:04:06.59" />
                    <SPLIT distance="250" swimtime="00:05:11.58" />
                    <SPLIT distance="300" swimtime="00:06:14.07" />
                    <SPLIT distance="350" swimtime="00:07:17.98" />
                    <SPLIT distance="450" swimtime="00:09:22.40" />
                    <SPLIT distance="500" swimtime="00:10:24.82" />
                    <SPLIT distance="550" swimtime="00:11:26.76" />
                    <SPLIT distance="650" swimtime="00:13:31.77" />
                    <SPLIT distance="750" swimtime="00:15:36.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="557" reactiontime="+111" swimtime="00:03:44.55" resultid="2419" heatid="4329" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.78" />
                    <SPLIT distance="100" swimtime="00:01:48.71" />
                    <SPLIT distance="150" swimtime="00:02:48.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="498" reactiontime="+97" swimtime="00:01:43.46" resultid="2420" heatid="4368" lane="1" entrytime="00:01:40.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="357" reactiontime="+72" swimtime="00:03:46.00" resultid="2421" heatid="4432" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="524" reactiontime="+103" swimtime="00:00:44.92" resultid="2422" heatid="4444" lane="4" entrytime="00:00:42.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1386" points="351" reactiontime="+69" swimtime="00:02:29.45" resultid="2450" heatid="4492" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:01:52.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2397" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2423" number="2" />
                    <RELAYPOSITION athleteid="2386" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2393" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" points="300" reactiontime="+81" swimtime="00:02:21.78" resultid="2455" heatid="4496" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:50.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2355" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2423" number="2" />
                    <RELAYPOSITION athleteid="2386" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2397" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1386" points="531" reactiontime="+92" swimtime="00:02:16.88" resultid="2451" heatid="4492" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:41.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4120" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="2435" number="2" />
                    <RELAYPOSITION athleteid="2346" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2379" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" points="470" reactiontime="+69" swimtime="00:02:06.34" resultid="2456" heatid="4495" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.47" />
                    <SPLIT distance="100" swimtime="00:01:04.26" />
                    <SPLIT distance="150" swimtime="00:01:31.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4120" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2435" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="2346" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2379" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1386" reactiontime="+96" swimtime="00:02:57.52" resultid="2452" heatid="4491" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.83" />
                    <SPLIT distance="100" swimtime="00:01:43.82" />
                    <SPLIT distance="150" swimtime="00:02:20.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2430" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="2417" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2370" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="2363" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" swimtime="00:02:37.58" resultid="2457" heatid="4495" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:01:22.04" />
                    <SPLIT distance="150" swimtime="00:02:03.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2363" number="1" />
                    <RELAYPOSITION athleteid="2430" number="2" />
                    <RELAYPOSITION athleteid="2417" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="2370" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1369" points="368" reactiontime="+85" swimtime="00:02:50.75" resultid="2448" heatid="4490" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.91" />
                    <SPLIT distance="100" swimtime="00:01:37.27" />
                    <SPLIT distance="150" swimtime="00:02:10.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2296" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="2408" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="2403" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="2439" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1542" points="332" reactiontime="+93" swimtime="00:02:37.40" resultid="2453" heatid="4494" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.72" />
                    <SPLIT distance="100" swimtime="00:01:24.95" />
                    <SPLIT distance="150" swimtime="00:02:04.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2408" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="2320" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2439" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2403" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1369" points="549" reactiontime="+79" swimtime="00:02:40.00" resultid="2449" heatid="4490" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:21.12" />
                    <SPLIT distance="150" swimtime="00:01:57.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2315" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2326" number="2" />
                    <RELAYPOSITION athleteid="2303" number="3" reactiontime="+84" />
                    <RELAYPOSITION athleteid="2320" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1542" points="585" reactiontime="+86" swimtime="00:02:18.75" resultid="2454" heatid="4494" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:13.80" />
                    <SPLIT distance="150" swimtime="00:01:47.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2303" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="2296" number="2" />
                    <RELAYPOSITION athleteid="2315" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2326" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" points="387" reactiontime="+102" swimtime="00:02:20.32" resultid="2445" heatid="4489" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="150" swimtime="00:01:52.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2423" number="1" reactiontime="+102" />
                    <RELAYPOSITION athleteid="2439" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2408" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="4120" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1714" points="573" reactiontime="+79" swimtime="00:02:16.31" resultid="2458" heatid="4499" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:01:45.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2303" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4120" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2346" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="2403" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1129" points="499" reactiontime="+74" swimtime="00:02:12.32" resultid="2446" heatid="4488" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:45.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2370" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2296" number="2" />
                    <RELAYPOSITION athleteid="2326" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="2346" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1714" points="328" reactiontime="+83" swimtime="00:02:53.91" resultid="2459" heatid="4498" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.67" />
                    <SPLIT distance="100" swimtime="00:01:35.17" />
                    <SPLIT distance="150" swimtime="00:02:11.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2417" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2296" number="2" />
                    <RELAYPOSITION athleteid="2423" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="2320" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1129" points="451" reactiontime="+85" swimtime="00:02:29.36" resultid="2447" heatid="4488" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                    <SPLIT distance="150" swimtime="00:01:54.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2315" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="2417" number="2" />
                    <RELAYPOSITION athleteid="2435" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2303" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1714" points="594" reactiontime="+80" swimtime="00:02:32.44" resultid="2460" heatid="4498" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:01:22.83" />
                    <SPLIT distance="150" swimtime="00:01:56.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2315" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2370" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="2326" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="2363" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3194" name="JK TEAM Kraków">
          <CONTACT name="Joanna Kwatera" phone="790611187" />
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Zając" birthdate="1984-01-01" gender="M" nation="POL" swrid="5468089" athleteid="3195">
              <RESULTS>
                <RESULT eventid="1076" points="251" reactiontime="+87" swimtime="00:00:36.06" resultid="3196" heatid="4277" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1301" points="259" reactiontime="+88" swimtime="00:01:19.70" resultid="3197" heatid="4345" lane="1" entrytime="00:01:23.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="160" reactiontime="+83" swimtime="00:00:44.51" resultid="3198" heatid="4379" lane="0" entrytime="00:00:45.26" entrycourse="LCM" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="3199" heatid="4402" lane="6" entrytime="00:02:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Tomczuk" birthdate="1980-01-01" gender="M" nation="POL" swrid="5484420" athleteid="3200">
              <RESULTS>
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="3201" heatid="4346" lane="1" entrytime="00:01:14.69" entrycourse="SCM" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="3202" heatid="4404" lane="1" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Wolak" birthdate="1987-01-01" gender="M" nation="POL" swrid="5468088" athleteid="3203">
              <RESULTS>
                <RESULT eventid="1076" points="530" reactiontime="+74" swimtime="00:00:28.12" resultid="3204" heatid="4283" lane="7" entrytime="00:00:27.86" entrycourse="SCM" />
                <RESULT eventid="1301" points="514" reactiontime="+71" swimtime="00:01:03.39" resultid="3205" heatid="4348" lane="5" entrytime="00:01:03.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="479" reactiontime="+75" swimtime="00:00:30.85" resultid="3206" heatid="4381" lane="6" entrytime="00:00:31.08" entrycourse="LCM" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="3207" heatid="4406" lane="5" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2751" name="Sopot Masters">
          <CONTACT name="Goździejewska" />
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Gorbaczow" birthdate="1958-01-01" gender="M" nation="POL" swrid="4191113" athleteid="2752">
              <RESULTS>
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="2753" heatid="4305" lane="2" entrytime="00:13:00.00" />
                <RESULT eventid="1267" points="606" reactiontime="+82" swimtime="00:00:36.15" resultid="2754" heatid="4322" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1301" points="570" reactiontime="+101" swimtime="00:01:09.71" resultid="2755" heatid="4347" lane="9" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="652" reactiontime="+83" swimtime="00:00:31.89" resultid="2756" heatid="4380" lane="1" entrytime="00:00:35.50" />
                <RESULT eventid="1525" points="489" reactiontime="+95" swimtime="00:02:42.02" resultid="2757" heatid="4403" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:17.66" />
                    <SPLIT distance="150" swimtime="00:02:01.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="423" reactiontime="+90" swimtime="00:03:14.67" resultid="2758" heatid="4435" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                    <SPLIT distance="100" swimtime="00:01:36.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3639" name="MOSiR Ostrowiec Św.">
          <CONTACT email="basen@mosir.ostrowiec.pl" name="Różalski Józef" />
          <ATHLETES>
            <ATHLETE firstname="Józef" lastname="Różalski" birthdate="1945-03-28" gender="M" nation="POL" license="501012700001" athleteid="3640">
              <RESULTS>
                <RESULT eventid="1076" points="537" reactiontime="+93" swimtime="00:00:35.92" resultid="3641" heatid="4277" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1112" points="394" reactiontime="+99" swimtime="00:04:02.32" resultid="3642" heatid="4292" lane="2" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.18" />
                    <SPLIT distance="100" swimtime="00:01:53.87" />
                    <SPLIT distance="150" swimtime="00:03:05.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="327" reactiontime="+117" swimtime="00:04:41.55" resultid="3643" heatid="4331" lane="9" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.30" />
                    <SPLIT distance="100" swimtime="00:02:10.98" />
                    <SPLIT distance="150" swimtime="00:03:27.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="383" reactiontime="+93" swimtime="00:01:31.47" resultid="3644" heatid="4344" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="300" reactiontime="+128" swimtime="00:02:11.03" resultid="3645" heatid="4367" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="389" reactiontime="+102" swimtime="00:00:43.48" resultid="3646" heatid="4379" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="1629" points="279" reactiontime="+103" swimtime="00:02:03.48" resultid="3647" heatid="4423" lane="7" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="432" reactiontime="+97" swimtime="00:00:51.65" resultid="3648" heatid="4444" lane="0" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" clubid="3865" name="MKP Szczecin">
          <CONTACT email="windmuhle@wp.pl" name="Kowalczyk Piotr" />
          <ATHLETES>
            <ATHLETE firstname="Szymon" lastname="Kluczyk" birthdate="1987-02-27" gender="M" nation="POL" athleteid="3866">
              <RESULTS>
                <RESULT eventid="1163" points="435" reactiontime="+90" swimtime="00:10:58.08" resultid="3867" heatid="4303" lane="0" entrytime="00:10:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                    <SPLIT distance="150" swimtime="00:03:10.23" />
                    <SPLIT distance="200" swimtime="00:02:30.11" />
                    <SPLIT distance="250" swimtime="00:05:55.39" />
                    <SPLIT distance="300" swimtime="00:03:50.62" />
                    <SPLIT distance="350" swimtime="00:07:20.69" />
                    <SPLIT distance="400" swimtime="00:05:13.07" />
                    <SPLIT distance="450" swimtime="00:08:47.46" />
                    <SPLIT distance="500" swimtime="00:06:37.68" />
                    <SPLIT distance="600" swimtime="00:08:03.37" />
                    <SPLIT distance="700" swimtime="00:09:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="338" reactiontime="+98" swimtime="00:02:55.94" resultid="3868" heatid="4357" lane="9" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                    <SPLIT distance="150" swimtime="00:02:10.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="519" reactiontime="+94" swimtime="00:05:44.22" resultid="3869" heatid="4414" lane="8" entrytime="00:05:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                    <SPLIT distance="150" swimtime="00:02:02.35" />
                    <SPLIT distance="200" swimtime="00:02:46.06" />
                    <SPLIT distance="250" swimtime="00:03:36.71" />
                    <SPLIT distance="300" swimtime="00:04:27.90" />
                    <SPLIT distance="350" swimtime="00:05:07.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="528" reactiontime="+87" swimtime="00:05:04.19" resultid="3870" heatid="4457" lane="1" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:47.80" />
                    <SPLIT distance="200" swimtime="00:02:26.61" />
                    <SPLIT distance="250" swimtime="00:03:06.39" />
                    <SPLIT distance="300" swimtime="00:03:46.14" />
                    <SPLIT distance="350" swimtime="00:04:26.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stefania" lastname="Noetzel" birthdate="1935-08-21" gender="F" nation="POL" athleteid="3876">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1233" points="213" swimtime="00:07:12.20" resultid="3877" heatid="4327" lane="9" entrytime="00:06:42.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:44.96" />
                    <SPLIT distance="100" swimtime="00:03:38.60" />
                    <SPLIT distance="150" swimtime="00:05:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1404" points="153" swimtime="00:03:35.02" resultid="3878" heatid="4363" lane="2" entrytime="00:03:16.80" />
                <RESULT eventid="1680" points="128" swimtime="00:01:42.72" resultid="3879" heatid="4439" lane="7" entrytime="00:01:22.08" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Serbin" birthdate="1966-08-10" gender="F" nation="POL" swrid="4302596" athleteid="3871">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters, Rekord Polski 800 m, 1500m w kat. masters" eventid="1180" points="671" reactiontime="+78" swimtime="00:21:15.24" resultid="3872" heatid="4308" lane="4" entrytime="00:21:01.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:17.08" />
                    <SPLIT distance="150" swimtime="00:01:58.63" />
                    <SPLIT distance="200" swimtime="00:02:40.52" />
                    <SPLIT distance="250" swimtime="00:03:22.77" />
                    <SPLIT distance="300" swimtime="00:04:04.93" />
                    <SPLIT distance="350" swimtime="00:04:47.33" />
                    <SPLIT distance="400" swimtime="00:05:29.79" />
                    <SPLIT distance="450" swimtime="00:06:12.26" />
                    <SPLIT distance="500" swimtime="00:06:54.60" />
                    <SPLIT distance="550" swimtime="00:07:36.93" />
                    <SPLIT distance="600" swimtime="00:08:19.80" />
                    <SPLIT distance="650" swimtime="00:09:02.38" />
                    <SPLIT distance="700" swimtime="00:09:45.12" />
                    <SPLIT distance="750" swimtime="00:10:27.77" />
                    <SPLIT distance="800" swimtime="00:11:10.44" />
                    <SPLIT distance="850" swimtime="00:11:53.62" />
                    <SPLIT distance="900" swimtime="00:12:36.55" />
                    <SPLIT distance="950" swimtime="00:13:19.63" />
                    <SPLIT distance="1000" swimtime="00:14:02.64" />
                    <SPLIT distance="1050" swimtime="00:14:45.54" />
                    <SPLIT distance="1100" swimtime="00:15:28.55" />
                    <SPLIT distance="1150" swimtime="00:16:12.09" />
                    <SPLIT distance="1200" swimtime="00:16:55.66" />
                    <SPLIT distance="1250" swimtime="00:17:39.13" />
                    <SPLIT distance="1300" swimtime="00:18:23.11" />
                    <SPLIT distance="1350" swimtime="00:19:07.10" />
                    <SPLIT distance="1400" swimtime="00:19:50.65" />
                    <SPLIT distance="1450" swimtime="00:20:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1284" points="654" reactiontime="+79" swimtime="00:01:11.44" resultid="3873" heatid="4339" lane="6" entrytime="00:01:13.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="689" reactiontime="+80" swimtime="00:02:34.30" resultid="3874" heatid="4398" lane="2" entrytime="00:02:32.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="150" swimtime="00:01:55.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="679" reactiontime="+79" swimtime="00:05:22.43" resultid="3875" heatid="4452" lane="6" entrytime="00:05:16.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:16.35" />
                    <SPLIT distance="150" swimtime="00:01:57.62" />
                    <SPLIT distance="200" swimtime="00:02:38.99" />
                    <SPLIT distance="250" swimtime="00:03:20.38" />
                    <SPLIT distance="300" swimtime="00:04:02.01" />
                    <SPLIT distance="350" swimtime="00:04:43.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Chmurski" birthdate="1987-09-23" gender="M" nation="POL" swrid="4060941" athleteid="3898">
              <RESULTS>
                <RESULT eventid="1076" points="613" reactiontime="+71" swimtime="00:00:26.80" resultid="3899" heatid="4286" lane="9" entrytime="00:00:26.00" />
                <RESULT eventid="1163" points="536" reactiontime="+83" swimtime="00:10:13.72" resultid="3900" heatid="4303" lane="9" entrytime="00:10:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:46.50" />
                    <SPLIT distance="200" swimtime="00:02:24.77" />
                    <SPLIT distance="250" swimtime="00:03:03.03" />
                    <SPLIT distance="300" swimtime="00:03:41.43" />
                    <SPLIT distance="350" swimtime="00:04:19.96" />
                    <SPLIT distance="400" swimtime="00:04:58.57" />
                    <SPLIT distance="450" swimtime="00:05:38.14" />
                    <SPLIT distance="500" swimtime="00:06:17.28" />
                    <SPLIT distance="550" swimtime="00:06:57.29" />
                    <SPLIT distance="600" swimtime="00:07:37.28" />
                    <SPLIT distance="650" swimtime="00:08:17.83" />
                    <SPLIT distance="700" swimtime="00:08:57.32" />
                    <SPLIT distance="750" swimtime="00:09:36.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="661" reactiontime="+82" swimtime="00:00:58.28" resultid="3901" heatid="4348" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" status="WDR" swimtime="00:00:00.00" resultid="3902" heatid="4406" lane="9" entrytime="00:02:16.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Chałupka" birthdate="1972-08-26" gender="M" nation="POL" athleteid="3903">
              <RESULTS>
                <RESULT eventid="1076" points="534" reactiontime="+89" swimtime="00:00:29.69" resultid="3904" heatid="4281" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1112" points="401" reactiontime="+92" swimtime="00:02:57.89" resultid="3905" heatid="4295" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:20.21" />
                    <SPLIT distance="150" swimtime="00:02:14.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="510" reactiontime="+74" swimtime="00:01:07.77" resultid="3906" heatid="4348" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="510" reactiontime="+84" swimtime="00:00:32.40" resultid="3907" heatid="4382" lane="9" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Szozda" birthdate="1960-01-12" gender="M" nation="POL" athleteid="3880">
              <RESULTS>
                <RESULT eventid="1112" points="387" reactiontime="+97" swimtime="00:03:14.82" resultid="3881" heatid="4294" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                    <SPLIT distance="100" swimtime="00:01:31.31" />
                    <SPLIT distance="150" swimtime="00:02:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="254" reactiontime="+105" swimtime="00:03:46.49" resultid="3882" heatid="4356" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.61" />
                    <SPLIT distance="100" swimtime="00:01:47.52" />
                    <SPLIT distance="150" swimtime="00:02:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="403" reactiontime="+82" swimtime="00:01:29.47" resultid="3883" heatid="4392" lane="0" entrytime="00:01:30.00" />
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="3885" heatid="4424" lane="7" entrytime="00:01:30.00" />
                <RESULT eventid="1697" status="DNS" swimtime="00:00:00.00" resultid="3886" heatid="4445" lane="9" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Kowalczyk" birthdate="1974-10-02" gender="M" nation="POL" swrid="4992788" athleteid="3892">
              <RESULTS>
                <RESULT eventid="1163" points="551" reactiontime="+81" swimtime="00:10:35.36" resultid="3893" heatid="4304" lane="4" entrytime="00:10:34.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                    <SPLIT distance="150" swimtime="00:01:54.55" />
                    <SPLIT distance="200" swimtime="00:02:34.53" />
                    <SPLIT distance="250" swimtime="00:03:13.98" />
                    <SPLIT distance="300" swimtime="00:03:54.33" />
                    <SPLIT distance="350" swimtime="00:04:34.55" />
                    <SPLIT distance="400" swimtime="00:05:14.83" />
                    <SPLIT distance="450" swimtime="00:05:55.05" />
                    <SPLIT distance="500" swimtime="00:06:35.76" />
                    <SPLIT distance="550" swimtime="00:07:16.08" />
                    <SPLIT distance="600" swimtime="00:07:57.30" />
                    <SPLIT distance="650" swimtime="00:08:37.51" />
                    <SPLIT distance="700" swimtime="00:09:18.08" />
                    <SPLIT distance="750" swimtime="00:09:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="523" reactiontime="+79" swimtime="00:01:04.82" resultid="3894" heatid="4348" lane="1" entrytime="00:01:05.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="584" reactiontime="+78" swimtime="00:02:20.87" resultid="3895" heatid="4405" lane="1" entrytime="00:02:20.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" status="WDR" swimtime="00:00:00.00" resultid="3896" heatid="4435" lane="3" entrytime="00:02:55.00" />
                <RESULT eventid="1748" points="577" reactiontime="+81" swimtime="00:05:01.52" resultid="3897" heatid="4458" lane="5" entrytime="00:05:03.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:13.33" />
                    <SPLIT distance="150" swimtime="00:01:51.88" />
                    <SPLIT distance="200" swimtime="00:02:30.95" />
                    <SPLIT distance="250" swimtime="00:03:09.63" />
                    <SPLIT distance="300" swimtime="00:03:48.41" />
                    <SPLIT distance="350" swimtime="00:04:25.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sławomir" lastname="Grzeszewski" birthdate="1953-09-25" gender="M" nation="POL" athleteid="3887">
              <RESULTS>
                <RESULT eventid="1112" points="310" reactiontime="+83" swimtime="00:03:34.64" resultid="3888" heatid="4293" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:01:44.18" />
                    <SPLIT distance="150" swimtime="00:02:44.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="355" reactiontime="+88" swimtime="00:03:48.14" resultid="3889" heatid="4331" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.11" />
                    <SPLIT distance="100" swimtime="00:01:52.57" />
                    <SPLIT distance="150" swimtime="00:02:51.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="406" reactiontime="+78" swimtime="00:01:40.98" resultid="3890" heatid="4368" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="483" reactiontime="+90" swimtime="00:00:42.43" resultid="3891" heatid="4444" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="100111" nation="POL" clubid="3365" name="UKS TRÓJKA Częstochowa">
          <CONTACT city="Częstochowa" email="trojkaczestochowa@o2.pl" name="Gawda" phone="511181791" state="ŚL" street="Schillera 5" zip="42-200" />
          <ATHLETES>
            <ATHLETE firstname="Wiktoria" lastname="Musik" birthdate="1997-08-04" gender="F" nation="POL" license="100111600053" athleteid="3392">
              <RESULTS>
                <RESULT eventid="1059" points="788" reactiontime="+72" swimtime="00:00:27.52" resultid="3393" heatid="4272" lane="5" entrytime="00:00:27.40" />
                <RESULT eventid="1094" points="719" reactiontime="+76" swimtime="00:02:37.09" resultid="3394" heatid="4290" lane="5" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="150" swimtime="00:01:59.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="581" reactiontime="+73" swimtime="00:00:34.02" resultid="3395" heatid="4316" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1284" points="828" reactiontime="+71" swimtime="00:01:00.67" resultid="3396" heatid="4340" lane="5" entrytime="00:01:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="646" reactiontime="+75" swimtime="00:00:30.44" resultid="3397" heatid="4375" lane="1" entrytime="00:00:31.30" />
                <RESULT eventid="1508" points="693" reactiontime="+75" swimtime="00:02:20.76" resultid="3398" heatid="4398" lane="4" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:06.50" />
                    <SPLIT distance="150" swimtime="00:01:44.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="601" reactiontime="+77" swimtime="00:01:11.10" resultid="3399" heatid="4421" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="607" reactiontime="+85" swimtime="00:00:37.32" resultid="3400" heatid="4441" lane="3" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Krogulec" birthdate="1991-07-31" gender="M" nation="POL" athleteid="3375">
              <RESULTS>
                <RESULT eventid="1112" status="DNS" swimtime="00:00:00.00" resultid="3376" heatid="4296" lane="7" entrytime="00:02:38.00" />
                <RESULT eventid="1163" points="364" reactiontime="+96" swimtime="00:11:24.37" resultid="3377" heatid="4304" lane="0" entrytime="00:11:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:03:22.66" />
                    <SPLIT distance="100" swimtime="00:01:16.10" />
                    <SPLIT distance="150" swimtime="00:09:13.91" />
                    <SPLIT distance="200" swimtime="00:02:39.76" />
                    <SPLIT distance="300" swimtime="00:04:05.34" />
                    <SPLIT distance="400" swimtime="00:05:33.05" />
                    <SPLIT distance="500" swimtime="00:07:00.84" />
                    <SPLIT distance="600" swimtime="00:08:29.46" />
                    <SPLIT distance="700" swimtime="00:09:58.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="498" swimtime="00:00:32.77" resultid="3378" heatid="4324" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1457" points="419" reactiontime="+86" swimtime="00:00:31.08" resultid="3379" heatid="4382" lane="7" entrytime="00:00:29.90" />
                <RESULT eventid="1491" points="458" reactiontime="+82" swimtime="00:01:12.55" resultid="3380" heatid="4394" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="458" reactiontime="+86" swimtime="00:02:39.30" resultid="3381" heatid="4437" lane="9" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:01:17.10" />
                    <SPLIT distance="150" swimtime="00:01:59.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="388" reactiontime="+82" swimtime="00:05:26.46" resultid="3382" heatid="4457" lane="0" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:53.56" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:03:18.37" />
                    <SPLIT distance="200" swimtime="00:02:35.31" />
                    <SPLIT distance="300" swimtime="00:04:01.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Warwas" birthdate="1995-07-13" gender="M" nation="POL" license="100111700100" swrid="4266133" athleteid="3409">
              <RESULTS>
                <RESULT eventid="1076" points="661" reactiontime="+70" swimtime="00:00:25.60" resultid="3410" heatid="4282" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1112" points="464" reactiontime="+70" swimtime="00:02:39.71" resultid="3411" heatid="4295" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:02:02.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="554" reactiontime="+73" swimtime="00:00:30.98" resultid="3412" heatid="4324" lane="7" entrytime="00:00:32.60" />
                <RESULT eventid="1491" points="464" reactiontime="+82" swimtime="00:01:11.14" resultid="3413" heatid="4394" lane="8" entrytime="00:01:09.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="370" reactiontime="+74" swimtime="00:06:16.11" resultid="3414" heatid="4414" lane="0" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="150" swimtime="00:02:05.92" />
                    <SPLIT distance="200" swimtime="00:02:58.43" />
                    <SPLIT distance="250" swimtime="00:03:54.24" />
                    <SPLIT distance="300" swimtime="00:04:50.20" />
                    <SPLIT distance="350" swimtime="00:05:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="441" reactiontime="+83" swimtime="00:02:41.31" resultid="3415" heatid="4437" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                    <SPLIT distance="100" swimtime="00:01:17.94" />
                    <SPLIT distance="150" swimtime="00:02:00.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="427" reactiontime="+82" swimtime="00:05:20.05" resultid="3416" heatid="4457" lane="7" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:07.58" />
                    <SPLIT distance="150" swimtime="00:01:45.77" />
                    <SPLIT distance="200" swimtime="00:02:25.51" />
                    <SPLIT distance="250" swimtime="00:03:08.14" />
                    <SPLIT distance="300" swimtime="00:03:51.49" />
                    <SPLIT distance="350" swimtime="00:04:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="640" reactiontime="+70" swimtime="00:00:58.54" resultid="4500" heatid="4352" lane="0" entrytime="00:00:55.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Gajda" birthdate="1995-04-23" gender="M" nation="POL" license="100111700062" athleteid="3366">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3367" heatid="4286" lane="2" entrytime="00:00:25.04" />
                <RESULT eventid="1163" points="544" reactiontime="+71" swimtime="00:10:18.34" resultid="3368" heatid="4303" lane="5" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                    <SPLIT distance="150" swimtime="00:01:42.81" />
                    <SPLIT distance="250" swimtime="00:02:58.49" />
                    <SPLIT distance="350" swimtime="00:04:15.32" />
                    <SPLIT distance="450" swimtime="00:05:34.11" />
                    <SPLIT distance="550" swimtime="00:06:54.73" />
                    <SPLIT distance="650" swimtime="00:08:16.49" />
                    <SPLIT distance="750" swimtime="00:09:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="516" reactiontime="+75" swimtime="00:00:31.71" resultid="3369" heatid="4325" lane="8" entrytime="00:00:31.10" />
                <RESULT eventid="1301" points="709" reactiontime="+71" swimtime="00:00:56.58" resultid="3370" heatid="4352" lane="9" entrytime="00:00:55.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="716" reactiontime="+70" swimtime="00:00:26.50" resultid="3371" heatid="4384" lane="2" entrytime="00:00:26.92" />
                <RESULT eventid="1525" points="676" reactiontime="+71" swimtime="00:02:06.18" resultid="3372" heatid="4407" lane="7" entrytime="00:02:06.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:01.45" />
                    <SPLIT distance="150" swimtime="00:01:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="684" reactiontime="+70" swimtime="00:01:00.26" resultid="3373" heatid="4427" lane="2" entrytime="00:01:00.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="568" reactiontime="+75" swimtime="00:04:50.90" resultid="3374" heatid="4456" lane="6" entrytime="00:04:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:48.39" />
                    <SPLIT distance="200" swimtime="00:02:26.48" />
                    <SPLIT distance="250" swimtime="00:03:04.42" />
                    <SPLIT distance="300" swimtime="00:03:42.39" />
                    <SPLIT distance="350" swimtime="00:04:18.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sonia" lastname="Nowak" birthdate="1996-05-23" gender="F" nation="POL" license="100111600092" athleteid="3401">
              <RESULTS>
                <RESULT eventid="1059" points="548" reactiontime="+86" swimtime="00:00:31.06" resultid="3402" heatid="4271" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1215" points="377" reactiontime="+82" swimtime="00:00:39.29" resultid="3403" heatid="4316" lane="7" entrytime="00:00:34.50" />
                <RESULT eventid="1335" points="529" reactiontime="+96" swimtime="00:02:46.98" resultid="3404" heatid="4354" lane="3" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:17.88" />
                    <SPLIT distance="150" swimtime="00:02:01.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="493" reactiontime="+86" swimtime="00:00:33.32" resultid="3405" heatid="4374" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1508" points="622" reactiontime="+94" swimtime="00:02:25.92" resultid="3406" heatid="4398" lane="3" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:11.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="554" reactiontime="+90" swimtime="00:01:13.05" resultid="3407" heatid="4421" lane="2" entrytime="00:01:11.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="528" reactiontime="+93" swimtime="00:05:20.02" resultid="3408" heatid="4452" lane="2" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:19.04" />
                    <SPLIT distance="150" swimtime="00:02:00.22" />
                    <SPLIT distance="200" swimtime="00:02:41.35" />
                    <SPLIT distance="250" swimtime="00:03:21.90" />
                    <SPLIT distance="300" swimtime="00:04:02.46" />
                    <SPLIT distance="350" swimtime="00:04:41.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kurek" birthdate="1994-07-11" gender="M" nation="POL" license="100111700097" athleteid="3383">
              <RESULTS>
                <RESULT eventid="1076" points="492" reactiontime="+61" swimtime="00:00:28.24" resultid="3384" heatid="4282" lane="0" entrytime="00:00:28.34" />
                <RESULT eventid="1197" points="424" reactiontime="+64" swimtime="00:21:35.75" resultid="3385" heatid="4309" lane="1" entrytime="00:19:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:01:58.10" />
                    <SPLIT distance="200" swimtime="00:02:39.27" />
                    <SPLIT distance="250" swimtime="00:03:21.76" />
                    <SPLIT distance="300" swimtime="00:04:04.17" />
                    <SPLIT distance="350" swimtime="00:04:46.58" />
                    <SPLIT distance="400" swimtime="00:05:29.64" />
                    <SPLIT distance="450" swimtime="00:06:12.90" />
                    <SPLIT distance="500" swimtime="00:06:57.07" />
                    <SPLIT distance="550" swimtime="00:07:40.60" />
                    <SPLIT distance="600" swimtime="00:09:53.86" />
                    <SPLIT distance="650" swimtime="00:09:08.99" />
                    <SPLIT distance="700" swimtime="00:11:22.67" />
                    <SPLIT distance="750" swimtime="00:10:38.72" />
                    <SPLIT distance="800" swimtime="00:12:50.67" />
                    <SPLIT distance="850" swimtime="00:12:06.68" />
                    <SPLIT distance="900" swimtime="00:14:18.66" />
                    <SPLIT distance="950" swimtime="00:13:34.84" />
                    <SPLIT distance="1000" swimtime="00:15:47.36" />
                    <SPLIT distance="1050" swimtime="00:15:02.98" />
                    <SPLIT distance="1100" swimtime="00:17:16.16" />
                    <SPLIT distance="1150" swimtime="00:16:31.60" />
                    <SPLIT distance="1200" swimtime="00:18:45.73" />
                    <SPLIT distance="1250" swimtime="00:18:01.46" />
                    <SPLIT distance="1350" swimtime="00:19:30.33" />
                    <SPLIT distance="1400" swimtime="00:20:13.93" />
                    <SPLIT distance="1450" swimtime="00:20:57.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="349" reactiontime="+74" swimtime="00:00:36.13" resultid="3386" heatid="4323" lane="5" entrytime="00:00:34.20" />
                <RESULT eventid="1301" points="493" reactiontime="+67" swimtime="00:01:03.85" resultid="3387" heatid="4349" lane="1" entrytime="00:01:02.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="390" reactiontime="+64" swimtime="00:00:32.44" resultid="3388" heatid="4381" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="1525" points="477" reactiontime="+60" swimtime="00:02:21.74" resultid="3389" heatid="4404" lane="3" entrytime="00:02:25.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:45.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="407" reactiontime="+69" swimtime="00:00:36.72" resultid="3390" heatid="4448" lane="8" entrytime="00:00:34.20" />
                <RESULT eventid="1748" points="420" reactiontime="+63" swimtime="00:05:21.73" resultid="3391" heatid="4458" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="150" swimtime="00:01:56.18" />
                    <SPLIT distance="200" swimtime="00:02:37.45" />
                    <SPLIT distance="250" swimtime="00:03:18.52" />
                    <SPLIT distance="300" swimtime="00:04:00.81" />
                    <SPLIT distance="350" swimtime="00:04:43.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Chowaniec" birthdate="1995-06-07" gender="M" nation="POL" license="100111700079" athleteid="3417">
              <RESULTS>
                <RESULT eventid="1112" points="534" reactiontime="+74" swimtime="00:02:32.38" resultid="3418" heatid="4296" lane="4" entrytime="00:02:28.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:10.45" />
                    <SPLIT distance="150" swimtime="00:01:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="511" reactiontime="+74" swimtime="00:02:44.86" resultid="3419" heatid="4334" lane="6" entrytime="00:02:33.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:16.74" />
                    <SPLIT distance="150" swimtime="00:02:00.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="559" reactiontime="+75" swimtime="00:01:13.32" resultid="3420" heatid="4371" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="577" reactiontime="+82" swimtime="00:05:24.40" resultid="3421" heatid="4414" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:13.78" />
                    <SPLIT distance="150" swimtime="00:01:56.37" />
                    <SPLIT distance="200" swimtime="00:02:37.59" />
                    <SPLIT distance="250" swimtime="00:03:21.99" />
                    <SPLIT distance="300" swimtime="00:04:07.78" />
                    <SPLIT distance="350" swimtime="00:04:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="599" reactiontime="+75" swimtime="00:00:32.28" resultid="3422" heatid="4449" lane="2" entrytime="00:00:31.57" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1559" points="672" reactiontime="+65" swimtime="00:01:44.96" resultid="3426" heatid="4497" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                    <SPLIT distance="100" swimtime="00:00:54.71" />
                    <SPLIT distance="150" swimtime="00:01:20.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3383" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="3417" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3409" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="3366" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1386" points="705" reactiontime="+79" swimtime="00:01:56.63" resultid="3429" heatid="4493" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:05.64" />
                    <SPLIT distance="150" swimtime="00:01:31.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3375" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="3417" number="2" />
                    <RELAYPOSITION athleteid="3366" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3409" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1714" points="748" reactiontime="+78" swimtime="00:02:03.39" resultid="3423" heatid="4499" lane="5" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:07.00" />
                    <SPLIT distance="150" swimtime="00:01:33.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3392" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3417" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3366" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="3401" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1129" points="763" reactiontime="+67" swimtime="00:01:50.76" resultid="3424" heatid="4489" lane="5" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="150" swimtime="00:01:24.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3409" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3401" number="2" reactiontime="+8" />
                    <RELAYPOSITION athleteid="3392" number="3" />
                    <RELAYPOSITION athleteid="3417" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="01" clubid="2125" name="KS Rekin Świebodzice">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Gajdowska" birthdate="1995-07-17" gender="F" nation="POL" license="102001600173" swrid="4258728" athleteid="2126">
              <RESULTS>
                <RESULT eventid="1059" points="737" reactiontime="+66" swimtime="00:00:28.14" resultid="2127" heatid="4272" lane="6" entrytime="00:00:27.94" entrycourse="LCM" />
                <RESULT eventid="1284" points="833" reactiontime="+67" swimtime="00:01:00.53" resultid="2128" heatid="4340" lane="3" entrytime="00:01:00.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="641" reactiontime="+66" swimtime="00:00:30.52" resultid="2129" heatid="4375" lane="6" entrytime="00:00:30.18" entrycourse="LCM" />
                <RESULT eventid="1508" points="741" reactiontime="+66" swimtime="00:02:17.64" resultid="2130" heatid="4396" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="100" swimtime="00:01:04.34" />
                    <SPLIT distance="150" swimtime="00:01:41.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="562" reactiontime="+69" swimtime="00:00:38.29" resultid="2131" heatid="4438" lane="4" />
                <RESULT eventid="1731" points="704" reactiontime="+68" swimtime="00:04:50.72" resultid="2132" heatid="4454" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="100" swimtime="00:01:08.67" />
                    <SPLIT distance="150" swimtime="00:03:02.11" />
                    <SPLIT distance="200" swimtime="00:02:24.39" />
                    <SPLIT distance="250" swimtime="00:04:17.58" />
                    <SPLIT distance="300" swimtime="00:03:40.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01514" nation="POL" region="14" clubid="2286" name="MPKS Orka Ciechanów">
          <ATHLETES>
            <ATHLETE firstname="Maja" lastname="Dyakowska" birthdate="1996-04-02" gender="F" nation="POL" license="101514600153" swrid="4195195" athleteid="2287">
              <RESULTS>
                <RESULT eventid="1059" points="727" reactiontime="+65" swimtime="00:00:28.27" resultid="2288" heatid="4272" lane="7" entrytime="00:00:28.73" entrycourse="LCM" />
                <RESULT eventid="1284" points="749" reactiontime="+68" swimtime="00:01:02.72" resultid="2289" heatid="4340" lane="6" entrytime="00:01:02.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="102705" nation="POL" clubid="2856" name="Olimpijczyk Tomaszów Mazowiecki Masters">
          <CONTACT email="olimpijczyktomaszow@gmail.com" name="Bucholz" phone="606135860" />
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Bucholz" birthdate="1972-01-26" gender="M" nation="POL" athleteid="2857">
              <RESULTS>
                <RESULT eventid="1112" points="329" reactiontime="+117" swimtime="00:03:09.93" resultid="2858" heatid="4295" lane="0" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                    <SPLIT distance="100" swimtime="00:01:30.60" />
                    <SPLIT distance="150" swimtime="00:02:25.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1197" points="486" reactiontime="+119" swimtime="00:21:47.78" resultid="2859" heatid="4310" lane="3" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="150" swimtime="00:02:03.09" />
                    <SPLIT distance="200" swimtime="00:02:45.71" />
                    <SPLIT distance="250" swimtime="00:03:27.56" />
                    <SPLIT distance="300" swimtime="00:04:09.83" />
                    <SPLIT distance="350" swimtime="00:04:54.09" />
                    <SPLIT distance="400" swimtime="00:05:37.87" />
                    <SPLIT distance="450" swimtime="00:06:21.31" />
                    <SPLIT distance="500" swimtime="00:07:05.07" />
                    <SPLIT distance="550" swimtime="00:07:48.31" />
                    <SPLIT distance="600" swimtime="00:08:32.51" />
                    <SPLIT distance="650" swimtime="00:09:16.95" />
                    <SPLIT distance="700" swimtime="00:10:01.09" />
                    <SPLIT distance="750" swimtime="00:10:45.37" />
                    <SPLIT distance="800" swimtime="00:11:29.88" />
                    <SPLIT distance="850" swimtime="00:12:13.23" />
                    <SPLIT distance="900" swimtime="00:12:56.85" />
                    <SPLIT distance="950" swimtime="00:13:42.34" />
                    <SPLIT distance="1000" swimtime="00:14:27.61" />
                    <SPLIT distance="1050" swimtime="00:15:12.57" />
                    <SPLIT distance="1100" swimtime="00:15:57.09" />
                    <SPLIT distance="1150" swimtime="00:16:40.47" />
                    <SPLIT distance="1200" swimtime="00:17:24.49" />
                    <SPLIT distance="1250" swimtime="00:18:09.47" />
                    <SPLIT distance="1300" swimtime="00:18:54.19" />
                    <SPLIT distance="1350" swimtime="00:19:38.71" />
                    <SPLIT distance="1400" swimtime="00:20:22.89" />
                    <SPLIT distance="1450" swimtime="00:21:06.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="438" reactiontime="+107" swimtime="00:02:36.17" resultid="2860" heatid="4403" lane="1" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:11.44" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="2861" heatid="4416" lane="2" entrytime="00:07:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4097" name="Qswim">
          <CONTACT name="Goździejewska" />
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Rudziński" birthdate="1974-02-12" gender="M" nation="POL" athleteid="4100">
              <RESULTS>
                <RESULT eventid="1197" points="173" reactiontime="+151" swimtime="00:29:51.58" resultid="4101" heatid="4311" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.24" />
                    <SPLIT distance="100" swimtime="00:01:48.07" />
                    <SPLIT distance="150" swimtime="00:02:45.48" />
                    <SPLIT distance="200" swimtime="00:03:43.08" />
                    <SPLIT distance="250" swimtime="00:04:45.59" />
                    <SPLIT distance="300" swimtime="00:05:44.54" />
                    <SPLIT distance="350" swimtime="00:06:45.08" />
                    <SPLIT distance="400" swimtime="00:07:45.28" />
                    <SPLIT distance="450" swimtime="00:08:45.91" />
                    <SPLIT distance="500" swimtime="00:09:45.39" />
                    <SPLIT distance="550" swimtime="00:10:44.99" />
                    <SPLIT distance="600" swimtime="00:11:44.57" />
                    <SPLIT distance="650" swimtime="00:12:44.01" />
                    <SPLIT distance="700" swimtime="00:13:43.00" />
                    <SPLIT distance="750" swimtime="00:14:43.32" />
                    <SPLIT distance="800" swimtime="00:15:43.31" />
                    <SPLIT distance="850" swimtime="00:16:44.09" />
                    <SPLIT distance="900" swimtime="00:17:43.74" />
                    <SPLIT distance="950" swimtime="00:18:45.57" />
                    <SPLIT distance="1000" swimtime="00:19:44.59" />
                    <SPLIT distance="1050" swimtime="00:20:45.02" />
                    <SPLIT distance="1100" swimtime="00:21:45.07" />
                    <SPLIT distance="1150" swimtime="00:22:45.82" />
                    <SPLIT distance="1200" swimtime="00:23:47.22" />
                    <SPLIT distance="1250" swimtime="00:24:48.62" />
                    <SPLIT distance="1300" swimtime="00:25:49.61" />
                    <SPLIT distance="1350" swimtime="00:26:50.45" />
                    <SPLIT distance="1400" swimtime="00:27:50.78" />
                    <SPLIT distance="1450" swimtime="00:28:53.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Kocząb" birthdate="1998-07-26" gender="F" nation="POL" athleteid="4098">
              <RESULTS>
                <RESULT eventid="1180" reactiontime="+136" swimtime="00:30:45.08" resultid="4099" heatid="4308" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.98" />
                    <SPLIT distance="100" swimtime="00:01:48.67" />
                    <SPLIT distance="150" swimtime="00:02:50.06" />
                    <SPLIT distance="200" swimtime="00:03:50.70" />
                    <SPLIT distance="250" swimtime="00:06:55.64" />
                    <SPLIT distance="300" swimtime="00:05:54.60" />
                    <SPLIT distance="350" swimtime="00:08:58.54" />
                    <SPLIT distance="400" swimtime="00:07:55.76" />
                    <SPLIT distance="450" swimtime="00:11:02.34" />
                    <SPLIT distance="500" swimtime="00:09:59.68" />
                    <SPLIT distance="550" swimtime="00:13:07.87" />
                    <SPLIT distance="600" swimtime="00:14:09.19" />
                    <SPLIT distance="650" swimtime="00:15:12.05" />
                    <SPLIT distance="700" swimtime="00:16:13.09" />
                    <SPLIT distance="750" swimtime="00:17:15.51" />
                    <SPLIT distance="800" swimtime="00:18:16.25" />
                    <SPLIT distance="850" swimtime="00:19:18.39" />
                    <SPLIT distance="900" swimtime="00:20:22.94" />
                    <SPLIT distance="950" swimtime="00:21:25.06" />
                    <SPLIT distance="1000" swimtime="00:22:27.66" />
                    <SPLIT distance="1050" swimtime="00:23:32.12" />
                    <SPLIT distance="1100" swimtime="00:24:33.20" />
                    <SPLIT distance="1150" swimtime="00:25:36.28" />
                    <SPLIT distance="1200" swimtime="00:26:39.21" />
                    <SPLIT distance="1250" swimtime="00:27:42.19" />
                    <SPLIT distance="1300" swimtime="00:28:44.17" />
                    <SPLIT distance="1350" swimtime="00:29:46.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="3060" name="Marijampoles &quot;TORPEDOS&quot;">
          <CONTACT email="klubastorpedos@gmail.com" name="Vilmantas Krasauskas" phone="+37068746068" street="R. Jukneviciaus mg.78-10" street2="Marijampole" />
          <ATHLETES>
            <ATHLETE firstname="Stasys" lastname="Grigas" birthdate="1941-03-14" gender="M" nation="LTU" athleteid="3061">
              <RESULTS>
                <RESULT eventid="1076" points="160" reactiontime="+134" swimtime="00:00:58.86" resultid="3062" heatid="4275" lane="3" entrytime="00:00:58.65" entrycourse="LCM" />
                <RESULT eventid="1163" status="WDR" swimtime="00:00:00.00" resultid="3063" heatid="4306" lane="7" entrytime="00:25:10.00" entrycourse="LCM" />
                <RESULT eventid="1267" points="139" reactiontime="+126" swimtime="00:01:13.65" resultid="3064" heatid="4320" lane="9" entrytime="00:01:12.91" entrycourse="LCM" />
                <RESULT eventid="1301" points="117" reactiontime="+116" swimtime="00:02:26.90" resultid="3065" heatid="4343" lane="4" entrytime="00:02:30.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="150" reactiontime="+122" swimtime="00:02:42.76" resultid="3066" heatid="4390" lane="0" entrytime="00:02:41.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="100" reactiontime="+120" swimtime="00:05:44.75" resultid="3067" heatid="4401" lane="2" entrytime="00:05:41.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.62" />
                    <SPLIT distance="100" swimtime="00:02:54.92" />
                    <SPLIT distance="150" swimtime="00:04:27.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="180" reactiontime="+119" swimtime="00:05:45.55" resultid="3068" heatid="4433" lane="2" entrytime="00:05:49.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.90" />
                    <SPLIT distance="100" swimtime="00:02:52.86" />
                    <SPLIT distance="150" swimtime="00:04:24.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="104" reactiontime="+116" swimtime="00:12:13.85" resultid="3069" heatid="4462" lane="5" entrytime="00:13:39.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.41" />
                    <SPLIT distance="100" swimtime="00:02:54.82" />
                    <SPLIT distance="150" swimtime="00:04:29.43" />
                    <SPLIT distance="200" swimtime="00:06:07.42" />
                    <SPLIT distance="250" swimtime="00:07:43.08" />
                    <SPLIT distance="300" swimtime="00:09:18.95" />
                    <SPLIT distance="350" swimtime="00:10:52.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laimute" lastname="Paludneviciene" birthdate="1963-01-21" gender="F" nation="LTU" athleteid="3080">
              <RESULTS>
                <RESULT eventid="1215" points="215" reactiontime="+83" swimtime="00:00:53.36" resultid="3081" heatid="4314" lane="1" entrytime="00:00:53.81" entrycourse="LCM" />
                <RESULT eventid="1680" points="305" reactiontime="+109" swimtime="00:00:53.40" resultid="3082" heatid="4440" lane="9" entrytime="00:00:53.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valdimaras" lastname="Paludnevicius" birthdate="1947-03-24" gender="M" nation="LTU" athleteid="3083">
              <RESULTS>
                <RESULT eventid="1076" points="364" reactiontime="+109" swimtime="00:00:40.88" resultid="3084" heatid="4276" lane="2" entrytime="00:00:44.00" entrycourse="LCM" />
                <RESULT eventid="1267" points="402" reactiontime="+83" swimtime="00:00:46.67" resultid="3085" heatid="4321" lane="0" entrytime="00:00:46.33" entrycourse="LCM" />
                <RESULT eventid="1491" points="411" reactiontime="+120" swimtime="00:01:43.79" resultid="3086" heatid="4391" lane="9" entrytime="00:01:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jurate" lastname="Pranckeviciene" birthdate="1975-05-04" gender="F" nation="LTU" athleteid="3070">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="3071" heatid="4270" lane="0" entrytime="00:00:35.08" entrycourse="LCM" />
                <RESULT eventid="1284" status="DNS" swimtime="00:00:00.00" resultid="3072" heatid="4338" lane="6" entrytime="00:01:20.16" entrycourse="LCM" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="3073" heatid="4397" lane="7" entrytime="00:03:04.78" entrycourse="LCM" />
                <RESULT eventid="1646" status="DNS" swimtime="00:00:00.00" resultid="3074" heatid="4430" lane="7" entrytime="00:03:50.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vilmantas" lastname="Krasauskas" birthdate="1964-07-31" gender="M" nation="LTU" athleteid="3075">
              <RESULTS>
                <RESULT eventid="1076" points="541" reactiontime="+80" swimtime="00:00:30.01" resultid="3076" heatid="4280" lane="7" entrytime="00:00:30.01" entrycourse="LCM" />
                <RESULT eventid="1301" points="615" reactiontime="+81" swimtime="00:01:05.86" resultid="3077" heatid="4348" lane="9" entrytime="00:01:05.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="567" reactiontime="+76" swimtime="00:02:29.80" resultid="3078" heatid="4404" lane="6" entrytime="00:02:25.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:12.64" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="553" reactiontime="+81" swimtime="00:05:19.78" resultid="3079" heatid="4459" lane="2" entrytime="00:05:25.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:15.86" />
                    <SPLIT distance="150" swimtime="00:01:55.79" />
                    <SPLIT distance="200" swimtime="00:02:37.02" />
                    <SPLIT distance="250" swimtime="00:03:18.33" />
                    <SPLIT distance="300" swimtime="00:04:00.08" />
                    <SPLIT distance="350" swimtime="00:04:41.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00905" nation="POL" clubid="3431" name="MKS Trójka Łódź">
          <CONTACT name="Melka" phone="600276930" />
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Szwedzki" birthdate="2000-12-12" gender="M" nation="POL" license="100905700604" swrid="4001538" athleteid="3432">
              <RESULTS>
                <RESULT eventid="1112" reactiontime="+70" swimtime="00:02:18.67" resultid="3433" heatid="4297" lane="6" entrytime="00:02:16.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:01:06.76" />
                    <SPLIT distance="150" swimtime="00:01:46.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1197" reactiontime="+75" swimtime="00:17:48.91" resultid="3434" heatid="4309" lane="5" entrytime="00:17:15.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:08.91" />
                    <SPLIT distance="150" swimtime="00:01:44.92" />
                    <SPLIT distance="200" swimtime="00:02:20.17" />
                    <SPLIT distance="250" swimtime="00:02:54.81" />
                    <SPLIT distance="300" swimtime="00:03:30.01" />
                    <SPLIT distance="350" swimtime="00:04:05.03" />
                    <SPLIT distance="400" swimtime="00:04:40.11" />
                    <SPLIT distance="450" swimtime="00:05:14.85" />
                    <SPLIT distance="500" swimtime="00:05:49.83" />
                    <SPLIT distance="550" swimtime="00:06:24.66" />
                    <SPLIT distance="600" swimtime="00:06:59.62" />
                    <SPLIT distance="650" swimtime="00:07:34.79" />
                    <SPLIT distance="700" swimtime="00:08:10.16" />
                    <SPLIT distance="750" swimtime="00:08:45.27" />
                    <SPLIT distance="800" swimtime="00:09:20.86" />
                    <SPLIT distance="850" swimtime="00:09:56.57" />
                    <SPLIT distance="900" swimtime="00:10:32.27" />
                    <SPLIT distance="950" swimtime="00:11:08.31" />
                    <SPLIT distance="1000" swimtime="00:11:44.34" />
                    <SPLIT distance="1050" swimtime="00:12:20.10" />
                    <SPLIT distance="1100" swimtime="00:12:56.68" />
                    <SPLIT distance="1150" swimtime="00:13:33.30" />
                    <SPLIT distance="1200" swimtime="00:14:09.58" />
                    <SPLIT distance="1250" swimtime="00:14:46.07" />
                    <SPLIT distance="1300" swimtime="00:15:22.59" />
                    <SPLIT distance="1350" swimtime="00:15:58.79" />
                    <SPLIT distance="1400" swimtime="00:16:35.19" />
                    <SPLIT distance="1450" swimtime="00:17:12.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" reactiontime="+73" swimtime="00:02:50.77" resultid="3435" heatid="4334" lane="2" entrytime="00:02:36.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                    <SPLIT distance="100" swimtime="00:01:22.20" />
                    <SPLIT distance="150" swimtime="00:02:06.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" reactiontime="+74" swimtime="00:02:25.05" resultid="3436" heatid="4357" lane="4" entrytime="00:02:17.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:08.85" />
                    <SPLIT distance="150" swimtime="00:01:47.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" reactiontime="+71" swimtime="00:02:04.86" resultid="3437" heatid="4407" lane="3" entrytime="00:02:03.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                    <SPLIT distance="100" swimtime="00:01:00.81" />
                    <SPLIT distance="150" swimtime="00:01:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" reactiontime="+80" swimtime="00:05:30.18" resultid="3438" heatid="4414" lane="3" entrytime="00:04:56.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:17.29" />
                    <SPLIT distance="150" swimtime="00:02:04.42" />
                    <SPLIT distance="200" swimtime="00:02:50.33" />
                    <SPLIT distance="250" swimtime="00:03:27.17" />
                    <SPLIT distance="300" swimtime="00:04:07.74" />
                    <SPLIT distance="350" swimtime="00:04:49.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" reactiontime="+72" swimtime="00:02:49.00" resultid="3439" heatid="4437" lane="6" entrytime="00:02:23.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:01:23.04" />
                    <SPLIT distance="150" swimtime="00:02:06.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" reactiontime="+69" swimtime="00:04:16.88" resultid="3440" heatid="4456" lane="3" entrytime="00:04:20.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                    <SPLIT distance="100" swimtime="00:04:36.59" />
                    <SPLIT distance="150" swimtime="00:01:33.44" />
                    <SPLIT distance="250" swimtime="00:02:39.84" />
                    <SPLIT distance="350" swimtime="00:03:47.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UKS SPARTA" nation="POL" clubid="3441" name="UKS Sparta Grodzisk Mazowicki">
          <CONTACT city="Grodzisk Mazowiecki" email="sherry@interia.pl" internet="www.spartiaci.pl" name="Wolnicki Robert" phone="533544534" state="MAZ" street="Zondka 6" zip="05-825" />
          <ATHLETES>
            <ATHLETE firstname="Karol" lastname="Zieliński" birthdate="1980-05-18" gender="M" nation="POL" athleteid="3442">
              <RESULTS>
                <RESULT eventid="1250" points="458" reactiontime="+91" swimtime="00:02:59.76" resultid="3443" heatid="4333" lane="2" entrytime="00:02:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:12.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K15" eventid="1406" reactiontime="+96" status="DSQ" swimtime="00:00:00.00" resultid="3444" heatid="4369" lane="4" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" status="DNS" swimtime="00:00:00.00" resultid="3445" heatid="4447" lane="7" entrytime="00:00:35.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Głowa" birthdate="1979-10-08" gender="M" nation="POL" athleteid="3446">
              <RESULTS>
                <RESULT eventid="1301" points="541" reactiontime="+84" swimtime="00:01:02.85" resultid="3447" heatid="4349" lane="0" entrytime="00:01:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="463" reactiontime="+86" swimtime="00:02:26.95" resultid="3448" heatid="4406" lane="8" entrytime="00:02:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                    <SPLIT distance="100" swimtime="00:01:10.37" />
                    <SPLIT distance="150" swimtime="00:01:47.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="4092" name="Dzukijos vandenis">
          <CONTACT name="Goździejewska" />
          <ATHLETES>
            <ATHLETE firstname="Sigitas" lastname="Katkevicius" birthdate="1957-08-05" gender="M" nation="LTU" swrid="4418116" athleteid="4093">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1250" points="736" reactiontime="+80" swimtime="00:02:58.94" resultid="4094" heatid="4333" lane="1" entrytime="00:02:58.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:27.27" />
                    <SPLIT distance="150" swimtime="00:02:14.17" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1525" points="709" reactiontime="+77" swimtime="00:02:25.08" resultid="4095" heatid="4403" lane="4" entrytime="00:02:30.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:10.55" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="734" reactiontime="+77" swimtime="00:00:36.91" resultid="4096" heatid="4447" lane="9" entrytime="00:00:36.78" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" clubid="2862" name="Uks Cityzen">
          <CONTACT name="Pietraszewski" phone="501648415" />
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Pietraszewski" birthdate="1955-04-07" gender="M" nation="POL" swrid="4187282" athleteid="2878">
              <RESULTS>
                <RESULT eventid="1112" points="300" reactiontime="+91" swimtime="00:03:37.00" resultid="2879" heatid="4293" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.69" />
                    <SPLIT distance="100" swimtime="00:01:43.42" />
                    <SPLIT distance="150" swimtime="00:02:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="360" reactiontime="+98" swimtime="00:14:19.38" resultid="2880" heatid="4305" lane="7" entrytime="00:13:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:37.11" />
                    <SPLIT distance="150" swimtime="00:02:30.06" />
                    <SPLIT distance="200" swimtime="00:03:23.46" />
                    <SPLIT distance="250" swimtime="00:04:16.80" />
                    <SPLIT distance="300" swimtime="00:05:10.67" />
                    <SPLIT distance="350" swimtime="00:06:04.75" />
                    <SPLIT distance="400" swimtime="00:06:59.78" />
                    <SPLIT distance="450" swimtime="00:07:54.09" />
                    <SPLIT distance="500" swimtime="00:08:48.31" />
                    <SPLIT distance="550" swimtime="00:09:44.97" />
                    <SPLIT distance="600" swimtime="00:10:40.60" />
                    <SPLIT distance="650" swimtime="00:11:35.80" />
                    <SPLIT distance="700" swimtime="00:12:30.51" />
                    <SPLIT distance="750" swimtime="00:13:27.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="284" reactiontime="+97" swimtime="00:00:47.07" resultid="2881" heatid="4321" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1491" points="385" reactiontime="+84" swimtime="00:01:35.96" resultid="2882" heatid="4391" lane="6" entrytime="00:01:35.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="2883" heatid="4416" lane="6" entrytime="00:07:15.00" />
                <RESULT eventid="1663" points="429" reactiontime="+98" swimtime="00:03:28.35" resultid="2884" heatid="4434" lane="6" entrytime="00:03:24.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.02" />
                    <SPLIT distance="100" swimtime="00:01:42.65" />
                    <SPLIT distance="150" swimtime="00:02:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="2885" heatid="4460" lane="9" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Matyszczak" birthdate="1970-12-14" gender="M" nation="POL" swrid="5471729" athleteid="2890">
              <RESULTS>
                <RESULT eventid="1076" points="461" reactiontime="+89" swimtime="00:00:31.18" resultid="2891" heatid="4280" lane="0" entrytime="00:00:30.99" entrycourse="LCM" />
                <RESULT eventid="1112" points="245" reactiontime="+99" swimtime="00:03:29.55" resultid="2892" heatid="4294" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:35.08" />
                    <SPLIT distance="150" swimtime="00:02:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="323" reactiontime="+89" swimtime="00:00:41.64" resultid="2893" heatid="4322" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1301" points="401" reactiontime="+94" swimtime="00:01:13.46" resultid="2894" heatid="4346" lane="6" entrytime="00:01:12.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="329" reactiontime="+96" swimtime="00:02:51.84" resultid="2896" heatid="4402" lane="4" entrytime="00:02:51.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:08.95" />
                    <SPLIT distance="100" swimtime="00:02:51.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="258" reactiontime="+96" swimtime="00:03:31.31" resultid="2897" heatid="4435" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:40.59" />
                    <SPLIT distance="150" swimtime="00:02:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="288" reactiontime="+101" swimtime="00:06:27.38" resultid="2898" heatid="4459" lane="8" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:13.27" />
                    <SPLIT distance="100" swimtime="00:03:03.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="300" reactiontime="+84" swimtime="00:01:31.98" resultid="3672" heatid="4391" lane="5" entrytime="00:01:33.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Rybak-Starczak" birthdate="1975-01-16" gender="F" nation="POL" swrid="5439532" athleteid="2868">
              <RESULTS>
                <RESULT eventid="1094" points="478" reactiontime="+96" swimtime="00:03:08.68" resultid="2869" heatid="4289" lane="6" entrytime="00:03:11.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                    <SPLIT distance="100" swimtime="00:01:31.72" />
                    <SPLIT distance="150" swimtime="00:02:26.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="482" reactiontime="+122" swimtime="00:03:28.83" resultid="2870" heatid="4328" lane="0" entrytime="00:03:24.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                    <SPLIT distance="100" swimtime="00:01:41.20" />
                    <SPLIT distance="150" swimtime="00:02:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="421" reactiontime="+119" swimtime="00:01:38.06" resultid="2871" heatid="4365" lane="9" entrytime="00:01:35.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Łutowicz" birthdate="1950-08-23" gender="F" nation="POL" swrid="4188428" athleteid="2863">
              <RESULTS>
                <RESULT eventid="1059" points="247" swimtime="00:00:48.95" resultid="2864" heatid="4269" lane="0" entrytime="00:00:43.39" entrycourse="LCM" />
                <RESULT eventid="1215" points="259" reactiontime="+61" swimtime="00:00:54.38" resultid="2865" heatid="4314" lane="0" entrytime="00:01:00.00" />
                <RESULT eventid="1284" points="261" swimtime="00:01:44.73" resultid="2866" heatid="4337" lane="2" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="268" swimtime="00:02:01.01" resultid="2867" heatid="4387" lane="1" entrytime="00:02:04.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Boryski" birthdate="1951-03-05" gender="M" nation="POL" swrid="4754708" athleteid="2872">
              <RESULTS>
                <RESULT eventid="1197" points="338" reactiontime="+103" swimtime="00:29:20.34" resultid="2873" heatid="4310" lane="8" entrytime="00:29:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.79" />
                    <SPLIT distance="100" swimtime="00:01:51.88" />
                    <SPLIT distance="150" swimtime="00:02:51.24" />
                    <SPLIT distance="200" swimtime="00:03:49.73" />
                    <SPLIT distance="250" swimtime="00:04:47.88" />
                    <SPLIT distance="300" swimtime="00:05:46.67" />
                    <SPLIT distance="350" swimtime="00:06:44.59" />
                    <SPLIT distance="400" swimtime="00:07:43.76" />
                    <SPLIT distance="450" swimtime="00:08:43.04" />
                    <SPLIT distance="500" swimtime="00:09:43.13" />
                    <SPLIT distance="550" swimtime="00:10:41.52" />
                    <SPLIT distance="600" swimtime="00:11:41.33" />
                    <SPLIT distance="650" swimtime="00:12:40.31" />
                    <SPLIT distance="700" swimtime="00:13:39.77" />
                    <SPLIT distance="750" swimtime="00:14:39.45" />
                    <SPLIT distance="800" swimtime="00:15:38.99" />
                    <SPLIT distance="850" swimtime="00:16:38.03" />
                    <SPLIT distance="900" swimtime="00:17:37.17" />
                    <SPLIT distance="950" swimtime="00:18:36.10" />
                    <SPLIT distance="1000" swimtime="00:19:35.39" />
                    <SPLIT distance="1050" swimtime="00:20:34.56" />
                    <SPLIT distance="1100" swimtime="00:21:34.99" />
                    <SPLIT distance="1150" swimtime="00:22:32.52" />
                    <SPLIT distance="1200" swimtime="00:23:31.17" />
                    <SPLIT distance="1250" swimtime="00:24:30.77" />
                    <SPLIT distance="1300" swimtime="00:25:30.30" />
                    <SPLIT distance="1350" swimtime="00:26:28.23" />
                    <SPLIT distance="1400" swimtime="00:27:27.35" />
                    <SPLIT distance="1450" swimtime="00:28:25.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="369" reactiontime="+82" swimtime="00:00:46.80" resultid="2874" heatid="4321" lane="1" entrytime="00:00:45.56" entrycourse="LCM" />
                <RESULT eventid="1491" points="286" reactiontime="+82" swimtime="00:01:51.48" resultid="2875" heatid="4391" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" status="DNS" swimtime="00:00:00.00" resultid="2876" heatid="4434" lane="0" entrytime="00:03:53.23" entrycourse="LCM" />
                <RESULT eventid="1748" points="314" reactiontime="+93" swimtime="00:07:26.63" resultid="2877" heatid="4461" lane="8" entrytime="00:07:39.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.64" />
                    <SPLIT distance="100" swimtime="00:01:42.61" />
                    <SPLIT distance="150" swimtime="00:02:40.73" />
                    <SPLIT distance="200" swimtime="00:03:38.43" />
                    <SPLIT distance="250" swimtime="00:04:36.12" />
                    <SPLIT distance="300" swimtime="00:05:33.34" />
                    <SPLIT distance="350" swimtime="00:06:31.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sławomir" lastname="Cybertowicz" birthdate="1966-01-12" gender="M" nation="POL" swrid="4269915" athleteid="2886">
              <RESULTS>
                <RESULT eventid="1250" points="374" reactiontime="+94" swimtime="00:03:29.04" resultid="2887" heatid="4332" lane="1" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:41.68" />
                    <SPLIT distance="150" swimtime="00:02:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="302" reactiontime="+90" swimtime="00:01:40.79" resultid="2888" heatid="4369" lane="8" entrytime="00:01:26.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="362" reactiontime="+91" swimtime="00:00:42.13" resultid="2889" heatid="4445" lane="4" entrytime="00:00:38.62" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1386" points="352" reactiontime="+77" swimtime="00:02:46.28" resultid="2899" heatid="4492" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.22" />
                    <SPLIT distance="100" swimtime="00:01:32.29" />
                    <SPLIT distance="150" swimtime="00:02:09.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2872" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2890" number="2" reactiontime="+6" />
                    <RELAYPOSITION athleteid="2886" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="2878" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" points="427" swimtime="00:02:32.09" resultid="2900" heatid="4488" lane="6" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.75" />
                    <SPLIT distance="100" swimtime="00:01:24.33" />
                    <SPLIT distance="150" swimtime="00:01:59.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2863" number="1" />
                    <RELAYPOSITION athleteid="2878" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="2868" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="2886" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="05806" nation="POL" region="06" clubid="1929" name="IKS Druga Strona Sportu">
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Rupp" birthdate="1956-03-06" gender="F" nation="POL" license="505806600021" swrid="5484417" athleteid="2708">
              <RESULTS>
                <RESULT eventid="1094" points="169" reactiontime="+110" swimtime="00:05:10.09" resultid="2709" heatid="4288" lane="6" entrytime="00:04:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.78" />
                    <SPLIT distance="100" swimtime="00:02:27.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="229" reactiontime="+128" swimtime="00:17:42.50" resultid="2710" heatid="4302" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.06" />
                    <SPLIT distance="100" swimtime="00:02:06.31" />
                    <SPLIT distance="150" swimtime="00:03:13.16" />
                    <SPLIT distance="200" swimtime="00:04:19.64" />
                    <SPLIT distance="250" swimtime="00:05:26.61" />
                    <SPLIT distance="300" swimtime="00:06:33.80" />
                    <SPLIT distance="350" swimtime="00:07:40.59" />
                    <SPLIT distance="400" swimtime="00:08:48.02" />
                    <SPLIT distance="450" swimtime="00:09:55.21" />
                    <SPLIT distance="500" swimtime="00:11:02.86" />
                    <SPLIT distance="550" swimtime="00:12:10.30" />
                    <SPLIT distance="600" swimtime="00:13:17.94" />
                    <SPLIT distance="650" swimtime="00:14:25.40" />
                    <SPLIT distance="700" swimtime="00:15:32.70" />
                    <SPLIT distance="750" swimtime="00:16:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="164" reactiontime="+87" swimtime="00:01:01.31" resultid="2711" heatid="4314" lane="9" entrytime="00:01:02.95" entrycourse="SCM" />
                <RESULT eventid="1284" points="172" reactiontime="+113" swimtime="00:01:56.75" resultid="2712" heatid="4337" lane="7" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="81" reactiontime="+119" swimtime="00:01:16.07" resultid="2713" heatid="4373" lane="8" entrytime="00:01:12.00" />
                <RESULT eventid="1474" points="165" reactiontime="+77" swimtime="00:02:15.74" resultid="2714" heatid="4387" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="203" reactiontime="+80" swimtime="00:04:45.25" resultid="2715" heatid="4430" lane="0" entrytime="00:08:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.11" />
                    <SPLIT distance="100" swimtime="00:02:22.90" />
                    <SPLIT distance="150" swimtime="00:03:34.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3248" name="Max Masters Karol Bartkowiak">
          <CONTACT city="Szamotuły" email="karolbartkowiak88@gmail.com" name="Bartkowiak" phone="721573722" state="WLKP" street="Wojska Polskiego 9b/14" zip="64-500" />
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Sędrowicz" birthdate="1997-05-17" gender="M" nation="POL" athleteid="3249">
              <RESULTS>
                <RESULT eventid="1076" points="459" reactiontime="+76" swimtime="00:00:28.91" resultid="3250" heatid="4281" lane="6" entrytime="00:00:29.00" />
                <RESULT comment="Z3G8" eventid="1112" reactiontime="+80" status="DSQ" swimtime="00:00:00.00" resultid="3251" heatid="4295" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                    <SPLIT distance="100" swimtime="00:03:05.65" />
                    <SPLIT distance="150" swimtime="00:02:16.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="333" reactiontime="+80" swimtime="00:03:10.03" resultid="3252" heatid="4333" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:30.11" />
                    <SPLIT distance="150" swimtime="00:02:20.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="394" reactiontime="+75" swimtime="00:01:08.80" resultid="3253" heatid="4347" lane="0" entrytime="00:01:10.00" />
                <RESULT eventid="1406" points="410" reactiontime="+74" swimtime="00:01:21.30" resultid="3254" heatid="4370" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="3255" heatid="4416" lane="5" entrytime="00:07:00.00" />
                <RESULT eventid="1663" status="DNS" swimtime="00:00:00.00" resultid="3256" heatid="4433" lane="3" entrytime="00:04:55.00" />
                <RESULT eventid="1697" points="437" reactiontime="+71" swimtime="00:00:35.85" resultid="3257" heatid="4448" lane="1" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02706" nation="POL" region="06" clubid="2533" name="UKS ,,Jasień&apos;&apos; Sucha Beskidzka">
          <ATHLETES>
            <ATHLETE firstname="Aneta" lastname="Pytel" birthdate="1979-02-03" gender="F" nation="POL" license="102706600133" athleteid="2534">
              <RESULTS>
                <RESULT eventid="1059" points="246" reactiontime="+73" swimtime="00:00:42.22" resultid="2535" heatid="4268" lane="0" />
                <RESULT comment="Z3/G8" eventid="1094" reactiontime="+74" status="DSQ" swimtime="00:00:00.00" resultid="2536" heatid="4287" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.75" />
                    <SPLIT distance="100" swimtime="00:01:56.93" />
                    <SPLIT distance="150" swimtime="00:03:05.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="197" reactiontime="+80" swimtime="00:00:50.92" resultid="2537" heatid="4313" lane="8" />
                <RESULT eventid="1284" points="185" reactiontime="+74" swimtime="00:01:41.92" resultid="2538" heatid="4336" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="267" reactiontime="+78" swimtime="00:01:52.92" resultid="2539" heatid="4363" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="192" reactiontime="+81" swimtime="00:01:52.20" resultid="2540" heatid="4385" lane="7" />
                <RESULT eventid="1680" points="278" reactiontime="+70" swimtime="00:00:49.76" resultid="2541" heatid="4438" lane="7" />
                <RESULT eventid="1731" points="177" reactiontime="+80" swimtime="00:07:48.08" resultid="2542" heatid="4455" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.67" />
                    <SPLIT distance="100" swimtime="00:01:46.51" />
                    <SPLIT distance="150" swimtime="00:02:44.37" />
                    <SPLIT distance="200" swimtime="00:03:44.89" />
                    <SPLIT distance="250" swimtime="00:04:46.88" />
                    <SPLIT distance="300" swimtime="00:05:48.52" />
                    <SPLIT distance="350" swimtime="00:06:50.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sabina" lastname="Sikora" birthdate="1984-10-03" gender="F" nation="POL" license="102706600159" swrid="5468086" athleteid="2543">
              <RESULTS>
                <RESULT eventid="1059" points="649" reactiontime="+79" swimtime="00:00:30.01" resultid="2544" heatid="4271" lane="1" entrytime="00:00:32.31" entrycourse="LCM" />
                <RESULT eventid="1094" points="441" reactiontime="+93" swimtime="00:03:05.79" resultid="2545" heatid="4288" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="150" swimtime="00:02:21.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="474" reactiontime="+98" swimtime="00:00:36.71" resultid="2546" heatid="4313" lane="1" />
                <RESULT eventid="1233" points="453" reactiontime="+68" swimtime="00:03:22.34" resultid="2547" heatid="4326" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="100" swimtime="00:01:37.84" />
                    <SPLIT distance="150" swimtime="00:02:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="576" reactiontime="+81" swimtime="00:01:26.95" resultid="2548" heatid="4365" lane="1" entrytime="00:01:34.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="406" reactiontime="+92" swimtime="00:01:23.36" resultid="2549" heatid="4386" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="688" reactiontime="+76" swimtime="00:00:37.01" resultid="2550" heatid="4441" lane="0" entrytime="00:00:42.21" entrycourse="LCM" />
                <RESULT eventid="1731" points="414" reactiontime="+68" swimtime="00:05:57.17" resultid="2551" heatid="4455" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                    <SPLIT distance="100" swimtime="00:01:25.16" />
                    <SPLIT distance="150" swimtime="00:02:10.87" />
                    <SPLIT distance="200" swimtime="00:02:57.13" />
                    <SPLIT distance="250" swimtime="00:03:43.71" />
                    <SPLIT distance="300" swimtime="00:04:30.36" />
                    <SPLIT distance="350" swimtime="00:05:16.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LCGW" nation="POL" clubid="3275" name="Landsberg Crew Gorzów Wlkp.">
          <CONTACT city="Os. Poznańskie" email="landsbergcrew@gmail.com" name="Kaczmarek" phone="600277732" state="LUB" street="Liliowa 9" zip="66-446" />
          <ATHLETES>
            <ATHLETE firstname="Stanislaw" lastname="Kaczmarek" birthdate="1979-01-26" gender="M" nation="POL" license="501304700001" swrid="4432188" athleteid="3276">
              <RESULTS>
                <RESULT eventid="1112" points="715" reactiontime="+74" swimtime="00:02:26.09" resultid="3277" heatid="4297" lane="1" entrytime="00:02:22.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="100" swimtime="00:01:09.80" />
                    <SPLIT distance="150" swimtime="00:01:52.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="650" reactiontime="+76" swimtime="00:09:55.58" resultid="3278" heatid="4303" lane="3" entrytime="00:09:29.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:11.89" />
                    <SPLIT distance="150" swimtime="00:01:49.61" />
                    <SPLIT distance="200" swimtime="00:02:27.63" />
                    <SPLIT distance="250" swimtime="00:03:06.13" />
                    <SPLIT distance="300" swimtime="00:03:44.08" />
                    <SPLIT distance="350" swimtime="00:04:22.45" />
                    <SPLIT distance="400" swimtime="00:05:00.60" />
                    <SPLIT distance="450" swimtime="00:05:38.40" />
                    <SPLIT distance="500" swimtime="00:06:16.39" />
                    <SPLIT distance="550" swimtime="00:06:54.12" />
                    <SPLIT distance="600" swimtime="00:07:31.11" />
                    <SPLIT distance="650" swimtime="00:08:07.37" />
                    <SPLIT distance="700" swimtime="00:08:44.13" />
                    <SPLIT distance="750" swimtime="00:09:20.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="545" reactiontime="+81" swimtime="00:02:49.66" resultid="3279" heatid="4334" lane="9" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                    <SPLIT distance="100" swimtime="00:01:20.40" />
                    <SPLIT distance="150" swimtime="00:02:04.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="531" reactiontime="+76" swimtime="00:02:35.08" resultid="3280" heatid="4357" lane="5" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:14.55" />
                    <SPLIT distance="150" swimtime="00:01:56.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="618" reactiontime="+75" swimtime="00:02:13.42" resultid="3281" heatid="4407" lane="8" entrytime="00:02:07.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                    <SPLIT distance="100" swimtime="00:01:04.65" />
                    <SPLIT distance="150" swimtime="00:01:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="679" reactiontime="+73" swimtime="00:05:21.95" resultid="3282" heatid="4414" lane="6" entrytime="00:05:12.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:10.33" />
                    <SPLIT distance="150" swimtime="00:01:56.28" />
                    <SPLIT distance="200" swimtime="00:02:39.35" />
                    <SPLIT distance="250" swimtime="00:03:26.06" />
                    <SPLIT distance="300" swimtime="00:04:12.76" />
                    <SPLIT distance="350" swimtime="00:04:48.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="588" reactiontime="+74" swimtime="00:00:34.42" resultid="3283" heatid="4448" lane="5" entrytime="00:00:33.33" />
                <RESULT eventid="1748" points="657" reactiontime="+76" swimtime="00:04:43.86" resultid="3284" heatid="4456" lane="2" entrytime="00:04:36.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:08.63" />
                    <SPLIT distance="150" swimtime="00:01:45.50" />
                    <SPLIT distance="200" swimtime="00:02:21.53" />
                    <SPLIT distance="250" swimtime="00:02:57.21" />
                    <SPLIT distance="300" swimtime="00:03:33.29" />
                    <SPLIT distance="350" swimtime="00:04:09.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="3995" name="Ukraine Swim Team">
          <ATHLETES>
            <ATHLETE firstname="DIANA" lastname="MILINKOVSKA" birthdate="1974-01-01" gender="F" nation="UKR" athleteid="3999">
              <RESULTS>
                <RESULT eventid="1094" points="650" reactiontime="+95" swimtime="00:02:50.32" resultid="4010" heatid="4290" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:20.03" />
                    <SPLIT distance="150" swimtime="00:02:11.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="553" reactiontime="+86" swimtime="00:01:21.70" resultid="4011" heatid="4388" lane="7" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="472" reactiontime="+88" swimtime="00:01:23.41" resultid="4012" heatid="4421" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1335" points="405" reactiontime="+93" swimtime="00:03:15.14" resultid="4013" heatid="4354" lane="7" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:32.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="WDR" swimtime="00:00:00.00" resultid="4014" entrytime="00:02:49.00" />
                <RESULT eventid="1646" points="550" reactiontime="+76" swimtime="00:02:55.81" resultid="5037" heatid="4431" lane="3" entrytime="00:02:49.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                    <SPLIT distance="100" swimtime="00:01:25.50" />
                    <SPLIT distance="150" swimtime="00:02:11.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="OLHA" lastname="TSETSENOVA" birthdate="1974-01-01" gender="F" nation="UKR" athleteid="4113">
              <RESULTS>
                <RESULT eventid="1146" points="199" reactiontime="+98" swimtime="00:15:44.97" resultid="5039" heatid="4302" lane="7" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                    <SPLIT distance="100" swimtime="00:01:41.49" />
                    <SPLIT distance="150" swimtime="00:02:39.06" />
                    <SPLIT distance="200" swimtime="00:03:38.72" />
                    <SPLIT distance="250" swimtime="00:04:39.42" />
                    <SPLIT distance="300" swimtime="00:05:40.15" />
                    <SPLIT distance="350" swimtime="00:06:40.75" />
                    <SPLIT distance="400" swimtime="00:07:41.22" />
                    <SPLIT distance="450" swimtime="00:08:40.55" />
                    <SPLIT distance="500" swimtime="00:09:42.00" />
                    <SPLIT distance="550" swimtime="00:10:42.91" />
                    <SPLIT distance="600" swimtime="00:11:43.75" />
                    <SPLIT distance="650" swimtime="00:12:43.52" />
                    <SPLIT distance="700" swimtime="00:13:43.87" />
                    <SPLIT distance="750" swimtime="00:14:46.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="324" reactiontime="+92" swimtime="00:03:58.38" resultid="5040" heatid="4327" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.51" />
                    <SPLIT distance="100" swimtime="00:01:55.86" />
                    <SPLIT distance="150" swimtime="00:02:58.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="285" reactiontime="+106" swimtime="00:01:51.65" resultid="5041" heatid="4364" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="263" reactiontime="+96" swimtime="00:03:23.13" resultid="5042" heatid="4396" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                    <SPLIT distance="100" swimtime="00:01:35.25" />
                    <SPLIT distance="150" swimtime="00:02:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="217" reactiontime="+100" swimtime="00:07:32.38" resultid="5043" heatid="4454" lane="4" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.59" />
                    <SPLIT distance="100" swimtime="00:01:46.42" />
                    <SPLIT distance="150" swimtime="00:02:44.30" />
                    <SPLIT distance="200" swimtime="00:03:42.88" />
                    <SPLIT distance="250" swimtime="00:04:41.89" />
                    <SPLIT distance="300" swimtime="00:05:40.96" />
                    <SPLIT distance="350" swimtime="00:06:41.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="IRYNA" lastname="ORIEKHOVA" birthdate="1988-01-01" gender="F" nation="UKR" athleteid="3996">
              <RESULTS>
                <RESULT eventid="1094" points="289" reactiontime="+86" swimtime="00:03:22.55" resultid="4015" heatid="4289" lane="1" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.84" />
                    <SPLIT distance="100" swimtime="00:01:33.90" />
                    <SPLIT distance="150" swimtime="00:02:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="281" reactiontime="+94" swimtime="00:03:47.44" resultid="4016" heatid="4327" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.70" />
                    <SPLIT distance="100" swimtime="00:01:50.96" />
                    <SPLIT distance="150" swimtime="00:02:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="267" reactiontime="+91" swimtime="00:03:09.97" resultid="4017" heatid="4397" lane="8" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                    <SPLIT distance="100" swimtime="00:01:28.92" />
                    <SPLIT distance="150" swimtime="00:02:20.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="246" reactiontime="+95" swimtime="00:06:52.70" resultid="4018" heatid="4453" lane="0" entrytime="00:06:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:24.93" />
                    <SPLIT distance="200" swimtime="00:03:19.67" />
                    <SPLIT distance="250" swimtime="00:04:13.83" />
                    <SPLIT distance="300" swimtime="00:05:07.64" />
                    <SPLIT distance="350" swimtime="00:06:01.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="OLENA" lastname="RUDNYTSKA" birthdate="1964-01-01" gender="F" nation="UKR" athleteid="3998">
              <RESULTS>
                <RESULT eventid="1508" points="201" reactiontime="+115" swimtime="00:03:52.70" resultid="4019" heatid="4396" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.96" />
                    <SPLIT distance="100" swimtime="00:01:46.67" />
                    <SPLIT distance="150" swimtime="00:02:50.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="196" reactiontime="+108" swimtime="00:08:07.94" resultid="4020" heatid="4454" lane="2" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.13" />
                    <SPLIT distance="100" swimtime="00:01:53.63" />
                    <SPLIT distance="150" swimtime="00:02:56.52" />
                    <SPLIT distance="200" swimtime="00:03:59.16" />
                    <SPLIT distance="250" swimtime="00:05:02.36" />
                    <SPLIT distance="300" swimtime="00:06:04.54" />
                    <SPLIT distance="350" swimtime="00:07:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="189" swimtime="00:16:59.49" resultid="4021" heatid="4301" lane="3" entrytime="00:16:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.72" />
                    <SPLIT distance="100" swimtime="00:01:52.47" />
                    <SPLIT distance="150" swimtime="00:02:55.78" />
                    <SPLIT distance="200" swimtime="00:03:59.08" />
                    <SPLIT distance="250" swimtime="00:05:02.75" />
                    <SPLIT distance="300" swimtime="00:08:16.42" />
                    <SPLIT distance="350" swimtime="00:07:10.58" />
                    <SPLIT distance="400" swimtime="00:12:36.93" />
                    <SPLIT distance="450" swimtime="00:09:20.13" />
                    <SPLIT distance="500" swimtime="00:14:46.97" />
                    <SPLIT distance="550" swimtime="00:11:31.44" />
                    <SPLIT distance="650" swimtime="00:13:41.72" />
                    <SPLIT distance="750" swimtime="00:15:51.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="IRYNA" lastname="DOMANOVA " birthdate="1982-01-01" gender="F" nation="UKR" athleteid="4000">
              <RESULTS>
                <RESULT eventid="1094" points="392" reactiontime="+102" swimtime="00:03:18.24" resultid="4001" heatid="4289" lane="2" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:32.85" />
                    <SPLIT distance="150" swimtime="00:02:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="358" reactiontime="+85" swimtime="00:00:41.72" resultid="4002" heatid="4315" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="1404" points="379" reactiontime="+89" swimtime="00:01:40.52" resultid="4003" heatid="4364" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="277" reactiontime="+107" swimtime="00:01:37.22" resultid="4004" heatid="4420" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="NATALIA" lastname="BORYSHKEVYCH" birthdate="1976-01-01" gender="F" nation="UKR" athleteid="3997">
              <RESULTS>
                <RESULT eventid="1180" points="460" reactiontime="+85" swimtime="00:22:39.98" resultid="4005" heatid="4308" lane="3" entrytime="00:23:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:21.50" />
                    <SPLIT distance="150" swimtime="00:02:06.32" />
                    <SPLIT distance="200" swimtime="00:02:51.46" />
                    <SPLIT distance="250" swimtime="00:03:37.67" />
                    <SPLIT distance="300" swimtime="00:04:23.17" />
                    <SPLIT distance="350" swimtime="00:06:41.96" />
                    <SPLIT distance="400" swimtime="00:05:55.40" />
                    <SPLIT distance="450" swimtime="00:08:14.57" />
                    <SPLIT distance="500" swimtime="00:07:27.94" />
                    <SPLIT distance="550" swimtime="00:09:47.56" />
                    <SPLIT distance="600" swimtime="00:09:00.64" />
                    <SPLIT distance="650" swimtime="00:11:20.02" />
                    <SPLIT distance="700" swimtime="00:10:33.81" />
                    <SPLIT distance="750" swimtime="00:12:52.29" />
                    <SPLIT distance="800" swimtime="00:12:06.03" />
                    <SPLIT distance="850" swimtime="00:14:24.78" />
                    <SPLIT distance="900" swimtime="00:13:38.53" />
                    <SPLIT distance="950" swimtime="00:15:57.73" />
                    <SPLIT distance="1000" swimtime="00:15:11.19" />
                    <SPLIT distance="1050" swimtime="00:17:29.63" />
                    <SPLIT distance="1100" swimtime="00:16:43.76" />
                    <SPLIT distance="1150" swimtime="00:19:02.16" />
                    <SPLIT distance="1200" swimtime="00:18:15.94" />
                    <SPLIT distance="1250" swimtime="00:20:32.22" />
                    <SPLIT distance="1300" swimtime="00:19:47.50" />
                    <SPLIT distance="1350" swimtime="00:21:59.40" />
                    <SPLIT distance="1400" swimtime="00:21:16.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="496" reactiontime="+73" swimtime="00:01:12.52" resultid="4006" heatid="4339" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="387" reactiontime="+79" swimtime="00:00:38.98" resultid="4007" heatid="4374" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1508" points="535" reactiontime="+63" swimtime="00:02:40.22" resultid="4008" heatid="4398" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:01:16.88" />
                    <SPLIT distance="150" swimtime="00:01:58.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" status="DNS" swimtime="00:00:00.00" resultid="4009" heatid="4452" lane="7" entrytime="00:05:25.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="4023" heatid="4495" lane="3" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1369" points="512" reactiontime="+84" swimtime="00:02:35.95" resultid="4022" heatid="4490" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:25.50" />
                    <SPLIT distance="150" swimtime="00:02:03.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4000" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3996" number="2" />
                    <RELAYPOSITION athleteid="3999" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3997" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1542" points="500" reactiontime="+62" swimtime="00:02:16.61" resultid="4024" heatid="4494" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:45.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3997" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4000" number="2" />
                    <RELAYPOSITION athleteid="3996" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3999" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4214" nation="POL" clubid="2901" name="Warsaw Masters team">
          <CONTACT email="marlena@masters.waw.pl" name="Dobrasiewicz-Iwaniuk" />
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Pfitzner" birthdate="1986-05-24" gender="M" nation="POL" athleteid="3023">
              <RESULTS>
                <RESULT eventid="1301" points="601" reactiontime="+73" swimtime="00:01:00.18" resultid="3024" heatid="4350" lane="5" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="536" reactiontime="+82" swimtime="00:01:11.27" resultid="3025" heatid="4393" lane="4" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="3026" heatid="4425" lane="2" entrytime="00:01:11.00" />
                <RESULT eventid="1748" points="578" reactiontime="+76" swimtime="00:04:55.16" resultid="3027" heatid="4457" lane="4" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:09.91" />
                    <SPLIT distance="150" swimtime="00:01:47.70" />
                    <SPLIT distance="200" swimtime="00:02:25.89" />
                    <SPLIT distance="250" swimtime="00:03:04.53" />
                    <SPLIT distance="300" swimtime="00:03:43.11" />
                    <SPLIT distance="350" swimtime="00:04:19.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Porada" birthdate="1983-06-10" gender="M" nation="POL" athleteid="2931">
              <RESULTS>
                <RESULT eventid="1076" points="511" reactiontime="+72" swimtime="00:00:28.46" resultid="2932" heatid="4282" lane="7" entrytime="00:00:28.18" />
                <RESULT eventid="1112" points="520" reactiontime="+71" swimtime="00:02:36.23" resultid="2933" heatid="4296" lane="9" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:15.68" />
                    <SPLIT distance="150" swimtime="00:01:59.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="597" reactiontime="+71" swimtime="00:02:46.62" resultid="2934" heatid="4333" lane="4" entrytime="00:02:47.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:19.47" />
                    <SPLIT distance="150" swimtime="00:02:02.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="561" reactiontime="+67" swimtime="00:01:15.66" resultid="2935" heatid="4370" lane="6" entrytime="00:01:16.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="567" reactiontime="+68" swimtime="00:00:34.40" resultid="2936" heatid="4448" lane="6" entrytime="00:00:33.65" />
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="2937" heatid="4458" lane="1" entrytime="00:05:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szymański" birthdate="1981-11-04" gender="M" nation="POL" athleteid="2954">
              <RESULTS>
                <RESULT eventid="1076" points="547" reactiontime="+83" swimtime="00:00:28.43" resultid="2955" heatid="4282" lane="9" entrytime="00:00:28.90" />
                <RESULT eventid="1267" points="431" reactiontime="+95" swimtime="00:00:35.92" resultid="2956" heatid="4323" lane="6" entrytime="00:00:34.50" />
                <RESULT eventid="1457" points="555" reactiontime="+83" swimtime="00:00:30.49" resultid="2957" heatid="4381" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1697" points="350" reactiontime="+89" swimtime="00:00:40.91" resultid="2958" heatid="4445" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Giejsztowt" birthdate="1978-06-13" gender="M" nation="POL" athleteid="2959">
              <RESULTS>
                <RESULT eventid="1076" points="554" reactiontime="+73" swimtime="00:00:28.31" resultid="2960" heatid="4281" lane="1" entrytime="00:00:29.20" />
                <RESULT eventid="1301" points="561" reactiontime="+69" swimtime="00:01:02.08" resultid="2961" heatid="4349" lane="7" entrytime="00:01:02.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="541" reactiontime="+70" swimtime="00:02:19.51" resultid="2962" heatid="4405" lane="6" entrytime="00:02:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:43.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="545" reactiontime="+72" swimtime="00:05:02.08" resultid="2963" heatid="4458" lane="4" entrytime="00:05:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="150" swimtime="00:01:51.27" />
                    <SPLIT distance="200" swimtime="00:02:30.18" />
                    <SPLIT distance="250" swimtime="00:03:09.12" />
                    <SPLIT distance="300" swimtime="00:03:48.53" />
                    <SPLIT distance="350" swimtime="00:04:26.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Burdelak" birthdate="1991-07-06" gender="F" nation="POL" athleteid="2976">
              <RESULTS>
                <RESULT eventid="1215" points="534" reactiontime="+63" swimtime="00:00:35.21" resultid="2977" heatid="4316" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1233" points="527" reactiontime="+69" swimtime="00:03:04.36" resultid="2978" heatid="4328" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:30.23" />
                    <SPLIT distance="150" swimtime="00:02:17.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="615" reactiontime="+68" swimtime="00:01:22.45" resultid="2979" heatid="4365" lane="3" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="634" reactiontime="+68" swimtime="00:00:31.98" resultid="2980" heatid="4375" lane="0" entrytime="00:00:31.80" />
                <RESULT eventid="1611" points="346" reactiontime="+73" swimtime="00:01:23.81" resultid="2981" heatid="4421" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="633" reactiontime="+68" swimtime="00:00:37.52" resultid="2982" heatid="4441" lane="5" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Nowak" birthdate="1952-12-17" gender="M" nation="POL" athleteid="3012">
              <RESULTS>
                <RESULT eventid="1112" points="478" reactiontime="+88" swimtime="00:03:28.40" resultid="3013" heatid="4293" lane="5" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                    <SPLIT distance="100" swimtime="00:01:47.97" />
                    <SPLIT distance="150" swimtime="00:02:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="658" reactiontime="+100" swimtime="00:03:32.48" resultid="3014" heatid="4332" lane="0" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.70" />
                    <SPLIT distance="100" swimtime="00:01:39.63" />
                    <SPLIT distance="150" swimtime="00:02:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="711" reactiontime="+97" swimtime="00:01:31.85" resultid="3015" heatid="4368" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="401" reactiontime="+93" swimtime="00:08:02.62" resultid="3016" heatid="4416" lane="1" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.72" />
                    <SPLIT distance="100" swimtime="00:02:02.88" />
                    <SPLIT distance="150" swimtime="00:05:12.78" />
                    <SPLIT distance="200" swimtime="00:04:13.57" />
                    <SPLIT distance="300" swimtime="00:06:14.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="781" reactiontime="+79" swimtime="00:00:39.32" resultid="3017" heatid="4445" lane="5" entrytime="00:00:38.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Kozak" birthdate="1986-02-13" gender="M" nation="POL" swrid="4992669" athleteid="2983">
              <RESULTS>
                <RESULT eventid="1250" points="516" reactiontime="+92" swimtime="00:02:54.88" resultid="2984" heatid="4333" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:26.87" />
                    <SPLIT distance="150" swimtime="00:02:12.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="596" reactiontime="+87" swimtime="00:01:14.14" resultid="2985" heatid="4369" lane="2" entrytime="00:01:22.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="674" reactiontime="+76" swimtime="00:00:32.47" resultid="2986" heatid="4447" lane="3" entrytime="00:00:34.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Jarecka-Skorykow" birthdate="1974-01-30" gender="F" nation="POL" swrid="4992672" athleteid="3043">
              <RESULTS>
                <RESULT eventid="1404" points="467" reactiontime="+82" swimtime="00:01:34.73" resultid="3044" heatid="4364" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Dargas-Miszczak" birthdate="1981-09-06" gender="F" nation="POL" athleteid="2987">
              <RESULTS>
                <RESULT eventid="1059" points="448" reactiontime="+80" swimtime="00:00:34.55" resultid="2988" heatid="4270" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1094" points="392" reactiontime="+83" swimtime="00:03:18.10" resultid="2989" heatid="4289" lane="0" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:01:39.74" />
                    <SPLIT distance="150" swimtime="00:02:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="446" reactiontime="+88" swimtime="00:01:15.97" resultid="2990" heatid="4338" lane="8" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="455" reactiontime="+84" swimtime="00:00:36.87" resultid="2991" heatid="4374" lane="0" entrytime="00:00:39.80" />
                <RESULT eventid="1508" points="411" reactiontime="+85" swimtime="00:02:53.89" resultid="2992" heatid="4397" lane="5" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:24.36" />
                    <SPLIT distance="150" swimtime="00:02:11.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="328" reactiontime="+74" swimtime="00:01:31.91" resultid="2993" heatid="4420" lane="7" entrytime="00:01:36.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="365" reactiontime="+88" swimtime="00:06:07.92" resultid="2994" heatid="4453" lane="6" entrytime="00:06:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:01:28.00" />
                    <SPLIT distance="150" swimtime="00:02:14.80" />
                    <SPLIT distance="200" swimtime="00:03:02.58" />
                    <SPLIT distance="250" swimtime="00:03:50.40" />
                    <SPLIT distance="300" swimtime="00:04:38.16" />
                    <SPLIT distance="350" swimtime="00:05:24.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Paluszak" birthdate="1967-02-17" gender="M" nation="POL" swrid="5471792" athleteid="2947">
              <RESULTS>
                <RESULT eventid="1112" points="246" reactiontime="+80" swimtime="00:03:44.57" resultid="2948" heatid="4293" lane="8" entrytime="00:03:50.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                    <SPLIT distance="100" swimtime="00:01:46.35" />
                    <SPLIT distance="150" swimtime="00:02:50.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="242" reactiontime="+75" swimtime="00:00:42.64" resultid="2950" heatid="4379" lane="1" entrytime="00:00:44.25" />
                <RESULT eventid="1593" points="239" reactiontime="+92" swimtime="00:08:06.26" resultid="2951" heatid="4417" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.13" />
                    <SPLIT distance="100" swimtime="00:01:58.75" />
                    <SPLIT distance="150" swimtime="00:03:04.57" />
                    <SPLIT distance="200" swimtime="00:04:10.30" />
                    <SPLIT distance="250" swimtime="00:05:12.30" />
                    <SPLIT distance="300" swimtime="00:06:15.56" />
                    <SPLIT distance="350" swimtime="00:07:10.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="2952" heatid="4423" lane="5" entrytime="00:01:46.31" />
                <RESULT eventid="1748" points="209" reactiontime="+81" swimtime="00:07:22.05" resultid="2953" heatid="4461" lane="1" entrytime="00:07:26.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                    <SPLIT distance="100" swimtime="00:01:43.95" />
                    <SPLIT distance="150" swimtime="00:02:39.59" />
                    <SPLIT distance="200" swimtime="00:03:35.40" />
                    <SPLIT distance="250" swimtime="00:04:32.15" />
                    <SPLIT distance="300" swimtime="00:05:28.62" />
                    <SPLIT distance="350" swimtime="00:06:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="232" reactiontime="+77" swimtime="00:01:31.16" resultid="4112" heatid="4343" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leszk" lastname="Madej" birthdate="1960-06-17" gender="M" nation="POL" athleteid="2902">
              <RESULTS>
                <RESULT eventid="1076" points="689" reactiontime="+80" swimtime="00:00:28.57" resultid="2903" heatid="4282" lane="2" entrytime="00:00:28.11" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1112" points="670" reactiontime="+83" swimtime="00:02:42.23" resultid="2904" heatid="4295" lane="3" entrytime="00:02:42.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="150" swimtime="00:02:03.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="592" reactiontime="+72" swimtime="00:00:36.44" resultid="2905" heatid="4323" lane="8" entrytime="00:00:35.21" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1301" points="796" reactiontime="+78" swimtime="00:01:02.35" resultid="2906" heatid="4348" lane="4" entrytime="00:01:03.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1525" points="777" reactiontime="+80" swimtime="00:02:18.90" resultid="2907" heatid="4405" lane="7" entrytime="00:02:20.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:08.51" />
                    <SPLIT distance="150" swimtime="00:01:43.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="2908" heatid="4415" lane="1" entrytime="00:06:15.37" />
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="2909" heatid="4425" lane="0" entrytime="00:01:14.21" />
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="2910" heatid="4458" lane="3" entrytime="00:05:05.71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" swrid="5506635" athleteid="3000">
              <RESULTS>
                <RESULT eventid="1076" points="693" reactiontime="+76" swimtime="00:00:26.61" resultid="3001" heatid="4284" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1301" points="623" reactiontime="+76" swimtime="00:01:01.17" resultid="3002" heatid="4349" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="672" reactiontime="+72" swimtime="00:01:13.93" resultid="3003" heatid="4370" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="480" reactiontime="+74" swimtime="00:02:30.37" resultid="3004" heatid="4404" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:50.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="689" reactiontime="+65" swimtime="00:00:33.09" resultid="3005" heatid="4449" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1748" points="415" reactiontime="+82" swimtime="00:05:36.72" resultid="3006" heatid="4459" lane="9" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                    <SPLIT distance="200" swimtime="00:02:43.64" />
                    <SPLIT distance="250" swimtime="00:03:27.64" />
                    <SPLIT distance="300" swimtime="00:04:10.98" />
                    <SPLIT distance="350" swimtime="00:04:55.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katharina" lastname="Szymańska" birthdate="1985-05-31" gender="F" nation="POL" athleteid="3033">
              <RESULTS>
                <RESULT eventid="1508" points="300" reactiontime="+93" swimtime="00:03:08.17" resultid="3034" heatid="4395" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:30.40" />
                    <SPLIT distance="150" swimtime="00:02:20.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1576" points="265" reactiontime="+96" swimtime="00:07:46.56" resultid="3035" heatid="4413" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.01" />
                    <SPLIT distance="150" swimtime="00:02:53.08" />
                    <SPLIT distance="200" swimtime="00:03:57.04" />
                    <SPLIT distance="250" swimtime="00:04:59.53" />
                    <SPLIT distance="300" swimtime="00:06:04.82" />
                    <SPLIT distance="350" swimtime="00:06:58.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="274" reactiontime="+95" swimtime="00:00:50.29" resultid="3036" heatid="4438" lane="3" />
                <RESULT eventid="1731" points="278" reactiontime="+94" swimtime="00:06:47.95" resultid="3037" heatid="4455" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                    <SPLIT distance="100" swimtime="00:01:36.07" />
                    <SPLIT distance="150" swimtime="00:02:27.28" />
                    <SPLIT distance="200" swimtime="00:03:20.29" />
                    <SPLIT distance="250" swimtime="00:04:12.64" />
                    <SPLIT distance="350" swimtime="00:05:59.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marlena" lastname="Dobrasiewicz-Iwaniuk" birthdate="1988-05-24" gender="F" nation="POL" athleteid="3045">
              <RESULTS>
                <RESULT eventid="1233" points="499" reactiontime="+89" swimtime="00:03:07.79" resultid="3046" heatid="4328" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:30.65" />
                    <SPLIT distance="150" swimtime="00:02:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="516" reactiontime="+87" swimtime="00:01:08.89" resultid="3047" heatid="4340" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="527" reactiontime="+90" swimtime="00:01:26.78" resultid="3048" heatid="4365" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="GALICA" birthdate="1985-11-25" gender="F" nation="POL" license="504214500057" athleteid="4243">
              <RESULTS>
                <RESULT eventid="1731" points="415" reactiontime="+77" swimtime="00:05:56.84" resultid="4244" heatid="4452" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="100" swimtime="00:01:17.29" />
                    <SPLIT distance="150" swimtime="00:02:02.82" />
                    <SPLIT distance="200" swimtime="00:02:49.00" />
                    <SPLIT distance="250" swimtime="00:03:35.81" />
                    <SPLIT distance="300" swimtime="00:04:23.04" />
                    <SPLIT distance="350" swimtime="00:05:10.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="4245" heatid="4397" lane="2" entrytime="00:03:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Saienko" birthdate="1994-08-03" gender="M" nation="UKR" athleteid="3038">
              <RESULTS>
                <RESULT eventid="1112" points="548" reactiontime="+79" swimtime="00:02:31.08" resultid="3039" heatid="4297" lane="9" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:54.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="669" reactiontime="+74" swimtime="00:00:57.67" resultid="3040" heatid="4351" lane="1" entrytime="00:00:57.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="625" reactiontime="+68" swimtime="00:02:09.56" resultid="3041" heatid="4406" lane="4" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                    <SPLIT distance="100" swimtime="00:01:02.17" />
                    <SPLIT distance="150" swimtime="00:01:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="570" reactiontime="+71" swimtime="00:01:04.02" resultid="3042" heatid="4426" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zenon" lastname="Kuliś" birthdate="1954-06-04" gender="M" nation="POL" athleteid="3007">
              <RESULTS>
                <RESULT eventid="1076" points="287" reactiontime="+122" swimtime="00:00:39.73" resultid="3008" heatid="4276" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1267" points="177" reactiontime="+93" swimtime="00:00:55.12" resultid="3009" heatid="4320" lane="4" entrytime="00:00:53.00" />
                <RESULT eventid="1301" points="259" reactiontime="+104" swimtime="00:01:33.38" resultid="3010" heatid="4344" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="3011" heatid="4462" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Skośkiewicz" birthdate="1966-05-05" gender="M" nation="POL" athleteid="2911">
              <RESULTS>
                <RESULT eventid="1076" points="648" reactiontime="+78" swimtime="00:00:28.25" resultid="2912" heatid="4281" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1112" points="701" reactiontime="+81" swimtime="00:02:38.37" resultid="2913" heatid="4296" lane="0" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:02:01.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="663" reactiontime="+74" swimtime="00:00:33.30" resultid="2914" heatid="4324" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1301" points="692" reactiontime="+86" swimtime="00:01:03.32" resultid="2915" heatid="4349" lane="9" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="703" reactiontime="+82" swimtime="00:00:29.87" resultid="2916" heatid="4381" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1491" points="677" reactiontime="+71" swimtime="00:01:12.30" resultid="2917" heatid="4393" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="655" reactiontime="+83" swimtime="00:01:09.74" resultid="2918" heatid="4425" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="630" reactiontime="+82" swimtime="00:02:44.29" resultid="2919" heatid="4436" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                    <SPLIT distance="150" swimtime="00:02:04.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Szymański" birthdate="1980-10-04" gender="M" nation="POL" athleteid="3028">
              <RESULTS>
                <RESULT eventid="1076" points="781" reactiontime="+73" swimtime="00:00:25.25" resultid="3029" heatid="4286" lane="1" entrytime="00:00:25.50" />
                <RESULT eventid="1267" points="822" reactiontime="+71" swimtime="00:00:28.96" resultid="3030" heatid="4325" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="3031" heatid="4384" lane="1" entrytime="00:00:27.30" />
                <RESULT eventid="1491" points="759" reactiontime="+73" swimtime="00:01:04.07" resultid="3032" heatid="4394" lane="3" entrytime="00:01:03.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Kośla" birthdate="1993-01-05" gender="F" nation="POL" athleteid="2971">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="2972" heatid="4271" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1215" points="608" reactiontime="+70" swimtime="00:00:33.52" resultid="2973" heatid="4316" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1474" points="575" reactiontime="+73" swimtime="00:01:14.09" resultid="2974" heatid="4388" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" status="DNS" swimtime="00:00:00.00" resultid="2975" heatid="4431" lane="4" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Sutowski" birthdate="1993-02-18" gender="M" nation="POL" athleteid="2938">
              <RESULTS>
                <RESULT eventid="1076" points="445" reactiontime="+75" swimtime="00:00:29.22" resultid="2939" heatid="4281" lane="7" entrytime="00:00:29.15" />
                <RESULT eventid="1301" points="424" reactiontime="+76" swimtime="00:01:07.14" resultid="2940" heatid="4347" lane="2" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="357" reactiontime="+70" swimtime="00:00:33.43" resultid="2941" heatid="4381" lane="9" entrytime="00:00:33.80" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="2942" heatid="4403" lane="2" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dymitr" lastname="Bielski" birthdate="1977-08-13" gender="M" nation="POL" athleteid="2925">
              <RESULTS>
                <RESULT eventid="1076" status="WDR" swimtime="00:00:00.00" resultid="2926" entrytime="00:00:30.00" />
                <RESULT eventid="1267" status="WDR" swimtime="00:00:00.00" resultid="2927" entrytime="00:00:37.00" />
                <RESULT eventid="1457" status="WDR" swimtime="00:00:00.00" resultid="2928" entrytime="00:00:33.00" />
                <RESULT eventid="1629" points="294" reactiontime="+85" swimtime="00:01:25.48" resultid="2929" heatid="4424" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="386" reactiontime="+82" swimtime="00:05:44.80" resultid="2930" heatid="4460" lane="3" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                    <SPLIT distance="200" swimtime="00:02:44.56" />
                    <SPLIT distance="250" swimtime="00:03:29.47" />
                    <SPLIT distance="300" swimtime="00:04:15.32" />
                    <SPLIT distance="350" swimtime="00:05:01.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luka" lastname="Crnjakovic" birthdate="1978-07-08" gender="M" nation="POL" athleteid="2943">
              <RESULTS>
                <RESULT eventid="1267" status="DNS" swimtime="00:00:00.00" resultid="2944" heatid="4323" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="2945" heatid="4405" lane="5" entrytime="00:02:18.00" />
                <RESULT eventid="1663" status="DNS" swimtime="00:00:00.00" resultid="2946" heatid="4436" lane="6" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Rogosz" birthdate="1976-04-28" gender="M" nation="POL" athleteid="2964">
              <RESULTS>
                <RESULT eventid="1112" points="522" reactiontime="+84" swimtime="00:02:41.53" resultid="2965" heatid="4295" lane="5" entrytime="00:02:41.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:02:41.53" />
                    <SPLIT distance="150" swimtime="00:02:05.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1197" points="489" reactiontime="+101" swimtime="00:21:07.98" resultid="2966" heatid="4309" lane="9" entrytime="00:22:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:18.72" />
                    <SPLIT distance="150" swimtime="00:02:01.94" />
                    <SPLIT distance="200" swimtime="00:02:44.27" />
                    <SPLIT distance="250" swimtime="00:03:26.94" />
                    <SPLIT distance="300" swimtime="00:04:10.02" />
                    <SPLIT distance="350" swimtime="00:04:52.36" />
                    <SPLIT distance="400" swimtime="00:05:35.19" />
                    <SPLIT distance="450" swimtime="00:06:17.36" />
                    <SPLIT distance="500" swimtime="00:06:59.65" />
                    <SPLIT distance="550" swimtime="00:07:42.39" />
                    <SPLIT distance="600" swimtime="00:08:24.82" />
                    <SPLIT distance="650" swimtime="00:09:06.94" />
                    <SPLIT distance="700" swimtime="00:09:49.03" />
                    <SPLIT distance="750" swimtime="00:10:31.53" />
                    <SPLIT distance="800" swimtime="00:11:13.92" />
                    <SPLIT distance="850" swimtime="00:11:56.49" />
                    <SPLIT distance="900" swimtime="00:12:39.02" />
                    <SPLIT distance="950" swimtime="00:13:21.82" />
                    <SPLIT distance="1000" swimtime="00:14:04.07" />
                    <SPLIT distance="1050" swimtime="00:14:47.12" />
                    <SPLIT distance="1100" swimtime="00:15:29.71" />
                    <SPLIT distance="1150" swimtime="00:16:12.21" />
                    <SPLIT distance="1200" swimtime="00:16:55.39" />
                    <SPLIT distance="1250" swimtime="00:17:38.10" />
                    <SPLIT distance="1300" swimtime="00:18:21.06" />
                    <SPLIT distance="1350" swimtime="00:19:03.69" />
                    <SPLIT distance="1400" swimtime="00:19:45.87" />
                    <SPLIT distance="1450" swimtime="00:20:27.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="504" reactiontime="+99" swimtime="00:02:55.23" resultid="2967" heatid="4333" lane="3" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="150" swimtime="00:02:11.27" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G4" eventid="1593" reactiontime="+81" status="DSQ" swimtime="00:00:00.00" resultid="2968" heatid="4414" lane="9" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:20.68" />
                    <SPLIT distance="150" swimtime="00:02:09.14" />
                    <SPLIT distance="200" swimtime="00:02:56.61" />
                    <SPLIT distance="250" swimtime="00:03:42.32" />
                    <SPLIT distance="300" swimtime="00:04:29.51" />
                    <SPLIT distance="350" swimtime="00:05:08.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="417" reactiontime="+92" swimtime="00:01:16.12" resultid="2969" heatid="4424" lane="5" entrytime="00:01:17.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="2970" heatid="4458" lane="9" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Szemberg" birthdate="1949-07-26" gender="F" nation="POL" athleteid="2995">
              <RESULTS>
                <RESULT eventid="1059" points="138" swimtime="00:00:59.46" resultid="2996" heatid="4268" lane="5" entrytime="00:00:57.00" />
                <RESULT eventid="1180" points="217" swimtime="00:37:06.22" resultid="2997" heatid="4308" lane="2" entrytime="00:38:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.31" />
                    <SPLIT distance="100" swimtime="00:02:20.44" />
                    <SPLIT distance="150" swimtime="00:03:36.44" />
                    <SPLIT distance="200" swimtime="00:04:49.07" />
                    <SPLIT distance="250" swimtime="00:06:03.23" />
                    <SPLIT distance="300" swimtime="00:07:17.61" />
                    <SPLIT distance="350" swimtime="00:08:32.80" />
                    <SPLIT distance="400" swimtime="00:09:46.98" />
                    <SPLIT distance="450" swimtime="00:11:01.85" />
                    <SPLIT distance="500" swimtime="00:12:16.35" />
                    <SPLIT distance="550" swimtime="00:13:30.04" />
                    <SPLIT distance="600" swimtime="00:14:44.92" />
                    <SPLIT distance="650" swimtime="00:15:59.51" />
                    <SPLIT distance="700" swimtime="00:17:13.78" />
                    <SPLIT distance="750" swimtime="00:18:28.26" />
                    <SPLIT distance="800" swimtime="00:19:42.50" />
                    <SPLIT distance="850" swimtime="00:20:57.96" />
                    <SPLIT distance="900" swimtime="00:22:12.81" />
                    <SPLIT distance="950" swimtime="00:23:27.78" />
                    <SPLIT distance="1000" swimtime="00:24:42.50" />
                    <SPLIT distance="1050" swimtime="00:25:58.13" />
                    <SPLIT distance="1100" swimtime="00:27:13.14" />
                    <SPLIT distance="1150" swimtime="00:28:28.70" />
                    <SPLIT distance="1200" swimtime="00:29:42.26" />
                    <SPLIT distance="1250" swimtime="00:30:57.42" />
                    <SPLIT distance="1300" swimtime="00:32:12.68" />
                    <SPLIT distance="1350" swimtime="00:33:26.71" />
                    <SPLIT distance="1400" swimtime="00:34:41.17" />
                    <SPLIT distance="1450" swimtime="00:35:54.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="122" swimtime="00:02:14.75" resultid="2998" heatid="4337" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="183" swimtime="00:09:32.79" resultid="2999" heatid="4454" lane="8" entrytime="00:09:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.97" />
                    <SPLIT distance="100" swimtime="00:02:16.67" />
                    <SPLIT distance="150" swimtime="00:03:29.92" />
                    <SPLIT distance="200" swimtime="00:04:43.12" />
                    <SPLIT distance="250" swimtime="00:05:56.48" />
                    <SPLIT distance="300" swimtime="00:07:10.15" />
                    <SPLIT distance="350" swimtime="00:08:23.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Olszewska" birthdate="1964-08-01" gender="F" nation="POL" athleteid="3018">
              <RESULTS>
                <RESULT eventid="1233" status="WDR" swimtime="00:00:00.00" resultid="3019" entrytime="00:03:40.00" />
                <RESULT eventid="1404" status="WDR" swimtime="00:00:00.00" resultid="3020" entrytime="00:01:44.00" />
                <RESULT eventid="1474" points="78" swimtime="00:02:42.87" resultid="3021" heatid="4387" lane="7" entrytime="00:01:56.00" />
                <RESULT eventid="1680" status="WDR" swimtime="00:00:00.00" resultid="3022" heatid="4440" lane="7" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Warchoł" birthdate="1953-08-30" gender="M" nation="POL" athleteid="2920">
              <RESULTS>
                <RESULT eventid="1076" points="554" reactiontime="+85" swimtime="00:00:31.92" resultid="2921" heatid="4279" lane="2" entrytime="00:00:31.55" />
                <RESULT eventid="1301" points="595" reactiontime="+87" swimtime="00:01:10.72" resultid="2922" heatid="4347" lane="7" entrytime="00:01:09.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="636" reactiontime="+81" swimtime="00:01:21.14" resultid="2923" heatid="4392" lane="2" entrytime="00:01:22.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="716" reactiontime="+81" swimtime="00:02:55.67" resultid="2924" heatid="4435" lane="5" entrytime="00:02:54.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:25.78" />
                    <SPLIT distance="150" swimtime="00:02:11.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1386" points="704" reactiontime="+64" swimtime="00:01:55.01" resultid="3051" heatid="4493" lane="3" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:00.99" />
                    <SPLIT distance="150" swimtime="00:01:28.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3028" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="3000" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3038" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3023" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1386" points="580" reactiontime="+79" swimtime="00:02:06.46" resultid="3052" heatid="4493" lane="8" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:07.17" />
                    <SPLIT distance="150" swimtime="00:01:37.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2911" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2983" number="2" />
                    <RELAYPOSITION athleteid="2954" number="3" reactiontime="+8" />
                    <RELAYPOSITION athleteid="2938" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1386" points="440" reactiontime="+80" swimtime="00:02:25.69" resultid="3053" heatid="4492" lane="5" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="150" swimtime="00:01:57.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2920" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2931" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="2947" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="2959" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="1559" points="746" reactiontime="+74" swimtime="00:01:42.38" resultid="3055" heatid="4497" lane="4" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.18" />
                    <SPLIT distance="100" swimtime="00:00:51.50" />
                    <SPLIT distance="150" swimtime="00:01:17.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3028" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="3023" number="2" />
                    <RELAYPOSITION athleteid="3000" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="3038" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1559" points="522" reactiontime="+83" swimtime="00:01:55.27" resultid="3056" heatid="4497" lane="1" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="100" swimtime="00:00:58.80" />
                    <SPLIT distance="150" swimtime="00:01:27.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2938" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2983" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="2959" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="2931" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="1559" points="549" reactiontime="+83" swimtime="00:01:59.97" resultid="3057" heatid="4497" lane="9" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                    <SPLIT distance="100" swimtime="00:00:59.34" />
                    <SPLIT distance="150" swimtime="00:01:28.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2954" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2925" number="2" />
                    <RELAYPOSITION athleteid="2911" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2920" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="2">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1369" points="706" reactiontime="+72" swimtime="00:02:17.39" resultid="3050" heatid="4490" lane="5" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:14.74" />
                    <SPLIT distance="150" swimtime="00:01:46.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2971" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="3043" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2976" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="3045" number="4" reactiontime="+77" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="6">
              <RESULTS>
                <RESULT eventid="1542" points="697" reactiontime="+75" swimtime="00:02:02.99" resultid="3054" heatid="4494" lane="5" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="100" swimtime="00:01:00.76" />
                    <SPLIT distance="150" swimtime="00:01:33.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2971" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3045" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3043" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="2976" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" points="730" reactiontime="+71" swimtime="00:01:51.20" resultid="3049" heatid="4489" lane="4" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.16" />
                    <SPLIT distance="100" swimtime="00:00:54.12" />
                    <SPLIT distance="150" swimtime="00:01:24.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3028" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="2976" number="2" />
                    <RELAYPOSITION athleteid="2971" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="3038" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="10">
              <RESULTS>
                <RESULT eventid="1714" points="722" reactiontime="+69" swimtime="00:02:03.49" resultid="3058" heatid="4499" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                    <SPLIT distance="100" swimtime="00:01:01.53" />
                    <SPLIT distance="150" swimtime="00:01:34.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3028" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3038" number="2" />
                    <RELAYPOSITION athleteid="2971" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2976" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="11">
              <RESULTS>
                <RESULT eventid="1714" reactiontime="+68" status="DSQ" swimtime="00:00:00.00" resultid="3059" heatid="4499" lane="2" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:11.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2931" number="1" reactiontime="+68" status="DSQ" />
                    <RELAYPOSITION athleteid="3000" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2987" number="3" reactiontime="+104" status="DSQ" />
                    <RELAYPOSITION athleteid="3033" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3208" name="Swim Tri Rzeszów">
          <CONTACT name="SWIM TRI RZESZÓW" />
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Sarna" birthdate="1975-10-31" gender="M" nation="POL" athleteid="3215">
              <RESULTS>
                <RESULT eventid="1076" points="617" reactiontime="+73" swimtime="00:00:27.67" resultid="3216" heatid="4285" lane="2" entrytime="00:00:26.44" />
                <RESULT eventid="1301" points="589" reactiontime="+71" swimtime="00:01:02.33" resultid="3217" heatid="4350" lane="6" entrytime="00:00:59.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="652" reactiontime="+74" swimtime="00:02:15.80" resultid="3218" heatid="4406" lane="2" entrytime="00:02:11.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:05.45" />
                    <SPLIT distance="150" swimtime="00:01:41.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="621" reactiontime="+80" swimtime="00:04:54.23" resultid="3219" heatid="4456" lane="9" entrytime="00:04:44.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:06.67" />
                    <SPLIT distance="150" swimtime="00:01:43.50" />
                    <SPLIT distance="200" swimtime="00:02:21.27" />
                    <SPLIT distance="250" swimtime="00:02:59.67" />
                    <SPLIT distance="300" swimtime="00:03:38.34" />
                    <SPLIT distance="350" swimtime="00:04:17.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Faff" birthdate="1963-11-15" gender="M" nation="POL" athleteid="3209">
              <RESULTS>
                <RESULT eventid="1076" points="600" reactiontime="+78" swimtime="00:00:28.99" resultid="3210" heatid="4282" lane="1" entrytime="00:00:28.28" />
                <RESULT eventid="1301" points="610" reactiontime="+76" swimtime="00:01:06.03" resultid="3211" heatid="4348" lane="8" entrytime="00:01:05.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="569" reactiontime="+84" swimtime="00:00:32.06" resultid="3212" heatid="4381" lane="8" entrytime="00:00:32.25" />
                <RESULT eventid="1525" points="543" reactiontime="+82" swimtime="00:02:32.04" resultid="3213" heatid="4404" lane="2" entrytime="00:02:26.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:52.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="491" reactiontime="+82" swimtime="00:05:32.80" resultid="3214" heatid="4458" lane="0" entrytime="00:05:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:56.12" />
                    <SPLIT distance="100" swimtime="00:01:13.37" />
                    <SPLIT distance="200" swimtime="00:02:40.11" />
                    <SPLIT distance="300" swimtime="00:04:07.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04002" nation="POL" region="02" clubid="2461" name="Stowarzyszenie AZS WSG">
          <ATHLETES>
            <ATHLETE firstname="Kinga" lastname="Paradowska" birthdate="2001-06-12" gender="F" nation="POL" license="104002600006" swrid="4411672" athleteid="2462">
              <RESULTS>
                <RESULT eventid="1094" reactiontime="+71" swimtime="00:02:26.59" resultid="2463" heatid="4290" lane="4" entrytime="00:02:19.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:11.75" />
                    <SPLIT distance="150" swimtime="00:01:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" reactiontime="+72" swimtime="00:09:22.04" resultid="2464" heatid="4300" lane="4" entrytime="00:09:10.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:10.05" />
                    <SPLIT distance="150" swimtime="00:01:46.15" />
                    <SPLIT distance="200" swimtime="00:02:22.61" />
                    <SPLIT distance="250" swimtime="00:02:58.63" />
                    <SPLIT distance="300" swimtime="00:03:34.63" />
                    <SPLIT distance="350" swimtime="00:04:10.30" />
                    <SPLIT distance="400" swimtime="00:04:46.33" />
                    <SPLIT distance="450" swimtime="00:05:21.20" />
                    <SPLIT distance="500" swimtime="00:05:56.46" />
                    <SPLIT distance="550" swimtime="00:06:31.35" />
                    <SPLIT distance="600" swimtime="00:07:06.40" />
                    <SPLIT distance="650" swimtime="00:07:40.88" />
                    <SPLIT distance="700" swimtime="00:08:15.73" />
                    <SPLIT distance="750" swimtime="00:08:48.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" reactiontime="+69" swimtime="00:02:44.94" resultid="2465" heatid="4328" lane="4" entrytime="00:02:33.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:20.36" />
                    <SPLIT distance="150" swimtime="00:02:03.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1335" reactiontime="+69" swimtime="00:02:23.12" resultid="2466" heatid="4354" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:10.15" />
                    <SPLIT distance="150" swimtime="00:01:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" reactiontime="+67" swimtime="00:01:18.86" resultid="2467" heatid="4365" lane="4" entrytime="00:01:13.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1576" reactiontime="+69" swimtime="00:05:22.10" resultid="2468" heatid="4412" lane="4" entrytime="00:04:54.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="150" swimtime="00:01:54.40" />
                    <SPLIT distance="200" swimtime="00:02:34.41" />
                    <SPLIT distance="250" swimtime="00:03:20.80" />
                    <SPLIT distance="300" swimtime="00:04:05.83" />
                    <SPLIT distance="350" swimtime="00:04:44.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" reactiontime="+69" swimtime="00:01:05.41" resultid="2469" heatid="4421" lane="5" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" reactiontime="+70" swimtime="00:04:35.08" resultid="2470" heatid="4452" lane="4" entrytime="00:04:31.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="150" swimtime="00:01:43.03" />
                    <SPLIT distance="200" swimtime="00:02:18.38" />
                    <SPLIT distance="250" swimtime="00:02:52.98" />
                    <SPLIT distance="300" swimtime="00:03:28.05" />
                    <SPLIT distance="350" swimtime="00:04:02.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrianna" lastname="Rzewuska" birthdate="1997-05-30" gender="F" nation="POL" license="504002600005" swrid="4261695" athleteid="2471">
              <RESULTS>
                <RESULT eventid="1215" points="552" reactiontime="+71" swimtime="00:00:34.60" resultid="2472" heatid="4312" lane="0" />
                <RESULT comment="G1" eventid="1474" reactiontime="+82" status="DSQ" swimtime="00:00:00.00" resultid="2473" heatid="4386" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="495" reactiontime="+75" swimtime="00:02:48.32" resultid="2474" heatid="4429" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:01:20.27" />
                    <SPLIT distance="150" swimtime="00:02:04.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Rutkowska" birthdate="1999-06-10" gender="F" nation="POL" license="104002600004" swrid="4411705" athleteid="2475">
              <RESULTS>
                <RESULT eventid="1335" reactiontime="+78" swimtime="00:02:35.08" resultid="2476" heatid="4353" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:12.47" />
                    <SPLIT distance="150" swimtime="00:01:53.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" reactiontime="+76" swimtime="00:02:40.92" resultid="2477" heatid="4429" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:18.12" />
                    <SPLIT distance="150" swimtime="00:01:59.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4025">
          <ATHLETES>
            <ATHLETE firstname="Aleksandra" lastname="CWOJDZIŃSKA" birthdate="1992-12-21" gender="F" nation="POL" swrid="4104697" athleteid="4261">
              <RESULTS>
                <RESULT eventid="1059" points="430" reactiontime="+67" swimtime="00:00:34.09" resultid="4262" heatid="4270" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1215" points="406" reactiontime="+68" swimtime="00:00:38.59" resultid="4263" heatid="4315" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1474" points="396" reactiontime="+61" swimtime="00:01:24.15" resultid="4264" heatid="4387" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="377" reactiontime="+71" swimtime="00:03:10.53" resultid="4265" heatid="4430" lane="4" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                    <SPLIT distance="150" swimtime="00:02:20.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="WIESŁAW" lastname="CIEKLIŃSKI" birthdate="1957-01-01" gender="M" nation="POL" athleteid="3751">
              <RESULTS>
                <RESULT eventid="1076" points="519" reactiontime="+90" swimtime="00:00:32.61" resultid="3752" heatid="4278" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1197" points="447" reactiontime="+87" swimtime="00:25:34.34" resultid="3753" heatid="4311" lane="8" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:30.00" />
                    <SPLIT distance="150" swimtime="00:02:19.79" />
                    <SPLIT distance="200" swimtime="00:03:09.85" />
                    <SPLIT distance="250" swimtime="00:04:01.35" />
                    <SPLIT distance="300" swimtime="00:06:36.63" />
                    <SPLIT distance="350" swimtime="00:05:44.43" />
                    <SPLIT distance="400" swimtime="00:11:48.00" />
                    <SPLIT distance="450" swimtime="00:07:28.48" />
                    <SPLIT distance="550" swimtime="00:09:12.06" />
                    <SPLIT distance="650" swimtime="00:10:56.97" />
                    <SPLIT distance="750" swimtime="00:12:38.80" />
                    <SPLIT distance="800" swimtime="00:15:13.45" />
                    <SPLIT distance="850" swimtime="00:14:22.88" />
                    <SPLIT distance="900" swimtime="00:16:55.45" />
                    <SPLIT distance="950" swimtime="00:16:03.54" />
                    <SPLIT distance="1000" swimtime="00:18:43.63" />
                    <SPLIT distance="1050" swimtime="00:19:36.51" />
                    <SPLIT distance="1100" swimtime="00:20:27.54" />
                    <SPLIT distance="1150" swimtime="00:21:19.04" />
                    <SPLIT distance="1200" swimtime="00:22:13.84" />
                    <SPLIT distance="1250" swimtime="00:23:06.42" />
                    <SPLIT distance="1300" swimtime="00:25:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="536" reactiontime="+88" swimtime="00:01:13.22" resultid="3754" heatid="4346" lane="7" entrytime="00:01:13.90" />
                <RESULT eventid="1525" points="426" reactiontime="+81" swimtime="00:02:52.00" resultid="3755" heatid="4402" lane="5" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                    <SPLIT distance="100" swimtime="00:01:23.00" />
                    <SPLIT distance="150" swimtime="00:02:10.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="367" reactiontime="+89" swimtime="00:06:27.93" resultid="3756" heatid="4460" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.87" />
                    <SPLIT distance="100" swimtime="00:01:28.41" />
                    <SPLIT distance="150" swimtime="00:02:19.21" />
                    <SPLIT distance="200" swimtime="00:03:11.99" />
                    <SPLIT distance="250" swimtime="00:04:03.39" />
                    <SPLIT distance="300" swimtime="00:04:54.20" />
                    <SPLIT distance="350" swimtime="00:05:44.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="ROBERT" lastname="KAMIŃSKI" birthdate="1965-01-01" gender="M" nation="POL" athleteid="3947" />
            <ATHLETE firstname="IZABELA" lastname="WYPYCH-STASZEWSKA" birthdate="1970-01-01" gender="F" nation="POL" athleteid="3837">
              <RESULTS>
                <RESULT eventid="1059" points="416" reactiontime="+69" swimtime="00:00:36.29" resultid="3838" heatid="4269" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1284" points="403" reactiontime="+72" swimtime="00:01:21.82" resultid="3839" heatid="4339" lane="9" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="407" reactiontime="+70" swimtime="00:00:40.23" resultid="3840" heatid="4373" lane="4" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="ALINA" lastname="PIEKARSKA" birthdate="1947-01-01" gender="F" nation="POL" athleteid="3993">
              <RESULTS>
                <RESULT eventid="1680" points="30" swimtime="00:02:21.54" resultid="3994" heatid="4439" lane="1" entrytime="00:02:11.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="WIKTOR" lastname="WIŚNIEWSKI" birthdate="1995-01-01" gender="M" nation="POL" athleteid="3861">
              <RESULTS>
                <RESULT eventid="1267" points="590" reactiontime="+77" swimtime="00:00:30.33" resultid="3862" heatid="4323" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1491" points="550" reactiontime="+79" swimtime="00:01:07.22" resultid="3863" heatid="4394" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="518" reactiontime="+77" swimtime="00:02:32.81" resultid="3864" heatid="4435" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:52.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="TOBIASZ" lastname="JANKOWSKI" birthdate="1983-01-01" gender="M" nation="POL" athleteid="3908">
              <RESULTS>
                <RESULT comment="Z3G8" eventid="1112" reactiontime="+73" status="DSQ" swimtime="00:00:00.00" resultid="3909" heatid="4294" lane="6" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="376" reactiontime="+75" swimtime="00:01:26.46" resultid="3910" heatid="4369" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="366" reactiontime="+68" swimtime="00:00:33.76" resultid="3911" heatid="4380" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1697" points="447" reactiontime="+71" swimtime="00:00:37.24" resultid="3912" heatid="4446" lane="0" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="MACIEJ" lastname="KORZUCHOWSKI" birthdate="1999-01-01" gender="M" nation="POL" swrid="4598470" athleteid="3937">
              <RESULTS>
                <RESULT eventid="1112" reactiontime="+79" swimtime="00:02:47.47" resultid="3940" heatid="4296" lane="8" entrytime="00:02:38.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="150" swimtime="00:02:09.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" status="DNS" swimtime="00:00:00.00" resultid="3941" heatid="4325" lane="0" entrytime="00:00:31.27" />
                <RESULT eventid="1250" status="DNS" swimtime="00:00:00.00" resultid="3942" heatid="4332" lane="5" entrytime="00:03:00.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3943" heatid="4394" lane="1" entrytime="00:01:09.00" />
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="3944" heatid="4415" lane="4" entrytime="00:05:45.00" />
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="3945" heatid="4426" lane="8" entrytime="00:01:07.42" />
                <RESULT eventid="1663" status="DNS" swimtime="00:00:00.00" resultid="3946" heatid="4436" lane="4" entrytime="00:02:37.00" />
                <RESULT eventid="1076" reactiontime="+67" swimtime="00:00:27.27" resultid="4119" heatid="4283" lane="5" entrytime="00:00:27.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="DOMINIKA" lastname="OPAŁKO" birthdate="1999-01-01" gender="F" nation="POL" swrid="4493246" athleteid="3852">
              <RESULTS>
                <RESULT eventid="1094" reactiontime="+78" swimtime="00:02:56.58" resultid="3853" heatid="4290" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                    <SPLIT distance="150" swimtime="00:02:12.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" reactiontime="+83" swimtime="00:03:27.38" resultid="3855" heatid="4328" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                    <SPLIT distance="100" swimtime="00:01:37.95" />
                    <SPLIT distance="150" swimtime="00:02:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1335" reactiontime="+86" swimtime="00:03:27.72" resultid="3856" heatid="4354" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:01:32.48" />
                    <SPLIT distance="150" swimtime="00:02:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="3857" heatid="4374" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1576" status="DNS" swimtime="00:00:00.00" resultid="3858" heatid="4412" lane="3" entrytime="00:06:00.00" />
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="3859" heatid="4421" lane="9" entrytime="00:01:23.00" />
                <RESULT eventid="1646" status="DNS" swimtime="00:00:00.00" resultid="3860" heatid="4431" lane="7" entrytime="00:03:05.00" />
                <RESULT eventid="1059" reactiontime="+73" swimtime="00:00:30.98" resultid="4194" heatid="4271" lane="5" entrytime="00:00:30.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="PRZEMYSŁAW" lastname="KUŚMIDER" birthdate="1989-01-01" gender="M" nation="POL" athleteid="3777">
              <RESULTS>
                <RESULT eventid="1076" points="459" reactiontime="+79" swimtime="00:00:28.68" resultid="3778" heatid="4280" lane="4" entrytime="00:00:29.90" />
                <RESULT eventid="1163" points="441" reactiontime="+90" swimtime="00:10:41.77" resultid="3779" heatid="4304" lane="1" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:52.86" />
                    <SPLIT distance="200" swimtime="00:02:32.81" />
                    <SPLIT distance="250" swimtime="00:03:13.55" />
                    <SPLIT distance="300" swimtime="00:03:54.58" />
                    <SPLIT distance="350" swimtime="00:04:35.25" />
                    <SPLIT distance="400" swimtime="00:05:15.84" />
                    <SPLIT distance="450" swimtime="00:05:56.12" />
                    <SPLIT distance="500" swimtime="00:06:37.32" />
                    <SPLIT distance="550" swimtime="00:07:18.20" />
                    <SPLIT distance="600" swimtime="00:07:59.25" />
                    <SPLIT distance="650" swimtime="00:08:40.29" />
                    <SPLIT distance="700" swimtime="00:09:21.88" />
                    <SPLIT distance="750" swimtime="00:10:02.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="445" reactiontime="+90" swimtime="00:01:05.21" resultid="3780" heatid="4348" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="456" reactiontime="+78" swimtime="00:02:22.30" resultid="3781" heatid="4404" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="150" swimtime="00:01:46.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="IZABELA" lastname="SKURCZYŃSKA" birthdate="1971-01-01" gender="F" nation="POL" athleteid="3810">
              <RESULTS>
                <RESULT eventid="1059" points="241" reactiontime="+88" swimtime="00:00:43.53" resultid="3811" heatid="4269" lane="9" entrytime="00:00:46.50" />
                <RESULT eventid="1404" points="283" reactiontime="+86" swimtime="00:01:54.94" resultid="3812" heatid="4364" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="156" reactiontime="+82" swimtime="00:00:55.37" resultid="3813" heatid="4372" lane="3" />
                <RESULT eventid="1680" points="284" reactiontime="+82" swimtime="00:00:52.01" resultid="3814" heatid="4440" lane="8" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="RAFAŁ" lastname="SZKLARZEWSKI" birthdate="1985-01-01" gender="M" nation="POL" athleteid="3841">
              <RESULTS>
                <RESULT eventid="1076" points="555" reactiontime="+59" swimtime="00:00:27.69" resultid="3842" heatid="4285" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="3843" heatid="4305" lane="5" entrytime="00:12:00.00" />
                <RESULT eventid="1301" points="527" reactiontime="+64" swimtime="00:01:02.85" resultid="3844" heatid="4350" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="422" reactiontime="+64" swimtime="00:00:32.19" resultid="3845" heatid="4383" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="3846" heatid="4405" lane="2" entrytime="00:02:20.00" />
                <RESULT eventid="1352" status="DNS" swimtime="00:00:00.00" resultid="3948" heatid="4357" lane="0" entrytime="00:02:50.00" />
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="3949" heatid="4425" lane="9" entrytime="00:01:15.00" />
                <RESULT eventid="1697" points="360" reactiontime="+63" swimtime="00:00:40.02" resultid="3950" heatid="4446" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1267" points="303" reactiontime="+61" swimtime="00:00:39.33" resultid="4242" heatid="4319" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="MICHAŁ" lastname="ANZORGE " birthdate="1982-01-01" gender="M" nation="POL" athleteid="3764">
              <RESULTS>
                <RESULT eventid="1076" points="427" reactiontime="+86" swimtime="00:00:30.88" resultid="3765" heatid="4285" lane="0" entrytime="00:00:26.60" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="3766" heatid="4351" lane="9" entrytime="00:00:58.70" />
                <RESULT eventid="1406" points="419" reactiontime="+77" swimtime="00:01:24.97" resultid="3767" heatid="4371" lane="7" entrytime="00:01:10.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="519" reactiontime="+71" swimtime="00:00:35.88" resultid="3768" heatid="4449" lane="7" entrytime="00:00:31.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="KAMIL" lastname="LUBIŃSKI" birthdate="1992-01-01" gender="M" nation="POL" athleteid="3961">
              <RESULTS>
                <RESULT eventid="1267" points="415" reactiontime="+89" swimtime="00:00:34.83" resultid="3962" heatid="4325" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1250" points="446" reactiontime="+84" swimtime="00:03:00.69" resultid="3963" heatid="4333" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:01:28.01" />
                    <SPLIT distance="150" swimtime="00:02:15.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="476" reactiontime="+76" swimtime="00:00:28.35" resultid="3966" heatid="4283" lane="3" entrytime="00:00:27.50" />
                <RESULT eventid="1163" points="361" reactiontime="+90" swimtime="00:11:26.02" resultid="3968" heatid="4304" lane="7" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:17.41" />
                    <SPLIT distance="150" swimtime="00:01:58.22" />
                    <SPLIT distance="200" swimtime="00:02:39.27" />
                    <SPLIT distance="250" swimtime="00:03:20.84" />
                    <SPLIT distance="300" swimtime="00:04:02.88" />
                    <SPLIT distance="350" swimtime="00:04:45.18" />
                    <SPLIT distance="400" swimtime="00:05:28.58" />
                    <SPLIT distance="450" swimtime="00:06:12.23" />
                    <SPLIT distance="500" swimtime="00:06:56.02" />
                    <SPLIT distance="550" swimtime="00:07:40.50" />
                    <SPLIT distance="650" swimtime="00:09:11.59" />
                    <SPLIT distance="750" swimtime="00:10:42.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="3969" heatid="4370" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1663" points="375" reactiontime="+89" swimtime="00:02:50.15" resultid="3970" heatid="4436" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                    <SPLIT distance="150" swimtime="00:02:08.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="414" reactiontime="+82" swimtime="00:05:19.55" resultid="3971" heatid="4458" lane="7" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                    <SPLIT distance="150" swimtime="00:01:53.07" />
                    <SPLIT distance="200" swimtime="00:02:33.50" />
                    <SPLIT distance="250" swimtime="00:03:14.06" />
                    <SPLIT distance="300" swimtime="00:05:19.55" />
                    <SPLIT distance="350" swimtime="00:04:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="383" reactiontime="+82" swimtime="00:05:59.16" resultid="4049" heatid="4415" lane="6" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                    <SPLIT distance="150" swimtime="00:02:05.39" />
                    <SPLIT distance="200" swimtime="00:02:54.32" />
                    <SPLIT distance="250" swimtime="00:03:45.29" />
                    <SPLIT distance="300" swimtime="00:04:36.44" />
                    <SPLIT distance="350" swimtime="00:05:18.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="JANUSZ" lastname="PŁONKA" birthdate="1948-01-01" gender="M" nation="POL" swrid="4754750" athleteid="3954">
              <RESULTS>
                <RESULT eventid="1112" points="117" reactiontime="+105" swimtime="00:05:33.01" resultid="3955" heatid="4292" lane="7" entrytime="00:05:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.21" />
                    <SPLIT distance="100" swimtime="00:02:48.52" />
                    <SPLIT distance="150" swimtime="00:04:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="120" reactiontime="+108" swimtime="00:06:14.62" resultid="3956" heatid="4330" lane="5" entrytime="00:05:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.64" />
                    <SPLIT distance="100" swimtime="00:03:02.81" />
                    <SPLIT distance="150" swimtime="00:04:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="76" reactiontime="+114" swimtime="00:06:33.80" resultid="3957" heatid="4355" lane="1" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.81" />
                    <SPLIT distance="100" swimtime="00:03:13.59" />
                    <SPLIT distance="150" swimtime="00:04:59.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="87" reactiontime="+102" swimtime="00:11:24.13" resultid="3958" heatid="4462" lane="4" entrytime="00:09:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.77" />
                    <SPLIT distance="100" swimtime="00:02:43.10" />
                    <SPLIT distance="150" swimtime="00:04:14.62" />
                    <SPLIT distance="200" swimtime="00:05:44.23" />
                    <SPLIT distance="250" swimtime="00:07:12.22" />
                    <SPLIT distance="300" swimtime="00:08:37.86" />
                    <SPLIT distance="350" swimtime="00:10:03.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="51" reactiontime="+116" swimtime="00:03:01.54" resultid="3959" heatid="4423" lane="8" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="103" reactiontime="+102" swimtime="00:12:38.39" resultid="3960" heatid="4417" lane="5" entrytime="00:10:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.08" />
                    <SPLIT distance="100" swimtime="00:03:00.56" />
                    <SPLIT distance="150" swimtime="00:04:51.80" />
                    <SPLIT distance="200" swimtime="00:06:29.06" />
                    <SPLIT distance="250" swimtime="00:08:15.97" />
                    <SPLIT distance="300" swimtime="00:09:58.87" />
                    <SPLIT distance="350" swimtime="00:11:21.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="74" reactiontime="+103" swimtime="00:01:11.29" resultid="4250" heatid="4378" lane="7" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="MONIKA" lastname="BORUCH" birthdate="1978-01-01" gender="F" nation="POL" athleteid="3799">
              <RESULTS>
                <RESULT eventid="1284" points="332" reactiontime="+79" swimtime="00:01:23.84" resultid="3800" heatid="4338" lane="9" entrytime="00:01:25.80" />
                <RESULT eventid="1440" points="333" reactiontime="+83" swimtime="00:00:40.92" resultid="3801" heatid="4373" lane="6" entrytime="00:00:42.43" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="3802" heatid="4397" lane="9" entrytime="00:03:18.90" />
                <RESULT eventid="1611" points="172" reactiontime="+71" swimtime="00:01:53.85" resultid="3803" heatid="4420" lane="8" entrytime="00:01:57.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="ADAM" lastname="ZIELEZIŃSKI" birthdate="1951-01-01" gender="M" nation="POL" athleteid="3830">
              <RESULTS>
                <RESULT eventid="1076" points="219" swimtime="00:00:45.97" resultid="3831" heatid="4276" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="1112" points="180" reactiontime="+119" swimtime="00:04:48.42" resultid="3832" heatid="4293" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.35" />
                    <SPLIT distance="150" swimtime="00:03:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="79" swimtime="00:01:18.40" resultid="3833" heatid="4320" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="3834" heatid="4344" lane="8" entrytime="00:01:50.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="3835" heatid="4378" lane="6" entrytime="00:00:59.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3836" heatid="4390" lane="3" entrytime="00:01:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="KRZYSZTOF" lastname="KUBIAK" birthdate="1989-01-01" gender="M" nation="POL" athleteid="3790">
              <RESULTS>
                <RESULT comment="Z3G8" eventid="1112" status="DSQ" swimtime="00:00:00.00" resultid="3791" heatid="4294" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.15" />
                    <SPLIT distance="100" swimtime="00:01:54.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="3792" heatid="4304" lane="9" entrytime="00:11:10.00" />
                <RESULT eventid="1250" points="149" reactiontime="+105" swimtime="00:04:20.28" resultid="3793" heatid="4331" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.89" />
                    <SPLIT distance="100" swimtime="00:02:08.32" />
                    <SPLIT distance="150" swimtime="00:03:14.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="133" reactiontime="+117" swimtime="00:04:01.69" resultid="3794" heatid="4356" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.41" />
                    <SPLIT distance="100" swimtime="00:01:54.60" />
                    <SPLIT distance="150" swimtime="00:02:57.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="122" reactiontime="+91" swimtime="00:00:46.95" resultid="3795" heatid="4380" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1593" points="179" swimtime="00:07:42.75" resultid="3796" heatid="4415" lane="0" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:05:10.83" />
                    <SPLIT distance="100" swimtime="00:01:58.77" />
                    <SPLIT distance="200" swimtime="00:04:05.08" />
                    <SPLIT distance="300" swimtime="00:06:15.94" />
                    <SPLIT distance="350" swimtime="00:06:58.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="97" swimtime="00:01:56.74" resultid="3797" heatid="4424" lane="2" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="295" swimtime="00:05:57.64" resultid="3798" heatid="4459" lane="7" entrytime="00:05:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:01:23.70" />
                    <SPLIT distance="150" swimtime="00:02:09.28" />
                    <SPLIT distance="200" swimtime="00:02:55.33" />
                    <SPLIT distance="250" swimtime="00:03:41.89" />
                    <SPLIT distance="300" swimtime="00:04:27.31" />
                    <SPLIT distance="350" swimtime="00:05:12.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="WILCZĘGA" birthdate="1981-01-01" gender="M" nation="POL" swrid="4992879" athleteid="4027">
              <RESULTS>
                <RESULT eventid="1076" points="541" reactiontime="+69" swimtime="00:00:28.54" resultid="4501" heatid="4284" lane="0" entrytime="00:00:27.18" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="MATEUSZ" lastname="KĘDZIOR" birthdate="1973-01-01" gender="M" nation="POL" athleteid="3769">
              <RESULTS>
                <RESULT comment="Z3G8" eventid="1112" reactiontime="+97" status="DSQ" swimtime="00:00:00.00" resultid="3782" heatid="4294" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                    <SPLIT distance="100" swimtime="00:01:36.42" />
                    <SPLIT distance="150" swimtime="00:02:47.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="315" reactiontime="+111" swimtime="00:12:45.12" resultid="3783" heatid="4305" lane="6" entrytime="00:12:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="100" swimtime="00:01:24.30" />
                    <SPLIT distance="150" swimtime="00:02:11.51" />
                    <SPLIT distance="200" swimtime="00:03:00.00" />
                    <SPLIT distance="250" swimtime="00:03:49.37" />
                    <SPLIT distance="300" swimtime="00:04:40.22" />
                    <SPLIT distance="350" swimtime="00:05:28.59" />
                    <SPLIT distance="400" swimtime="00:06:18.23" />
                    <SPLIT distance="450" swimtime="00:07:05.58" />
                    <SPLIT distance="500" swimtime="00:07:54.14" />
                    <SPLIT distance="550" swimtime="00:08:43.68" />
                    <SPLIT distance="600" swimtime="00:09:32.14" />
                    <SPLIT distance="650" swimtime="00:10:21.56" />
                    <SPLIT distance="700" swimtime="00:11:10.95" />
                    <SPLIT distance="750" swimtime="00:11:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="332" reactiontime="+71" swimtime="00:00:39.89" resultid="3784" heatid="4321" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1301" points="329" reactiontime="+92" swimtime="00:01:15.65" resultid="3785" heatid="4346" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="250" reactiontime="+95" swimtime="00:01:35.46" resultid="3786" heatid="4391" lane="3" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="301" reactiontime="+93" swimtime="00:02:55.66" resultid="3787" heatid="4403" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:21.49" />
                    <SPLIT distance="150" swimtime="00:02:08.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="222" reactiontime="+103" swimtime="00:03:37.17" resultid="3788" heatid="4434" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.84" />
                    <SPLIT distance="100" swimtime="00:01:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="312" reactiontime="+103" swimtime="00:06:10.13" resultid="3789" heatid="4460" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:02:07.75" />
                    <SPLIT distance="200" swimtime="00:02:55.96" />
                    <SPLIT distance="250" swimtime="00:03:44.14" />
                    <SPLIT distance="300" swimtime="00:04:32.71" />
                    <SPLIT distance="350" swimtime="00:05:21.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="ALEKSANDRA" lastname="SAC" birthdate="1999-01-01" gender="F" nation="POL" athleteid="3932">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:03:09.60" resultid="3933" heatid="4289" lane="5" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="100" swimtime="00:01:30.22" />
                    <SPLIT distance="150" swimtime="00:02:25.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" swimtime="00:22:43.35" resultid="3934" heatid="4308" lane="5" entrytime="00:22:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:22.49" />
                    <SPLIT distance="150" swimtime="00:02:06.55" />
                    <SPLIT distance="200" swimtime="00:02:50.88" />
                    <SPLIT distance="250" swimtime="00:03:35.81" />
                    <SPLIT distance="300" swimtime="00:04:20.97" />
                    <SPLIT distance="350" swimtime="00:05:06.07" />
                    <SPLIT distance="400" swimtime="00:05:52.05" />
                    <SPLIT distance="450" swimtime="00:06:37.26" />
                    <SPLIT distance="500" swimtime="00:07:23.31" />
                    <SPLIT distance="550" swimtime="00:08:09.16" />
                    <SPLIT distance="600" swimtime="00:08:55.61" />
                    <SPLIT distance="650" swimtime="00:09:41.47" />
                    <SPLIT distance="700" swimtime="00:10:27.58" />
                    <SPLIT distance="750" swimtime="00:11:13.96" />
                    <SPLIT distance="800" swimtime="00:12:00.11" />
                    <SPLIT distance="850" swimtime="00:12:45.65" />
                    <SPLIT distance="900" swimtime="00:13:30.85" />
                    <SPLIT distance="950" swimtime="00:14:16.46" />
                    <SPLIT distance="1000" swimtime="00:15:02.53" />
                    <SPLIT distance="1050" swimtime="00:15:49.17" />
                    <SPLIT distance="1100" swimtime="00:16:35.64" />
                    <SPLIT distance="1150" swimtime="00:17:22.40" />
                    <SPLIT distance="1200" swimtime="00:18:09.57" />
                    <SPLIT distance="1250" swimtime="00:18:56.70" />
                    <SPLIT distance="1300" swimtime="00:19:43.90" />
                    <SPLIT distance="1350" swimtime="00:20:30.04" />
                    <SPLIT distance="1400" swimtime="00:21:16.17" />
                    <SPLIT distance="1450" swimtime="00:22:00.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1576" reactiontime="+73" swimtime="00:06:39.20" resultid="3935" heatid="4412" lane="6" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                    <SPLIT distance="100" swimtime="00:01:32.42" />
                    <SPLIT distance="150" swimtime="00:02:24.72" />
                    <SPLIT distance="200" swimtime="00:03:16.39" />
                    <SPLIT distance="250" swimtime="00:04:13.59" />
                    <SPLIT distance="300" swimtime="00:05:11.85" />
                    <SPLIT distance="350" swimtime="00:05:57.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" reactiontime="+77" swimtime="00:05:54.59" resultid="3936" heatid="4452" lane="8" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:24.29" />
                    <SPLIT distance="150" swimtime="00:02:09.44" />
                    <SPLIT distance="200" swimtime="00:02:55.49" />
                    <SPLIT distance="250" swimtime="00:03:41.69" />
                    <SPLIT distance="300" swimtime="00:04:27.30" />
                    <SPLIT distance="350" swimtime="00:05:12.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="DARIUSZ" lastname="SEWERYŃSKI" birthdate="1961-01-01" gender="M" nation="POL" athleteid="3977">
              <RESULTS>
                <RESULT eventid="1076" points="439" reactiontime="+103" swimtime="00:00:33.20" resultid="3978" heatid="4278" lane="2" entrytime="00:00:33.40" />
                <RESULT eventid="1301" points="374" reactiontime="+108" swimtime="00:01:20.24" resultid="3979" heatid="4344" lane="5" entrytime="00:01:32.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="299" reactiontime="+104" swimtime="00:03:32.29" resultid="3980" heatid="4293" lane="6" entrytime="00:03:30.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:01:43.46" />
                    <SPLIT distance="150" swimtime="00:02:45.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="325" reactiontime="+83" swimtime="00:03:52.99" resultid="3981" heatid="4332" lane="8" entrytime="00:03:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                    <SPLIT distance="100" swimtime="00:01:45.46" />
                    <SPLIT distance="150" swimtime="00:02:48.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="375" reactiontime="+97" swimtime="00:01:39.49" resultid="3982" heatid="4368" lane="3" entrytime="00:01:35.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="380" reactiontime="+103" swimtime="00:00:38.18" resultid="3983" heatid="4380" lane="8" entrytime="00:00:36.49" />
                <RESULT eventid="1629" points="250" reactiontime="+116" swimtime="00:01:38.47" resultid="3984" heatid="4424" lane="8" entrytime="00:01:32.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="446" reactiontime="+104" swimtime="00:00:42.92" resultid="3985" heatid="4445" lane="8" entrytime="00:00:41.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="ALICJA" lastname="GRUCA" birthdate="2000-01-01" gender="F" nation="POL" swrid="4647670" athleteid="3923">
              <RESULTS>
                <RESULT eventid="1094" reactiontime="+66" swimtime="00:02:52.75" resultid="3924" heatid="4290" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:20.21" />
                    <SPLIT distance="150" swimtime="00:02:09.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" reactiontime="+72" swimtime="00:03:09.06" resultid="3925" heatid="4328" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:01:29.70" />
                    <SPLIT distance="150" swimtime="00:02:19.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" reactiontime="+74" swimtime="00:01:27.01" resultid="3926" heatid="4365" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" reactiontime="+76" swimtime="00:00:33.97" resultid="3927" heatid="4374" lane="9" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="KATARZYNA" lastname="TYBURCZYK" birthdate="1977-01-01" gender="F" nation="POL" athleteid="3758">
              <RESULTS>
                <RESULT eventid="1059" points="43" swimtime="00:01:15.71" resultid="3762" heatid="4269" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1215" points="285" reactiontime="+76" swimtime="00:00:47.11" resultid="3763" heatid="4314" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="MAREK" lastname="MŁYNARCZYK" birthdate="1957-01-01" gender="M" nation="POL" athleteid="3757">
              <RESULTS>
                <RESULT eventid="1076" points="416" reactiontime="+78" swimtime="00:00:35.10" resultid="3759" heatid="4277" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1267" points="520" reactiontime="+71" swimtime="00:00:38.48" resultid="3760" heatid="4321" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3761" heatid="4391" lane="1" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="MICHAŁ" lastname="KOTULSKI" birthdate="1981-01-01" gender="M" nation="POL" athleteid="3824">
              <RESULTS>
                <RESULT eventid="1076" points="348" reactiontime="+82" swimtime="00:00:33.04" resultid="3825" heatid="4278" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1301" points="314" reactiontime="+78" swimtime="00:01:15.34" resultid="3826" heatid="4345" lane="6" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="412" reactiontime="+77" swimtime="00:00:33.68" resultid="3827" heatid="4380" lane="6" entrytime="00:00:34.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="MACIEJ" lastname="RYBICKI" birthdate="1963-01-01" gender="M" nation="POL" athleteid="3951">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3952" heatid="4279" lane="5" entrytime="00:00:31.20" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="3953" heatid="4380" lane="0" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="TOMASZ" lastname="BOCHEŃ" birthdate="1999-01-01" gender="M" nation="POL" athleteid="3730">
              <RESULTS>
                <RESULT eventid="1267" reactiontime="+66" swimtime="00:00:29.60" resultid="3731" heatid="4325" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1301" reactiontime="+65" swimtime="00:00:57.76" resultid="3732" heatid="4351" lane="6" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" reactiontime="+63" swimtime="00:00:26.43" resultid="3733" heatid="4384" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="1406" reactiontime="+62" swimtime="00:01:18.93" resultid="3734" heatid="4370" lane="0" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" reactiontime="+62" swimtime="00:00:59.57" resultid="3735" heatid="4427" lane="6" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" reactiontime="+63" swimtime="00:00:31.57" resultid="3736" heatid="4449" lane="0" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="KINGA" lastname="PARADOWSKA" birthdate="2001-01-01" gender="F" nation="POL" athleteid="3823" />
            <ATHLETE firstname="ŁUKASZ" lastname="BOGUSIAK" birthdate="1982-01-01" gender="M" nation="POL" athleteid="3928">
              <RESULTS>
                <RESULT eventid="1076" points="293" reactiontime="+85" swimtime="00:00:35.01" resultid="3929" heatid="4277" lane="4" entrytime="00:00:34.60" />
                <RESULT eventid="1301" points="281" reactiontime="+83" swimtime="00:01:18.18" resultid="3930" heatid="4345" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="3931" heatid="4402" lane="8" entrytime="00:02:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="ALEKSANDRA" lastname="HEBEL" birthdate="1987-01-01" gender="F" nation="POL" athleteid="3847">
              <RESULTS>
                <RESULT eventid="1059" points="436" reactiontime="+102" swimtime="00:00:34.26" resultid="3848" heatid="4270" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1284" points="415" reactiontime="+100" swimtime="00:01:17.85" resultid="3849" heatid="4339" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="380" reactiontime="+106" swimtime="00:02:53.89" resultid="3850" heatid="4398" lane="9" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="150" swimtime="00:02:08.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="325" reactiontime="+106" swimtime="00:03:20.98" resultid="3851" heatid="4431" lane="9" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                    <SPLIT distance="100" swimtime="00:01:38.18" />
                    <SPLIT distance="150" swimtime="00:02:30.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="EWELINA" lastname="CUCH" birthdate="1979-01-01" gender="F" nation="POL" athleteid="3815">
              <RESULTS>
                <RESULT eventid="1146" status="DNS" swimtime="00:00:00.00" resultid="3816" heatid="4300" lane="9" entrytime="00:13:45.00" />
                <RESULT eventid="1233" points="386" reactiontime="+95" swimtime="00:03:37.66" resultid="3817" heatid="4327" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                    <SPLIT distance="100" swimtime="00:01:39.37" />
                    <SPLIT distance="150" swimtime="00:02:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="389" reactiontime="+89" swimtime="00:01:19.53" resultid="3818" heatid="4335" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="426" reactiontime="+84" swimtime="00:01:36.64" resultid="3819" heatid="4364" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="459" reactiontime="+85" swimtime="00:00:36.76" resultid="3820" heatid="4374" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1680" points="392" reactiontime="+79" swimtime="00:00:44.37" resultid="3821" heatid="4440" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1731" points="338" reactiontime="+91" swimtime="00:06:17.51" resultid="3822" heatid="4453" lane="1" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:01:29.42" />
                    <SPLIT distance="150" swimtime="00:02:17.09" />
                    <SPLIT distance="200" swimtime="00:03:04.88" />
                    <SPLIT distance="250" swimtime="00:03:52.25" />
                    <SPLIT distance="300" swimtime="00:04:40.45" />
                    <SPLIT distance="350" swimtime="00:05:30.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="ROBERT" lastname="KAMIŃSKI " birthdate="1965-01-01" gender="M" nation="POL" athleteid="3804">
              <RESULTS>
                <RESULT eventid="1076" points="362" reactiontime="+86" swimtime="00:00:34.32" resultid="3805" heatid="4276" lane="5" entrytime="00:00:39.45" />
                <RESULT eventid="1267" points="397" reactiontime="+81" swimtime="00:00:39.51" resultid="3806" heatid="4321" lane="7" entrytime="00:00:44.45" />
                <RESULT eventid="1301" points="395" reactiontime="+91" swimtime="00:01:16.34" resultid="3807" heatid="4346" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="372" reactiontime="+85" swimtime="00:01:28.27" resultid="3808" heatid="4391" lane="7" entrytime="00:01:38.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="357" swimtime="00:03:18.58" resultid="3809" heatid="4434" lane="3" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                    <SPLIT distance="100" swimtime="00:03:18.58" />
                    <SPLIT distance="150" swimtime="00:02:24.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="ANDRZEJ" lastname="ŁOPUSZYŃSKI" birthdate="1969-01-01" gender="M" nation="POL" athleteid="3972">
              <RESULTS>
                <RESULT eventid="1112" points="155" reactiontime="+113" swimtime="00:04:04.10" resultid="3973" heatid="4292" lane="5" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.18" />
                    <SPLIT distance="100" swimtime="00:04:04.10" />
                    <SPLIT distance="150" swimtime="00:03:07.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="162" reactiontime="+113" swimtime="00:08:44.34" resultid="3974" heatid="4416" lane="9" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.35" />
                    <SPLIT distance="100" swimtime="00:01:54.50" />
                    <SPLIT distance="150" swimtime="00:03:08.61" />
                    <SPLIT distance="200" swimtime="00:04:27.17" />
                    <SPLIT distance="250" swimtime="00:05:35.22" />
                    <SPLIT distance="300" swimtime="00:06:45.93" />
                    <SPLIT distance="350" swimtime="00:07:45.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="161" reactiontime="+96" swimtime="00:04:05.27" resultid="3975" heatid="4355" lane="3" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.62" />
                    <SPLIT distance="100" swimtime="00:01:52.45" />
                    <SPLIT distance="150" swimtime="00:02:58.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="138" reactiontime="+101" swimtime="00:01:50.66" resultid="3976" heatid="4423" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="PAULINA" lastname="ZYGA" birthdate="1994-01-01" gender="F" nation="POL" athleteid="3750" />
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2725" name="iSwim Białystok">
          <CONTACT city="Białystok" email="biuro@iswim.bialystok.pl" name="Humbla Sebastian" phone="535309915" state="PDL" street="Wierzbowa 3C" zip="15-743" />
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Humbla" birthdate="1979-01-24" gender="M" nation="POL" swrid="4046250" athleteid="2726">
              <RESULTS>
                <RESULT eventid="1076" points="645" reactiontime="+72" swimtime="00:00:26.91" resultid="2727" heatid="4283" lane="2" entrytime="00:00:27.65" entrycourse="LCM" />
                <RESULT eventid="1267" points="570" reactiontime="+70" swimtime="00:00:32.73" resultid="2728" heatid="4324" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1457" points="620" reactiontime="+67" swimtime="00:00:29.39" resultid="2729" heatid="4383" lane="7" entrytime="00:00:28.90" />
                <RESULT eventid="1697" status="DNS" swimtime="00:00:00.00" resultid="2730" heatid="4447" lane="2" entrytime="00:00:35.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elżbieta" lastname="Piwowarczyk" birthdate="1966-01-06" gender="F" nation="POL" swrid="4186247" athleteid="2736">
              <RESULTS>
                <RESULT eventid="1059" points="534" reactiontime="+63" swimtime="00:00:34.86" resultid="2737" heatid="4269" lane="5" entrytime="00:00:36.50" />
                <RESULT eventid="1215" points="381" reactiontime="+78" swimtime="00:00:44.14" resultid="2738" heatid="4314" lane="5" entrytime="00:00:45.50" />
                <RESULT eventid="1284" points="510" reactiontime="+75" swimtime="00:01:17.61" resultid="2739" heatid="4338" lane="1" entrytime="00:01:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="420" reactiontime="+91" swimtime="00:01:33.05" resultid="2740" heatid="4387" lane="3" entrytime="00:01:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="474" reactiontime="+78" swimtime="00:02:54.75" resultid="2741" heatid="4397" lane="3" entrytime="00:02:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                    <SPLIT distance="150" swimtime="00:02:10.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" status="DNS" swimtime="00:00:00.00" resultid="2742" heatid="4430" lane="3" entrytime="00:03:25.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Świderski" birthdate="1979-02-13" gender="M" nation="POL" swrid="5422007" athleteid="2731">
              <RESULTS>
                <RESULT eventid="1076" points="673" reactiontime="+74" swimtime="00:00:26.53" resultid="2732" heatid="4285" lane="1" entrytime="00:00:26.49" />
                <RESULT eventid="1301" points="616" reactiontime="+81" swimtime="00:01:00.20" resultid="2733" heatid="4349" lane="4" entrytime="00:01:00.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="693" reactiontime="+75" swimtime="00:00:28.32" resultid="2734" heatid="4383" lane="3" entrytime="00:00:28.16" entrycourse="LCM" />
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="2735" heatid="4426" lane="6" entrytime="00:01:04.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3722" name="Szczytno">
          <ATHLETES>
            <ATHLETE firstname="ZDZISŁAW" lastname="CHOROSZEWSKI" birthdate="1947-01-01" gender="M" nation="POL" athleteid="3723">
              <RESULTS>
                <RESULT eventid="1076" points="242" reactiontime="+95" swimtime="00:00:46.86" resultid="3724" heatid="4276" lane="0" entrytime="00:00:46.00" />
                <RESULT eventid="1197" points="221" swimtime="00:34:48.99" resultid="3725" heatid="4311" lane="7" entrytime="00:40:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.89" />
                    <SPLIT distance="100" swimtime="00:02:07.93" />
                    <SPLIT distance="150" swimtime="00:03:19.66" />
                    <SPLIT distance="200" swimtime="00:04:31.44" />
                    <SPLIT distance="250" swimtime="00:05:42.63" />
                    <SPLIT distance="300" swimtime="00:06:51.73" />
                    <SPLIT distance="350" swimtime="00:08:01.82" />
                    <SPLIT distance="400" swimtime="00:09:12.55" />
                    <SPLIT distance="450" swimtime="00:10:23.37" />
                    <SPLIT distance="500" swimtime="00:11:32.16" />
                    <SPLIT distance="550" swimtime="00:12:40.83" />
                    <SPLIT distance="600" swimtime="00:13:51.43" />
                    <SPLIT distance="650" swimtime="00:15:00.81" />
                    <SPLIT distance="700" swimtime="00:16:10.51" />
                    <SPLIT distance="750" swimtime="00:17:21.27" />
                    <SPLIT distance="800" swimtime="00:18:31.24" />
                    <SPLIT distance="850" swimtime="00:19:42.65" />
                    <SPLIT distance="900" swimtime="00:20:50.87" />
                    <SPLIT distance="950" swimtime="00:22:02.11" />
                    <SPLIT distance="1000" swimtime="00:23:13.68" />
                    <SPLIT distance="1050" swimtime="00:24:25.11" />
                    <SPLIT distance="1100" swimtime="00:25:34.46" />
                    <SPLIT distance="1150" swimtime="00:26:46.74" />
                    <SPLIT distance="1200" swimtime="00:27:55.77" />
                    <SPLIT distance="1250" swimtime="00:29:06.92" />
                    <SPLIT distance="1300" swimtime="00:30:17.71" />
                    <SPLIT distance="1350" swimtime="00:31:28.99" />
                    <SPLIT distance="1400" swimtime="00:32:36.83" />
                    <SPLIT distance="1450" swimtime="00:33:47.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="201" reactiontime="+85" swimtime="00:01:53.33" resultid="3726" heatid="4344" lane="0" entrytime="00:01:52.00" />
                <RESULT eventid="1525" points="167" reactiontime="+104" swimtime="00:04:24.40" resultid="3727" heatid="4401" lane="6" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.44" />
                    <SPLIT distance="100" swimtime="00:02:12.27" />
                    <SPLIT distance="150" swimtime="00:03:23.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="202" reactiontime="+89" swimtime="00:09:01.57" resultid="3728" heatid="4461" lane="9" entrytime="00:09:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.21" />
                    <SPLIT distance="100" swimtime="00:02:08.00" />
                    <SPLIT distance="150" swimtime="00:03:20.53" />
                    <SPLIT distance="200" swimtime="00:04:31.72" />
                    <SPLIT distance="250" swimtime="00:05:42.81" />
                    <SPLIT distance="300" swimtime="00:06:52.28" />
                    <SPLIT distance="350" swimtime="00:08:01.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00305" nation="POL" region="05" clubid="2615" name="UKS Nawa Skierniewice">
          <ATHLETES>
            <ATHLETE firstname="Pamela" lastname="Broniarek" birthdate="1995-11-21" gender="F" nation="POL" license="100305600178" athleteid="2637">
              <RESULTS>
                <RESULT eventid="1146" points="500" reactiontime="+127" swimtime="00:11:02.66" resultid="2638" heatid="4301" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:02:00.46" />
                    <SPLIT distance="200" swimtime="00:02:42.48" />
                    <SPLIT distance="250" swimtime="00:03:25.45" />
                    <SPLIT distance="300" swimtime="00:04:06.57" />
                    <SPLIT distance="350" swimtime="00:04:49.42" />
                    <SPLIT distance="400" swimtime="00:05:31.68" />
                    <SPLIT distance="450" swimtime="00:06:13.55" />
                    <SPLIT distance="500" swimtime="00:06:55.33" />
                    <SPLIT distance="550" swimtime="00:07:37.63" />
                    <SPLIT distance="600" swimtime="00:08:19.24" />
                    <SPLIT distance="650" swimtime="00:09:01.19" />
                    <SPLIT distance="700" swimtime="00:09:41.76" />
                    <SPLIT distance="750" swimtime="00:10:23.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Białkowska" birthdate="1997-02-13" gender="F" nation="POL" license="100305600117" swrid="4287915" athleteid="2616">
              <RESULTS>
                <RESULT eventid="1059" status="WDR" swimtime="00:00:00.00" resultid="2617" />
                <RESULT eventid="1215" points="426" reactiontime="+81" swimtime="00:00:37.74" resultid="2618" heatid="4312" lane="7" />
                <RESULT eventid="1284" points="508" reactiontime="+85" swimtime="00:01:11.39" resultid="2619" heatid="4336" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="427" reactiontime="+85" swimtime="00:01:21.80" resultid="2620" heatid="4385" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Sarna" birthdate="1998-12-02" gender="F" nation="POL" license="100305600120" swrid="4476652" athleteid="2631">
              <RESULTS>
                <RESULT eventid="1094" status="WDR" swimtime="00:00:00.00" resultid="2632" />
                <RESULT eventid="1215" reactiontime="+71" swimtime="00:00:34.49" resultid="2633" heatid="4312" lane="1" />
                <RESULT eventid="1440" reactiontime="+80" swimtime="00:00:33.45" resultid="2635" heatid="4373" lane="0" />
                <RESULT eventid="1611" reactiontime="+86" swimtime="00:01:18.32" resultid="2636" heatid="4419" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Dębski" birthdate="1998-08-01" gender="M" nation="POL" license="100305700340" swrid="4476651" athleteid="2621">
              <RESULTS>
                <RESULT eventid="1076" reactiontime="+73" swimtime="00:00:26.88" resultid="2622" heatid="4273" lane="3" />
                <RESULT eventid="1301" status="WDR" swimtime="00:00:00.00" resultid="2623" />
                <RESULT eventid="1457" reactiontime="+73" swimtime="00:00:28.88" resultid="2624" heatid="4376" lane="3" />
                <RESULT eventid="1629" reactiontime="+72" swimtime="00:01:11.80" resultid="2625" heatid="4422" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Zyga" birthdate="1994-12-15" gender="F" nation="POL" license="100305600193" swrid="4806433" athleteid="2626">
              <RESULTS>
                <RESULT eventid="1094" status="WDR" swimtime="00:00:00.00" resultid="2627" entrytime="00:03:00.00" />
                <RESULT eventid="1284" points="503" reactiontime="+69" swimtime="00:01:11.61" resultid="2628" heatid="4339" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="449" reactiontime="+72" swimtime="00:02:42.69" resultid="2629" heatid="4398" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:01:59.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="407" reactiontime="+79" swimtime="00:02:59.70" resultid="2630" heatid="4431" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                    <SPLIT distance="100" swimtime="00:01:27.31" />
                    <SPLIT distance="150" swimtime="00:02:14.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1542" status="DNS" swimtime="00:00:00.00" resultid="2641" heatid="4494" lane="1" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="GER" clubid="2743" name="SG Erkelenz-Kuckelhoven">
          <CONTACT name="Gożdziejewska" />
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Andrzejczak" birthdate="1967-01-29" gender="M" nation="GER" athleteid="2744">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1076" points="761" reactiontime="+77" swimtime="00:00:26.78" resultid="2745" heatid="4284" lane="4" entrytime="00:00:26.68" />
                <RESULT eventid="1267" points="656" reactiontime="+65" swimtime="00:00:33.41" resultid="2746" heatid="4323" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1301" points="808" reactiontime="+80" swimtime="00:01:00.12" resultid="2747" heatid="4349" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="730" reactiontime="+81" swimtime="00:00:29.50" resultid="2748" heatid="4382" lane="6" entrytime="00:00:29.22" />
                <RESULT eventid="1525" points="696" reactiontime="+83" swimtime="00:02:19.94" resultid="2749" heatid="4406" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:06.50" />
                    <SPLIT distance="150" swimtime="00:01:43.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="638" reactiontime="+84" swimtime="00:00:34.88" resultid="2750" heatid="4448" lane="9" entrytime="00:00:34.72" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3649" name="MKS Juvenia Białystok">
          <CONTACT email="wzmasters@wp.pl" name="Żmiejko" phone="797309140" />
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Żmiejko" birthdate="1963-01-01" gender="M" nation="POL" license="500309700377" swrid="4186249" athleteid="3655">
              <RESULTS>
                <RESULT eventid="1076" points="576" reactiontime="+76" swimtime="00:00:29.38" resultid="3656" heatid="4281" lane="8" entrytime="00:00:29.35" />
                <RESULT eventid="1112" points="595" reactiontime="+78" swimtime="00:02:47.22" resultid="3657" heatid="4295" lane="1" entrytime="00:02:47.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:18.11" />
                    <SPLIT distance="150" swimtime="00:02:07.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="641" reactiontime="+77" swimtime="00:01:04.96" resultid="3658" heatid="4348" lane="0" entrytime="00:01:05.83" entrycourse="LCM" />
                <RESULT eventid="1457" points="620" reactiontime="+78" swimtime="00:00:31.15" resultid="3659" heatid="4381" lane="2" entrytime="00:00:31.10" entrycourse="LCM" />
                <RESULT eventid="1491" points="504" reactiontime="+84" swimtime="00:01:19.81" resultid="3660" heatid="4392" lane="6" entrytime="00:01:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="533" reactiontime="+79" swimtime="00:01:14.71" resultid="3661" heatid="4425" lane="8" entrytime="00:01:12.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="491" reactiontime="+78" swimtime="00:00:38.06" resultid="3662" heatid="4446" lane="7" entrytime="00:00:37.75" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Michalik" birthdate="1979-01-01" gender="F" nation="POL" license="500309600228" swrid="4595750" athleteid="3650">
              <RESULTS>
                <RESULT eventid="1146" points="570" reactiontime="+79" swimtime="00:10:50.07" resultid="3651" heatid="4300" lane="3" entrytime="00:10:24.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                    <SPLIT distance="150" swimtime="00:01:56.68" />
                    <SPLIT distance="200" swimtime="00:02:38.16" />
                    <SPLIT distance="250" swimtime="00:03:19.47" />
                    <SPLIT distance="300" swimtime="00:04:00.47" />
                    <SPLIT distance="350" swimtime="00:04:42.00" />
                    <SPLIT distance="400" swimtime="00:05:23.49" />
                    <SPLIT distance="450" swimtime="00:06:04.40" />
                    <SPLIT distance="500" swimtime="00:06:45.40" />
                    <SPLIT distance="550" swimtime="00:07:26.30" />
                    <SPLIT distance="600" swimtime="00:08:06.90" />
                    <SPLIT distance="650" swimtime="00:08:47.32" />
                    <SPLIT distance="700" swimtime="00:09:29.39" />
                    <SPLIT distance="750" swimtime="00:10:10.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="693" reactiontime="+66" swimtime="00:01:05.58" resultid="3652" heatid="4340" lane="7" entrytime="00:01:04.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="718" reactiontime="+75" swimtime="00:02:24.36" resultid="3653" heatid="4398" lane="5" entrytime="00:02:22.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:48.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="599" reactiontime="+77" swimtime="00:05:11.89" resultid="3654" heatid="4452" lane="3" entrytime="00:05:01.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:52.41" />
                    <SPLIT distance="200" swimtime="00:02:32.28" />
                    <SPLIT distance="250" swimtime="00:03:12.13" />
                    <SPLIT distance="300" swimtime="00:03:52.83" />
                    <SPLIT distance="350" swimtime="00:04:33.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TMT" nation="POL" clubid="3522" name="Toruń Multisport Team">
          <CONTACT city="Toruń" email="g.arentewicz@onet.pl" name="Arentewicz" phone="535-763-476" state="KUJ-P" zip="87-100" />
          <ATHLETES>
            <ATHLETE firstname="Anita" lastname="Śliwa" birthdate="1972-09-24" gender="F" nation="POL" athleteid="3531">
              <RESULTS>
                <RESULT eventid="1094" points="247" reactiontime="+96" swimtime="00:04:00.69" resultid="3532" heatid="4288" lane="5" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.86" />
                    <SPLIT distance="100" swimtime="00:01:51.87" />
                    <SPLIT distance="150" swimtime="00:03:05.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="236" reactiontime="+102" swimtime="00:15:28.48" resultid="3533" heatid="4302" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.83" />
                    <SPLIT distance="100" swimtime="00:01:40.55" />
                    <SPLIT distance="150" swimtime="00:02:38.48" />
                    <SPLIT distance="200" swimtime="00:03:37.71" />
                    <SPLIT distance="250" swimtime="00:04:36.68" />
                    <SPLIT distance="300" swimtime="00:05:36.58" />
                    <SPLIT distance="350" swimtime="00:06:35.68" />
                    <SPLIT distance="400" swimtime="00:07:35.04" />
                    <SPLIT distance="450" swimtime="00:08:34.27" />
                    <SPLIT distance="500" swimtime="00:09:33.95" />
                    <SPLIT distance="550" swimtime="00:10:33.58" />
                    <SPLIT distance="600" swimtime="00:11:33.54" />
                    <SPLIT distance="650" swimtime="00:12:34.10" />
                    <SPLIT distance="700" swimtime="00:13:33.63" />
                    <SPLIT distance="750" swimtime="00:14:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="276" reactiontime="+101" swimtime="00:00:48.49" resultid="3534" heatid="4314" lane="3" entrytime="00:00:47.00" />
                <RESULT eventid="1284" points="269" reactiontime="+99" swimtime="00:01:33.54" resultid="3535" heatid="4337" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="260" reactiontime="+92" swimtime="00:01:46.78" resultid="3536" heatid="4387" lane="2" entrytime="00:01:44.00" />
                <RESULT eventid="1646" points="265" reactiontime="+92" swimtime="00:03:48.23" resultid="3537" heatid="4430" lane="2" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                    <SPLIT distance="100" swimtime="00:01:50.80" />
                    <SPLIT distance="150" swimtime="00:02:51.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="249" reactiontime="+103" swimtime="00:07:26.32" resultid="3538" heatid="4454" lane="5" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:41.53" />
                    <SPLIT distance="150" swimtime="00:02:39.00" />
                    <SPLIT distance="200" swimtime="00:03:37.28" />
                    <SPLIT distance="250" swimtime="00:04:35.96" />
                    <SPLIT distance="300" swimtime="00:05:34.38" />
                    <SPLIT distance="350" swimtime="00:06:32.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Gołembiewski" birthdate="1986-10-28" gender="M" nation="POL" athleteid="3523">
              <RESULTS>
                <RESULT eventid="1112" points="493" reactiontime="+82" swimtime="00:02:39.07" resultid="3524" heatid="4296" lane="1" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:02.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="476" reactiontime="+87" swimtime="00:10:38.23" resultid="3525" heatid="4303" lane="1" entrytime="00:10:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                    <SPLIT distance="100" swimtime="00:01:11.15" />
                    <SPLIT distance="150" swimtime="00:01:49.69" />
                    <SPLIT distance="200" swimtime="00:02:29.51" />
                    <SPLIT distance="250" swimtime="00:03:09.79" />
                    <SPLIT distance="300" swimtime="00:03:50.83" />
                    <SPLIT distance="350" swimtime="00:04:31.92" />
                    <SPLIT distance="400" swimtime="00:05:13.49" />
                    <SPLIT distance="450" swimtime="00:05:54.81" />
                    <SPLIT distance="500" swimtime="00:06:36.27" />
                    <SPLIT distance="550" swimtime="00:07:17.71" />
                    <SPLIT distance="600" swimtime="00:07:59.17" />
                    <SPLIT distance="650" swimtime="00:08:39.77" />
                    <SPLIT distance="700" swimtime="00:09:20.15" />
                    <SPLIT distance="750" swimtime="00:09:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="592" reactiontime="+76" swimtime="00:02:47.05" resultid="3526" heatid="4334" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:03.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="653" reactiontime="+79" swimtime="00:01:11.91" resultid="3527" heatid="4371" lane="1" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="3528" heatid="4406" lane="6" entrytime="00:02:11.00" />
                <RESULT eventid="1697" points="617" reactiontime="+83" swimtime="00:00:33.44" resultid="3529" heatid="4449" lane="8" entrytime="00:00:32.40" />
                <RESULT eventid="1748" points="527" reactiontime="+77" swimtime="00:05:04.44" resultid="3530" heatid="4457" lane="5" entrytime="00:04:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                    <SPLIT distance="150" swimtime="00:01:47.33" />
                    <SPLIT distance="200" swimtime="00:02:25.58" />
                    <SPLIT distance="250" swimtime="00:03:04.56" />
                    <SPLIT distance="300" swimtime="00:03:44.62" />
                    <SPLIT distance="350" swimtime="00:04:25.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Kordowski" birthdate="1997-10-11" gender="M" nation="POL" athleteid="3562">
              <RESULTS>
                <RESULT eventid="1076" points="568" reactiontime="+69" swimtime="00:00:26.92" resultid="3563" heatid="4284" lane="5" entrytime="00:00:26.70" />
                <RESULT eventid="1301" points="582" reactiontime="+76" swimtime="00:01:00.43" resultid="3564" heatid="4350" lane="8" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="548" reactiontime="+74" swimtime="00:00:28.98" resultid="3565" heatid="4382" lane="3" entrytime="00:00:29.20" />
                <RESULT eventid="1629" points="407" reactiontime="+73" swimtime="00:01:11.63" resultid="3566" heatid="4425" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Bilski" birthdate="1984-08-01" gender="M" nation="POL" athleteid="3581">
              <RESULTS>
                <RESULT eventid="1163" points="196" reactiontime="+143" swimtime="00:14:17.40" resultid="3582" heatid="4306" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                    <SPLIT distance="100" swimtime="00:01:39.11" />
                    <SPLIT distance="150" swimtime="00:02:32.58" />
                    <SPLIT distance="200" swimtime="00:03:26.55" />
                    <SPLIT distance="250" swimtime="00:04:21.07" />
                    <SPLIT distance="300" swimtime="00:05:15.36" />
                    <SPLIT distance="350" swimtime="00:06:11.27" />
                    <SPLIT distance="400" swimtime="00:07:06.53" />
                    <SPLIT distance="450" swimtime="00:08:01.21" />
                    <SPLIT distance="500" swimtime="00:08:55.45" />
                    <SPLIT distance="550" swimtime="00:09:49.82" />
                    <SPLIT distance="600" swimtime="00:10:43.86" />
                    <SPLIT distance="650" swimtime="00:11:39.17" />
                    <SPLIT distance="700" swimtime="00:12:33.36" />
                    <SPLIT distance="750" swimtime="00:13:27.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henryk" lastname="Zientara" birthdate="1946-03-03" gender="M" nation="POL" swrid="4754680" athleteid="3573">
              <RESULTS>
                <RESULT eventid="1076" points="211" reactiontime="+106" swimtime="00:00:49.01" resultid="3574" heatid="4276" lane="6" entrytime="00:00:42.12" />
                <RESULT eventid="1267" points="220" reactiontime="+89" swimtime="00:00:57.04" resultid="3575" heatid="4321" lane="9" entrytime="00:00:52.35" />
                <RESULT eventid="1250" points="230" reactiontime="+96" swimtime="00:05:16.46" resultid="3576" heatid="4331" lane="0" entrytime="00:04:31.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.09" />
                    <SPLIT distance="100" swimtime="00:02:30.89" />
                    <SPLIT distance="150" swimtime="00:03:57.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="248" reactiontime="+99" swimtime="00:02:19.71" resultid="3577" heatid="4367" lane="2" entrytime="00:02:06.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="154" reactiontime="+94" swimtime="00:02:24.02" resultid="3578" heatid="4390" lane="1" entrytime="00:02:21.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="135" reactiontime="+103" swimtime="00:05:31.73" resultid="3579" heatid="4433" lane="5" entrytime="00:04:51.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.21" />
                    <SPLIT distance="100" swimtime="00:02:44.30" />
                    <SPLIT distance="150" swimtime="00:04:10.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="266" reactiontime="+93" swimtime="00:01:00.74" resultid="3580" heatid="4444" lane="8" entrytime="00:00:49.08" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucyna" lastname="Serożyńska" birthdate="1955-06-29" gender="F" nation="POL" athleteid="3553">
              <RESULTS>
                <RESULT eventid="1059" points="178" reactiontime="+109" swimtime="00:00:51.76" resultid="3554" heatid="4268" lane="4" entrytime="00:00:54.27" />
                <RESULT eventid="1146" reactiontime="+143" status="DNS" swimtime="00:00:00.00" resultid="3555" heatid="4301" lane="2" entrytime="00:20:00.00" />
                <RESULT eventid="1215" points="153" reactiontime="+103" swimtime="00:01:02.85" resultid="3556" heatid="4313" lane="4" entrytime="00:01:03.00" />
                <RESULT eventid="1284" points="145" reactiontime="+120" swimtime="00:02:03.53" resultid="3557" heatid="4337" lane="1" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="277" reactiontime="+112" swimtime="00:02:18.52" resultid="3558" heatid="4363" lane="5" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="162" reactiontime="+97" swimtime="00:02:16.62" resultid="3559" heatid="4387" lane="0" entrytime="00:02:19.00" />
                <RESULT eventid="1646" points="201" reactiontime="+113" swimtime="00:04:46.24" resultid="3560" heatid="4430" lane="8" entrytime="00:04:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.98" />
                    <SPLIT distance="100" swimtime="00:02:21.27" />
                    <SPLIT distance="150" swimtime="00:03:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="223" reactiontime="+120" swimtime="00:08:36.12" resultid="3561" heatid="4454" lane="1" entrytime="00:08:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.95" />
                    <SPLIT distance="100" swimtime="00:02:09.46" />
                    <SPLIT distance="150" swimtime="00:03:19.04" />
                    <SPLIT distance="200" swimtime="00:04:29.02" />
                    <SPLIT distance="250" swimtime="00:05:39.21" />
                    <SPLIT distance="300" swimtime="00:06:52.18" />
                    <SPLIT distance="350" swimtime="00:08:02.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Lietz" birthdate="1952-04-23" gender="M" nation="POL" athleteid="3546">
              <RESULTS>
                <RESULT eventid="1076" points="507" reactiontime="+83" swimtime="00:00:34.76" resultid="3547" heatid="4278" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1163" points="385" reactiontime="+94" swimtime="00:14:36.85" resultid="3548" heatid="4305" lane="1" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                    <SPLIT distance="100" swimtime="00:01:39.61" />
                    <SPLIT distance="150" swimtime="00:02:35.57" />
                    <SPLIT distance="200" swimtime="00:03:31.89" />
                    <SPLIT distance="250" swimtime="00:04:27.99" />
                    <SPLIT distance="300" swimtime="00:05:23.85" />
                    <SPLIT distance="350" swimtime="00:06:19.82" />
                    <SPLIT distance="400" swimtime="00:07:17.23" />
                    <SPLIT distance="450" swimtime="00:08:13.59" />
                    <SPLIT distance="500" swimtime="00:09:10.68" />
                    <SPLIT distance="550" swimtime="00:10:07.02" />
                    <SPLIT distance="600" swimtime="00:11:03.80" />
                    <SPLIT distance="650" swimtime="00:11:59.64" />
                    <SPLIT distance="700" swimtime="00:12:55.34" />
                    <SPLIT distance="750" swimtime="00:13:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="470" reactiontime="+77" swimtime="00:01:21.45" resultid="3549" heatid="4346" lane="9" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="406" reactiontime="+78" swimtime="00:00:40.49" resultid="3550" heatid="4380" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1525" points="446" reactiontime="+84" swimtime="00:03:07.60" resultid="3551" heatid="4402" lane="1" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:01:31.95" />
                    <SPLIT distance="150" swimtime="00:02:22.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="402" reactiontime="+88" swimtime="00:06:51.29" resultid="3552" heatid="4460" lane="0" entrytime="00:06:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.68" />
                    <SPLIT distance="100" swimtime="00:01:35.59" />
                    <SPLIT distance="200" swimtime="00:03:22.32" />
                    <SPLIT distance="250" swimtime="00:04:17.03" />
                    <SPLIT distance="300" swimtime="00:05:10.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Lisiecki" birthdate="1982-01-28" gender="M" nation="POL" athleteid="3539">
              <RESULTS>
                <RESULT eventid="1112" points="388" reactiontime="+91" swimtime="00:02:59.16" resultid="3540" heatid="4291" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:22.20" />
                    <SPLIT distance="150" swimtime="00:02:15.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="358" reactiontime="+100" swimtime="00:12:06.44" resultid="3541" heatid="4307" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="100" swimtime="00:01:22.60" />
                    <SPLIT distance="150" swimtime="00:02:07.90" />
                    <SPLIT distance="200" swimtime="00:02:53.56" />
                    <SPLIT distance="250" swimtime="00:03:39.61" />
                    <SPLIT distance="300" swimtime="00:04:25.97" />
                    <SPLIT distance="350" swimtime="00:05:12.06" />
                    <SPLIT distance="400" swimtime="00:05:58.57" />
                    <SPLIT distance="450" swimtime="00:06:44.16" />
                    <SPLIT distance="500" swimtime="00:07:30.29" />
                    <SPLIT distance="550" swimtime="00:08:16.60" />
                    <SPLIT distance="600" swimtime="00:09:02.92" />
                    <SPLIT distance="650" swimtime="00:09:49.61" />
                    <SPLIT distance="700" swimtime="00:10:35.59" />
                    <SPLIT distance="750" swimtime="00:11:21.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="333" reactiontime="+93" swimtime="00:01:24.30" resultid="3542" heatid="4392" lane="1" entrytime="00:01:24.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="402" reactiontime="+98" swimtime="00:06:23.58" resultid="3543" heatid="4418" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                    <SPLIT distance="100" swimtime="00:01:29.78" />
                    <SPLIT distance="150" swimtime="00:02:17.07" />
                    <SPLIT distance="200" swimtime="00:03:05.31" />
                    <SPLIT distance="250" swimtime="00:04:00.17" />
                    <SPLIT distance="300" swimtime="00:04:55.65" />
                    <SPLIT distance="350" swimtime="00:05:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="365" reactiontime="+90" swimtime="00:02:59.16" resultid="3544" heatid="4435" lane="1" entrytime="00:03:02.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:26.36" />
                    <SPLIT distance="150" swimtime="00:02:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="360" reactiontime="+93" swimtime="00:05:46.70" resultid="3545" heatid="4459" lane="1" entrytime="00:05:38.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="150" swimtime="00:02:02.22" />
                    <SPLIT distance="200" swimtime="00:02:47.15" />
                    <SPLIT distance="250" swimtime="00:03:32.49" />
                    <SPLIT distance="300" swimtime="00:04:17.93" />
                    <SPLIT distance="350" swimtime="00:05:03.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Korolko" birthdate="1940-10-13" gender="M" nation="POL" athleteid="3567">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3568" heatid="4276" lane="7" entrytime="00:00:44.80" />
                <RESULT eventid="1267" status="DNS" swimtime="00:00:00.00" resultid="3569" heatid="4320" lane="0" entrytime="00:01:05.20" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="3570" heatid="4344" lane="1" entrytime="00:01:45.65" />
                <RESULT eventid="1491" points="114" swimtime="00:02:58.15" resultid="3571" heatid="4390" lane="2" entrytime="00:02:12.15" />
                <RESULT eventid="1663" status="DNS" swimtime="00:00:00.00" resultid="3572" heatid="4433" lane="6" entrytime="00:05:09.45" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" points="257" reactiontime="+81" swimtime="00:03:00.20" resultid="3583" heatid="4488" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.38" />
                    <SPLIT distance="100" swimtime="00:01:44.53" />
                    <SPLIT distance="150" swimtime="00:02:19.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3573" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3553" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="3546" number="3" reactiontime="-80" />
                    <RELAYPOSITION athleteid="3531" number="4" reactiontime="+82" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="11514" nation="POL" region="14" clubid="2488" name="Stowarzyszenie Pływackie Sebastiana Karasia">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Karczewski" birthdate="1974-07-07" gender="M" nation="POL" license="511514700195" athleteid="2497">
              <RESULTS>
                <RESULT eventid="1076" points="351" reactiontime="+83" swimtime="00:00:33.40" resultid="2498" heatid="4274" lane="2" />
                <RESULT eventid="1301" points="277" reactiontime="+82" swimtime="00:01:20.18" resultid="2499" heatid="4342" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="2500" heatid="4401" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Witek" birthdate="1984-09-22" gender="M" nation="POL" license="511514700194" athleteid="2514">
              <RESULTS>
                <RESULT eventid="1748" points="325" reactiontime="+74" swimtime="00:05:57.61" resultid="2515" heatid="4463" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:16.96" />
                    <SPLIT distance="150" swimtime="00:02:02.67" />
                    <SPLIT distance="200" swimtime="00:02:52.14" />
                    <SPLIT distance="250" swimtime="00:03:41.24" />
                    <SPLIT distance="300" swimtime="00:04:29.23" />
                    <SPLIT distance="350" swimtime="00:05:14.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Frąckowiak" birthdate="1980-12-04" gender="M" nation="POL" license="511514700192" athleteid="2501">
              <RESULTS>
                <RESULT eventid="1076" points="442" reactiontime="+78" swimtime="00:00:30.53" resultid="2502" heatid="4275" lane="1" />
                <RESULT eventid="1301" points="428" reactiontime="+77" swimtime="00:01:07.93" resultid="2503" heatid="4343" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="384" reactiontime="+80" swimtime="00:05:39.48" resultid="2504" heatid="4463" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:02:02.22" />
                    <SPLIT distance="200" swimtime="00:02:46.62" />
                    <SPLIT distance="250" swimtime="00:03:30.84" />
                    <SPLIT distance="300" swimtime="00:04:15.12" />
                    <SPLIT distance="350" swimtime="00:04:58.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Łukasiuk" birthdate="1980-01-02" gender="F" nation="POL" license="511514600187" athleteid="2489">
              <RESULTS>
                <RESULT eventid="1059" points="524" reactiontime="+67" swimtime="00:00:32.80" resultid="2490" heatid="4267" lane="8" />
                <RESULT eventid="1284" status="DNS" swimtime="00:00:00.00" resultid="2491" heatid="4336" lane="4" />
                <RESULT eventid="1404" points="478" reactiontime="+77" swimtime="00:01:33.04" resultid="2492" heatid="4362" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="517" reactiontime="+77" swimtime="00:00:40.45" resultid="2493" heatid="4439" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Bistron" birthdate="1989-06-30" gender="M" nation="POL" license="511514700191" athleteid="2507">
              <RESULTS>
                <RESULT eventid="1250" status="DNS" swimtime="00:00:00.00" resultid="2508" heatid="4329" lane="6" />
                <RESULT eventid="1352" points="172" reactiontime="+77" swimtime="00:03:41.74" resultid="2509" heatid="4355" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="100" swimtime="00:01:40.79" />
                    <SPLIT distance="150" swimtime="00:02:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="68" swimtime="00:02:16.73" resultid="2510" heatid="4389" lane="8" />
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="2511" heatid="4418" lane="6" />
                <RESULT eventid="1663" status="DNS" swimtime="00:00:00.00" resultid="2512" heatid="4432" lane="2" />
                <RESULT eventid="1697" status="DNS" swimtime="00:00:00.00" resultid="2513" heatid="4442" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Fuliński" birthdate="1982-06-03" gender="M" nation="POL" license="111514700186" swrid="4992686" athleteid="2494">
              <RESULTS>
                <RESULT eventid="1076" points="641" reactiontime="+77" swimtime="00:00:26.97" resultid="2495" heatid="4284" lane="3" entrytime="00:00:26.73" />
                <RESULT eventid="1301" points="651" reactiontime="+82" swimtime="00:00:59.10" resultid="2496" heatid="4350" lane="3" entrytime="00:00:59.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Diaby - Lipka" birthdate="1980-08-30" gender="F" nation="POL" license="111514600193" athleteid="2505">
              <RESULTS>
                <RESULT eventid="1215" points="571" reactiontime="+75" swimtime="00:00:35.71" resultid="2506" heatid="4312" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1559" points="548" reactiontime="+81" swimtime="00:01:55.97" resultid="2516" heatid="4496" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                    <SPLIT distance="100" swimtime="00:00:58.73" />
                    <SPLIT distance="150" swimtime="00:01:28.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2494" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2497" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="2501" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="2514" number="4" reactiontime="+5" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1714" points="545" reactiontime="+94" swimtime="00:02:18.64" resultid="2517" heatid="4499" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:15.68" />
                    <SPLIT distance="150" swimtime="00:01:45.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2505" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="2494" number="2" />
                    <RELAYPOSITION athleteid="2489" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="2497" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" clubid="2818" name="Uczniowski Klub Sportowy Wodnik 29 Katowice">
          <CONTACT name="Skoczylas" phone="662297707" />
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Koenig" birthdate="1987-04-21" gender="F" nation="POL" athleteid="2824">
              <RESULTS>
                <RESULT eventid="1059" points="82" reactiontime="+80" swimtime="00:00:59.91" resultid="2825" heatid="4268" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1233" status="DNS" swimtime="00:00:00.00" resultid="2826" heatid="4327" lane="8" entrytime="00:04:40.00" />
                <RESULT eventid="1404" points="177" reactiontime="+84" swimtime="00:02:08.86" resultid="2827" heatid="4364" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="171" reactiontime="+92" swimtime="00:00:58.91" resultid="2828" heatid="4439" lane="3" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Mroziński" birthdate="1959-12-28" gender="M" nation="POL" swrid="4877351" athleteid="2819">
              <RESULTS>
                <RESULT eventid="1076" points="452" reactiontime="+82" swimtime="00:00:32.87" resultid="2820" heatid="4279" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1250" points="546" reactiontime="+92" swimtime="00:03:15.98" resultid="2821" heatid="4332" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                    <SPLIT distance="100" swimtime="00:01:33.39" />
                    <SPLIT distance="150" swimtime="00:02:25.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="594" reactiontime="+82" swimtime="00:01:25.30" resultid="2822" heatid="4369" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="724" reactiontime="+79" swimtime="00:00:36.52" resultid="2823" heatid="4447" lane="8" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ilnicki" birthdate="1956-03-22" gender="M" nation="POL" athleteid="2829">
              <RESULTS>
                <RESULT eventid="1112" status="DNS" swimtime="00:00:00.00" resultid="2830" heatid="4292" lane="4" entrytime="00:04:00.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="2831" heatid="4368" lane="9" entrytime="00:01:46.00" />
                <RESULT eventid="1697" status="DNS" swimtime="00:00:00.00" resultid="2832" heatid="4444" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3152" name="SMT Szczecin">
          <CONTACT email="kamila.gebka@gmail.com" name="Robert Zając" phone="501186428" />
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Moskalenko" birthdate="2000-12-01" gender="F" nation="POL" athleteid="3163">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+71" swimtime="00:00:34.06" resultid="3164" heatid="4271" lane="0" entrytime="00:00:32.80" />
                <RESULT eventid="1146" reactiontime="+77" swimtime="00:13:02.05" resultid="3165" heatid="4300" lane="2" entrytime="00:12:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:25.05" />
                    <SPLIT distance="150" swimtime="00:02:12.83" />
                    <SPLIT distance="200" swimtime="00:03:00.91" />
                    <SPLIT distance="250" swimtime="00:03:51.01" />
                    <SPLIT distance="300" swimtime="00:04:40.63" />
                    <SPLIT distance="350" swimtime="00:05:30.63" />
                    <SPLIT distance="400" swimtime="00:06:21.16" />
                    <SPLIT distance="450" swimtime="00:07:12.01" />
                    <SPLIT distance="500" swimtime="00:08:03.06" />
                    <SPLIT distance="550" swimtime="00:08:53.44" />
                    <SPLIT distance="600" swimtime="00:09:44.12" />
                    <SPLIT distance="650" swimtime="00:10:34.48" />
                    <SPLIT distance="700" swimtime="00:11:24.29" />
                    <SPLIT distance="750" swimtime="00:12:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" reactiontime="+74" swimtime="00:01:16.73" resultid="3166" heatid="4338" lane="2" entrytime="00:01:20.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" reactiontime="+75" swimtime="00:02:53.14" resultid="3167" heatid="4398" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:21.35" />
                    <SPLIT distance="150" swimtime="00:02:09.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Kramek" birthdate="1992-02-04" gender="M" nation="POL" athleteid="3158">
              <RESULTS>
                <RESULT eventid="1076" points="593" reactiontime="+72" swimtime="00:00:26.34" resultid="3159" heatid="4283" lane="4" entrytime="00:00:27.20" />
                <RESULT eventid="1301" points="529" reactiontime="+78" swimtime="00:01:01.58" resultid="3160" heatid="4350" lane="2" entrytime="00:00:59.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="479" reactiontime="+81" swimtime="00:00:29.73" resultid="3161" heatid="4382" lane="1" entrytime="00:00:29.90" />
                <RESULT eventid="1697" points="523" reactiontime="+74" swimtime="00:00:34.70" resultid="3162" heatid="4447" lane="1" entrytime="00:00:35.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iwona" lastname="Damljanovic Waclawik" birthdate="1965-04-21" gender="F" nation="POL" athleteid="3183">
              <RESULTS>
                <RESULT eventid="1094" points="308" reactiontime="+91" swimtime="00:03:44.46" resultid="3184" heatid="4288" lane="4" entrytime="00:03:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                    <SPLIT distance="100" swimtime="00:01:49.10" />
                    <SPLIT distance="150" swimtime="00:02:51.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="319" reactiontime="+97" swimtime="00:14:16.15" resultid="3185" heatid="4300" lane="1" entrytime="00:13:15.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:38.82" />
                    <SPLIT distance="150" swimtime="00:02:32.16" />
                    <SPLIT distance="200" swimtime="00:03:26.49" />
                    <SPLIT distance="250" swimtime="00:04:20.23" />
                    <SPLIT distance="300" swimtime="00:05:14.44" />
                    <SPLIT distance="350" swimtime="00:06:08.45" />
                    <SPLIT distance="400" swimtime="00:07:02.99" />
                    <SPLIT distance="450" swimtime="00:07:57.73" />
                    <SPLIT distance="500" swimtime="00:08:52.54" />
                    <SPLIT distance="550" swimtime="00:09:46.62" />
                    <SPLIT distance="600" swimtime="00:10:41.94" />
                    <SPLIT distance="650" swimtime="00:11:35.85" />
                    <SPLIT distance="700" swimtime="00:12:30.59" />
                    <SPLIT distance="750" swimtime="00:13:24.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="476" reactiontime="+94" swimtime="00:03:49.07" resultid="3186" heatid="4327" lane="3" entrytime="00:03:45.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.08" />
                    <SPLIT distance="100" swimtime="00:01:51.21" />
                    <SPLIT distance="150" swimtime="00:02:50.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="401" reactiontime="+92" swimtime="00:01:48.35" resultid="3187" heatid="4364" lane="3" entrytime="00:01:42.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="403" reactiontime="+86" swimtime="00:00:48.67" resultid="3188" heatid="4440" lane="4" entrytime="00:00:47.50" />
                <RESULT eventid="1731" points="308" swimtime="00:06:59.56" resultid="3189" heatid="4453" lane="9" entrytime="00:06:50.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.19" />
                    <SPLIT distance="100" swimtime="00:01:37.02" />
                    <SPLIT distance="150" swimtime="00:02:30.63" />
                    <SPLIT distance="200" swimtime="00:03:24.14" />
                    <SPLIT distance="250" swimtime="00:04:18.94" />
                    <SPLIT distance="300" swimtime="00:05:13.36" />
                    <SPLIT distance="350" swimtime="00:06:07.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Rożek" birthdate="1984-05-09" gender="M" nation="POL" athleteid="3173">
              <RESULTS>
                <RESULT eventid="1163" points="227" reactiontime="+88" swimtime="00:13:37.65" resultid="3175" heatid="4306" lane="4" entrytime="00:13:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:32.50" />
                    <SPLIT distance="150" swimtime="00:02:23.29" />
                    <SPLIT distance="200" swimtime="00:03:14.67" />
                    <SPLIT distance="250" swimtime="00:04:06.19" />
                    <SPLIT distance="300" swimtime="00:04:58.91" />
                    <SPLIT distance="350" swimtime="00:05:51.80" />
                    <SPLIT distance="400" swimtime="00:06:44.37" />
                    <SPLIT distance="450" swimtime="00:07:36.42" />
                    <SPLIT distance="500" swimtime="00:08:28.87" />
                    <SPLIT distance="550" swimtime="00:09:21.21" />
                    <SPLIT distance="600" swimtime="00:10:13.70" />
                    <SPLIT distance="650" swimtime="00:11:05.57" />
                    <SPLIT distance="700" swimtime="00:11:57.91" />
                    <SPLIT distance="750" swimtime="00:12:48.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="313" reactiontime="+82" swimtime="00:01:14.83" resultid="3176" heatid="4345" lane="5" entrytime="00:01:17.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="264" reactiontime="+82" swimtime="00:02:55.89" resultid="3177" heatid="4402" lane="7" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:02:55.89" />
                    <SPLIT distance="150" swimtime="00:02:11.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="247" reactiontime="+86" swimtime="00:06:31.75" resultid="4240" heatid="4460" lane="8" entrytime="00:06:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:01:29.13" />
                    <SPLIT distance="250" swimtime="00:04:01.28" />
                    <SPLIT distance="300" swimtime="00:04:53.08" />
                    <SPLIT distance="350" swimtime="00:05:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="262" reactiontime="+77" swimtime="00:00:37.71" resultid="4241" heatid="4379" lane="4" entrytime="00:00:39.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Kotowska" birthdate="1994-08-12" gender="F" nation="POL" athleteid="3153">
              <RESULTS>
                <RESULT eventid="1059" points="377" reactiontime="+89" swimtime="00:00:35.19" resultid="3154" heatid="4269" lane="6" entrytime="00:00:38.02" />
                <RESULT eventid="1215" points="230" reactiontime="+68" swimtime="00:00:46.33" resultid="3155" heatid="4315" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1284" points="359" reactiontime="+81" swimtime="00:01:20.13" resultid="3156" heatid="4338" lane="7" entrytime="00:01:21.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="208" reactiontime="+70" swimtime="00:01:43.90" resultid="3157" heatid="4387" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="240" reactiontime="+86" swimtime="00:06:56.26" resultid="5105" heatid="4455" lane="5" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:29.82" />
                    <SPLIT distance="150" swimtime="00:02:21.40" />
                    <SPLIT distance="200" swimtime="00:03:15.90" />
                    <SPLIT distance="250" swimtime="00:04:11.06" />
                    <SPLIT distance="300" swimtime="00:05:07.02" />
                    <SPLIT distance="350" swimtime="00:06:03.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Zieliński" birthdate="1992-09-02" gender="M" nation="POL" athleteid="3179">
              <RESULTS>
                <RESULT eventid="1076" points="723" reactiontime="+72" swimtime="00:00:24.66" resultid="3180" heatid="4285" lane="5" entrytime="00:00:26.02" />
                <RESULT eventid="1301" points="771" reactiontime="+76" swimtime="00:00:54.32" resultid="3181" heatid="4352" lane="1" entrytime="00:00:55.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="641" reactiontime="+75" swimtime="00:00:26.98" resultid="3182" heatid="4383" lane="1" entrytime="00:00:28.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Zając" birthdate="1966-06-30" gender="M" nation="POL" athleteid="3168">
              <RESULTS>
                <RESULT eventid="1076" points="460" reactiontime="+91" swimtime="00:00:31.68" resultid="3169" heatid="4278" lane="4" entrytime="00:00:32.30" />
                <RESULT eventid="1301" points="410" reactiontime="+99" swimtime="00:01:15.38" resultid="3170" heatid="4346" lane="0" entrytime="00:01:15.02" />
                <RESULT eventid="1457" points="439" reactiontime="+95" swimtime="00:00:34.95" resultid="3171" heatid="4380" lane="2" entrytime="00:00:34.80" />
                <RESULT eventid="1697" status="DNS" swimtime="00:00:00.00" resultid="3172" heatid="4445" lane="1" entrytime="00:00:41.20" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1386" points="469" reactiontime="+87" swimtime="00:02:11.68" resultid="3191" heatid="4491" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="150" swimtime="00:01:39.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3179" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3158" number="2" />
                    <RELAYPOSITION athleteid="3168" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3173" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" points="552" reactiontime="+78" swimtime="00:01:53.18" resultid="3192" heatid="4496" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.10" />
                    <SPLIT distance="100" swimtime="00:00:56.85" />
                    <SPLIT distance="150" swimtime="00:01:28.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3158" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3168" number="2" />
                    <RELAYPOSITION athleteid="3173" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="3179" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" points="394" reactiontime="+84" swimtime="00:02:19.45" resultid="3190" heatid="4489" lane="7" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="150" swimtime="00:01:48.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3173" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3183" number="2" />
                    <RELAYPOSITION athleteid="3153" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="3168" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1714" points="354" reactiontime="+87" swimtime="00:02:40.04" resultid="3193" heatid="4498" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:28.32" />
                    <SPLIT distance="150" swimtime="00:02:05.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3168" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3183" number="2" />
                    <RELAYPOSITION athleteid="3173" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="3153" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" clubid="3468" name="Ks Extreme Team Oborniki">
          <CONTACT city="OBORNIKI" email="JANWOL2212@GMAIL.COM" name="WOLNIEWICZ" phone="791064667" state="WIE" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Wolniewicz" birthdate="1948-12-22" gender="M" nation="POL" swrid="4754624" athleteid="3469">
              <RESULTS>
                <RESULT eventid="1076" points="361" reactiontime="+83" swimtime="00:00:38.93" resultid="3470" heatid="4277" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1197" points="245" reactiontime="+98" swimtime="00:32:39.01" resultid="3471" heatid="4310" lane="0" entrytime="00:30:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.75" />
                    <SPLIT distance="100" swimtime="00:01:53.43" />
                    <SPLIT distance="150" swimtime="00:02:55.57" />
                    <SPLIT distance="200" swimtime="00:04:00.66" />
                    <SPLIT distance="250" swimtime="00:05:03.85" />
                    <SPLIT distance="300" swimtime="00:06:08.62" />
                    <SPLIT distance="350" swimtime="00:07:13.84" />
                    <SPLIT distance="400" swimtime="00:08:17.65" />
                    <SPLIT distance="450" swimtime="00:09:23.32" />
                    <SPLIT distance="500" swimtime="00:10:29.44" />
                    <SPLIT distance="550" swimtime="00:11:34.86" />
                    <SPLIT distance="600" swimtime="00:12:41.24" />
                    <SPLIT distance="650" swimtime="00:13:46.48" />
                    <SPLIT distance="700" swimtime="00:14:51.84" />
                    <SPLIT distance="750" swimtime="00:15:58.86" />
                    <SPLIT distance="800" swimtime="00:17:07.25" />
                    <SPLIT distance="850" swimtime="00:18:11.76" />
                    <SPLIT distance="900" swimtime="00:19:18.81" />
                    <SPLIT distance="950" swimtime="00:20:24.67" />
                    <SPLIT distance="1000" swimtime="00:21:31.26" />
                    <SPLIT distance="1050" swimtime="00:22:37.48" />
                    <SPLIT distance="1100" swimtime="00:23:46.79" />
                    <SPLIT distance="1150" swimtime="00:24:52.56" />
                    <SPLIT distance="1200" swimtime="00:25:59.36" />
                    <SPLIT distance="1250" swimtime="00:27:06.58" />
                    <SPLIT distance="1300" swimtime="00:28:14.39" />
                    <SPLIT distance="1350" swimtime="00:29:21.22" />
                    <SPLIT distance="1400" swimtime="00:30:28.99" />
                    <SPLIT distance="1450" swimtime="00:31:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="315" reactiontime="+94" swimtime="00:01:33.06" resultid="3472" heatid="4344" lane="6" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="3473" heatid="4378" lane="3" entrytime="00:00:54.00" />
                <RESULT eventid="1525" points="243" reactiontime="+96" swimtime="00:03:49.60" resultid="3474" heatid="4401" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.85" />
                    <SPLIT distance="100" swimtime="00:01:49.93" />
                    <SPLIT distance="150" swimtime="00:02:52.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="226" reactiontime="+93" swimtime="00:08:18.57" resultid="3475" heatid="4461" lane="0" entrytime="00:07:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.48" />
                    <SPLIT distance="200" swimtime="00:04:00.07" />
                    <SPLIT distance="300" swimtime="00:06:09.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06306" nation="POL" region="06" clubid="2047" name="Ks Korona 1919">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Orlewicz- Musiał" birthdate="1960-05-29" gender="F" nation="POL" license="506306600054" swrid="5352178" athleteid="2108">
              <RESULTS>
                <RESULT eventid="1094" points="179" reactiontime="+106" swimtime="00:04:52.04" resultid="2109" heatid="4287" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.65" />
                    <SPLIT distance="100" swimtime="00:02:16.06" />
                    <SPLIT distance="150" swimtime="00:03:45.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="181" swimtime="00:35:08.19" resultid="2110" heatid="4308" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.65" />
                    <SPLIT distance="100" swimtime="00:01:57.74" />
                    <SPLIT distance="150" swimtime="00:03:04.21" />
                    <SPLIT distance="200" swimtime="00:04:11.67" />
                    <SPLIT distance="250" swimtime="00:05:20.05" />
                    <SPLIT distance="300" swimtime="00:06:28.93" />
                    <SPLIT distance="350" swimtime="00:07:40.00" />
                    <SPLIT distance="400" swimtime="00:08:49.72" />
                    <SPLIT distance="450" swimtime="00:10:00.50" />
                    <SPLIT distance="500" swimtime="00:11:09.58" />
                    <SPLIT distance="550" swimtime="00:12:19.61" />
                    <SPLIT distance="600" swimtime="00:13:29.49" />
                    <SPLIT distance="650" swimtime="00:14:39.55" />
                    <SPLIT distance="700" swimtime="00:15:49.84" />
                    <SPLIT distance="750" swimtime="00:16:59.69" />
                    <SPLIT distance="800" swimtime="00:18:09.41" />
                    <SPLIT distance="850" swimtime="00:19:20.12" />
                    <SPLIT distance="900" swimtime="00:20:32.11" />
                    <SPLIT distance="950" swimtime="00:21:44.02" />
                    <SPLIT distance="1000" swimtime="00:22:55.75" />
                    <SPLIT distance="1050" swimtime="00:24:07.27" />
                    <SPLIT distance="1100" swimtime="00:25:20.17" />
                    <SPLIT distance="1150" swimtime="00:26:34.28" />
                    <SPLIT distance="1200" swimtime="00:27:47.25" />
                    <SPLIT distance="1250" swimtime="00:28:59.78" />
                    <SPLIT distance="1300" swimtime="00:30:12.83" />
                    <SPLIT distance="1350" swimtime="00:31:29.19" />
                    <SPLIT distance="1400" swimtime="00:32:43.28" />
                    <SPLIT distance="1450" swimtime="00:33:58.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="155" reactiontime="+86" swimtime="00:01:02.98" resultid="2111" heatid="4313" lane="5" entrytime="00:01:03.81" entrycourse="LCM" />
                <RESULT eventid="1335" points="113" reactiontime="+111" swimtime="00:05:32.88" resultid="2112" heatid="4353" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.45" />
                    <SPLIT distance="100" swimtime="00:02:29.48" />
                    <SPLIT distance="150" swimtime="00:04:01.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="115" swimtime="00:01:03.95" resultid="2113" heatid="4373" lane="9" />
                <RESULT eventid="1576" points="180" reactiontime="+104" swimtime="00:10:30.65" resultid="2114" heatid="4413" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.09" />
                    <SPLIT distance="100" swimtime="00:02:34.30" />
                    <SPLIT distance="150" swimtime="00:03:51.65" />
                    <SPLIT distance="200" swimtime="00:05:11.19" />
                    <SPLIT distance="250" swimtime="00:06:40.67" />
                    <SPLIT distance="300" swimtime="00:08:11.38" />
                    <SPLIT distance="350" swimtime="00:09:20.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="158" reactiontime="+80" swimtime="00:04:58.60" resultid="2115" heatid="4428" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.88" />
                    <SPLIT distance="100" swimtime="00:02:25.34" />
                    <SPLIT distance="150" swimtime="00:03:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="165" swimtime="00:09:06.78" resultid="2116" heatid="4454" lane="7" entrytime="00:08:35.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.38" />
                    <SPLIT distance="100" swimtime="00:02:02.56" />
                    <SPLIT distance="150" swimtime="00:03:12.25" />
                    <SPLIT distance="200" swimtime="00:04:21.09" />
                    <SPLIT distance="250" swimtime="00:05:32.17" />
                    <SPLIT distance="300" swimtime="00:06:43.47" />
                    <SPLIT distance="350" swimtime="00:07:57.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Waldemar" lastname="Piszczek" birthdate="1962-11-10" gender="M" nation="POL" license="506306700055" swrid="4992814" athleteid="2085">
              <RESULTS>
                <RESULT eventid="1076" points="548" reactiontime="+89" swimtime="00:00:30.84" resultid="2086" heatid="4274" lane="5" />
                <RESULT eventid="1112" status="DNS" swimtime="00:00:00.00" resultid="2087" heatid="4292" lane="8" />
                <RESULT eventid="1267" points="643" reactiontime="+81" swimtime="00:00:35.44" resultid="2088" heatid="4319" lane="1" />
                <RESULT eventid="1250" points="542" reactiontime="+96" swimtime="00:03:16.42" resultid="2089" heatid="4330" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="100" swimtime="00:01:32.66" />
                    <SPLIT distance="150" swimtime="00:02:26.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1457" points="701" reactiontime="+91" swimtime="00:00:31.13" resultid="2090" heatid="4377" lane="2" />
                <RESULT eventid="1491" points="580" reactiontime="+79" swimtime="00:01:19.23" resultid="2091" heatid="4389" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="2092" heatid="4423" lane="9" />
                <RESULT eventid="1663" points="564" reactiontime="+76" swimtime="00:02:56.85" resultid="2093" heatid="4432" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:24.30" />
                    <SPLIT distance="150" swimtime="00:02:12.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Leńczowska" birthdate="1982-01-15" gender="F" nation="POL" license="506306600071" swrid="4992907" athleteid="2055">
              <RESULTS>
                <RESULT eventid="1059" points="606" reactiontime="+85" swimtime="00:00:31.24" resultid="2056" heatid="4271" lane="9" entrytime="00:00:33.99" entrycourse="LCM" />
                <RESULT eventid="1094" points="560" reactiontime="+92" swimtime="00:02:56.00" resultid="2057" heatid="4288" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:23.68" />
                    <SPLIT distance="150" swimtime="00:02:14.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="527" reactiontime="+66" swimtime="00:00:36.68" resultid="2058" heatid="4315" lane="2" entrytime="00:00:38.42" entrycourse="LCM" />
                <RESULT eventid="1284" points="483" reactiontime="+82" swimtime="00:01:13.99" resultid="2059" heatid="4335" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="530" reactiontime="+79" swimtime="00:00:35.04" resultid="2060" heatid="4372" lane="7" />
                <RESULT eventid="1474" points="472" reactiontime="+81" swimtime="00:01:23.07" resultid="2061" heatid="4388" lane="8" entrytime="00:01:23.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="505" reactiontime="+70" swimtime="00:02:59.84" resultid="2062" heatid="4431" lane="8" entrytime="00:03:09.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:28.95" />
                    <SPLIT distance="150" swimtime="00:02:16.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="450" reactiontime="+94" swimtime="00:00:42.36" resultid="2063" heatid="4438" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariola" lastname="Kuliś" birthdate="1966-07-27" gender="F" nation="POL" license="506306600043" swrid="4992797" athleteid="2048">
              <RESULTS>
                <RESULT eventid="1059" points="731" reactiontime="+72" swimtime="00:00:31.40" resultid="2049" heatid="4271" lane="7" entrytime="00:00:31.92" entrycourse="LCM" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1215" points="618" reactiontime="+69" swimtime="00:00:37.56" resultid="2050" heatid="4315" lane="3" entrytime="00:00:37.83" entrycourse="LCM" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1284" points="636" reactiontime="+77" swimtime="00:01:12.10" resultid="2051" heatid="4336" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="669" reactiontime="+79" swimtime="00:01:31.35" resultid="2052" heatid="4364" lane="5" entrytime="00:01:41.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1474" points="565" reactiontime="+83" swimtime="00:01:24.28" resultid="2053" heatid="4388" lane="9" entrytime="00:01:25.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="750" reactiontime="+80" swimtime="00:00:39.55" resultid="2054" heatid="4441" lane="8" entrytime="00:00:40.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogusław" lastname="Kwiatkowski" birthdate="1956-07-24" gender="M" nation="POL" license="506306700044" swrid="5468084" athleteid="2078">
              <RESULTS>
                <RESULT comment="O11" eventid="1076" reactiontime="+116" status="DSQ" swimtime="00:00:00.00" resultid="2079" heatid="4275" lane="4" entrytime="00:00:52.70" entrycourse="LCM" />
                <RESULT eventid="1267" points="125" reactiontime="+94" swimtime="00:01:01.92" resultid="2080" heatid="4320" lane="7" entrytime="00:01:02.52" entrycourse="LCM" />
                <RESULT eventid="1301" points="124" reactiontime="+110" swimtime="00:01:59.22" resultid="2081" heatid="4344" lane="9" entrytime="00:02:05.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="92" reactiontime="+105" swimtime="00:02:45.39" resultid="2082" heatid="4367" lane="1" entrytime="00:02:37.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="97" reactiontime="+113" swimtime="00:04:41.14" resultid="2083" heatid="4399" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.27" />
                    <SPLIT distance="100" swimtime="00:02:11.26" />
                    <SPLIT distance="150" swimtime="00:03:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="106" reactiontime="+116" swimtime="00:01:10.28" resultid="2084" heatid="4443" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Zygmuntowicz" birthdate="1982-10-17" gender="F" nation="POL" license="506306600077" athleteid="2071">
              <RESULTS>
                <RESULT eventid="1059" points="509" reactiontime="+82" swimtime="00:00:33.12" resultid="2072" heatid="4266" lane="4" />
                <RESULT eventid="1094" points="444" reactiontime="+73" swimtime="00:03:10.04" resultid="2073" heatid="4287" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:29.18" />
                    <SPLIT distance="150" swimtime="00:02:26.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="424" reactiontime="+86" swimtime="00:01:17.26" resultid="2074" heatid="4335" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="488" reactiontime="+82" swimtime="00:00:36.02" resultid="2075" heatid="4372" lane="5" />
                <RESULT eventid="1508" points="432" reactiontime="+88" swimtime="00:02:51.08" resultid="2076" heatid="4395" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="100" swimtime="00:01:24.18" />
                    <SPLIT distance="150" swimtime="00:02:10.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="414" reactiontime="+89" swimtime="00:01:25.02" resultid="2077" heatid="4419" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" license="506306600048" swrid="4992827" athleteid="2099">
              <RESULTS>
                <RESULT eventid="1094" points="558" swimtime="00:03:19.93" resultid="2100" heatid="4289" lane="7" entrytime="00:03:18.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:01:35.66" />
                    <SPLIT distance="150" swimtime="00:02:36.56" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1146" points="510" swimtime="00:13:05.71" resultid="2101" heatid="4302" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="150" swimtime="00:02:19.07" />
                    <SPLIT distance="250" swimtime="00:03:58.86" />
                    <SPLIT distance="350" swimtime="00:05:39.47" />
                    <SPLIT distance="450" swimtime="00:07:20.07" />
                    <SPLIT distance="550" swimtime="00:09:00.58" />
                    <SPLIT distance="650" swimtime="00:10:40.66" />
                    <SPLIT distance="750" swimtime="00:12:20.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="541" reactiontime="+102" swimtime="00:01:18.35" resultid="2102" heatid="4338" lane="3" entrytime="00:01:20.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1335" points="427" swimtime="00:03:33.84" resultid="2103" heatid="4353" lane="4" entrytime="00:03:30.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                    <SPLIT distance="100" swimtime="00:01:38.63" />
                    <SPLIT distance="150" swimtime="00:02:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="480" reactiontime="+82" swimtime="00:01:35.13" resultid="2104" heatid="4385" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1508" points="521" swimtime="00:02:55.26" resultid="2105" heatid="4397" lane="4" entrytime="00:02:55.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:26.14" />
                    <SPLIT distance="150" swimtime="00:02:12.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="443" reactiontime="+92" swimtime="00:01:34.50" resultid="2106" heatid="4420" lane="3" entrytime="00:01:32.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="493" swimtime="00:06:19.57" resultid="2107" heatid="4455" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                    <SPLIT distance="100" swimtime="00:01:28.30" />
                    <SPLIT distance="150" swimtime="00:02:17.37" />
                    <SPLIT distance="200" swimtime="00:03:06.17" />
                    <SPLIT distance="250" swimtime="00:03:55.72" />
                    <SPLIT distance="300" swimtime="00:04:44.93" />
                    <SPLIT distance="350" swimtime="00:05:33.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Bielańska" birthdate="1984-04-20" gender="F" nation="POL" license="506306600072" swrid="5468078" athleteid="2064">
              <RESULTS>
                <RESULT eventid="1059" points="144" reactiontime="+114" swimtime="00:00:49.53" resultid="2065" heatid="4268" lane="8" />
                <RESULT eventid="1215" points="151" reactiontime="+96" swimtime="00:00:53.77" resultid="2066" heatid="4314" lane="8" entrytime="00:00:53.99" entrycourse="LCM" />
                <RESULT eventid="1233" points="145" reactiontime="+105" swimtime="00:04:55.76" resultid="2067" heatid="4326" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.93" />
                    <SPLIT distance="100" swimtime="00:02:25.73" />
                    <SPLIT distance="150" swimtime="00:03:43.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="131" reactiontime="+101" swimtime="00:02:22.44" resultid="2068" heatid="4362" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="133" reactiontime="+109" swimtime="00:02:00.95" resultid="2069" heatid="4386" lane="0" />
                <RESULT eventid="1680" points="149" reactiontime="+102" swimtime="00:01:01.63" resultid="2070" heatid="4438" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Borek" birthdate="1991-01-01" gender="M" nation="POL" license="506306700069" swrid="5468079" athleteid="2117">
              <RESULTS>
                <RESULT eventid="1267" points="467" reactiontime="+62" swimtime="00:00:33.48" resultid="2118" heatid="4319" lane="5" />
                <RESULT eventid="1491" points="426" reactiontime="+62" swimtime="00:01:14.36" resultid="2119" heatid="4392" lane="4" entrytime="00:01:17.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="395" reactiontime="+73" swimtime="00:00:38.09" resultid="2120" heatid="4446" lane="9" entrytime="00:00:38.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Baranik" birthdate="1969-06-29" gender="M" nation="POL" license="506306700027" swrid="4992740" athleteid="2094">
              <RESULTS>
                <RESULT eventid="1076" points="713" reactiontime="+74" swimtime="00:00:26.95" resultid="2095" heatid="4284" lane="1" entrytime="00:00:27.02" entrycourse="LCM" />
                <RESULT eventid="1301" points="672" reactiontime="+75" swimtime="00:01:01.81" resultid="2096" heatid="4349" lane="3" entrytime="00:01:01.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="727" reactiontime="+70" swimtime="00:00:28.78" resultid="2097" heatid="4382" lane="5" entrytime="00:00:29.15" entrycourse="LCM" />
                <RESULT eventid="1697" points="661" reactiontime="+74" swimtime="00:00:34.62" resultid="2098" heatid="4448" lane="2" entrytime="00:00:33.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1386" points="410" reactiontime="+64" swimtime="00:02:29.22" resultid="2122" heatid="4492" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:10.03" />
                    <SPLIT distance="150" swimtime="00:01:38.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2117" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2085" number="2" />
                    <RELAYPOSITION athleteid="2094" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2078" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1542" points="541" reactiontime="+78" swimtime="00:02:13.05" resultid="2123" heatid="4494" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:07.12" />
                    <SPLIT distance="150" swimtime="00:01:41.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2048" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="2099" number="2" />
                    <RELAYPOSITION athleteid="2071" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="2055" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" points="672" reactiontime="+77" swimtime="00:01:59.86" resultid="2121" heatid="4488" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:01.19" />
                    <SPLIT distance="150" swimtime="00:01:33.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2048" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2085" number="2" />
                    <RELAYPOSITION athleteid="2055" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="2094" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1714" points="530" reactiontime="+87" swimtime="00:02:19.93" resultid="2124" heatid="4498" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:18.26" />
                    <SPLIT distance="150" swimtime="00:01:49.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2055" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="2048" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2071" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2099" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3220" name="Gdynia Masters">
          <CONTACT name="Mysiak" />
          <ATHLETES>
            <ATHLETE firstname="Jan Maciej" lastname="Boboli" birthdate="1948-01-01" gender="M" nation="POL" swrid="4754700" athleteid="3226">
              <RESULTS>
                <RESULT eventid="1076" points="367" reactiontime="+85" swimtime="00:00:38.70" resultid="3227" heatid="4276" lane="4" entrytime="00:00:39.38" entrycourse="LCM" />
                <RESULT eventid="1301" points="237" reactiontime="+87" swimtime="00:01:42.38" resultid="3228" heatid="4344" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="180" reactiontime="+88" swimtime="00:00:53.11" resultid="3229" heatid="4378" lane="2" entrytime="00:00:59.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grażyna" lastname="Heisler" birthdate="1951-01-01" gender="F" nation="POL" swrid="4191114" athleteid="3241">
              <RESULTS>
                <RESULT eventid="1059" points="324" reactiontime="+100" swimtime="00:00:44.75" resultid="3242" heatid="4267" lane="2" />
                <RESULT eventid="1404" points="324" reactiontime="+108" swimtime="00:02:19.70" resultid="3243" heatid="4363" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="191" reactiontime="+86" swimtime="00:02:15.41" resultid="3244" heatid="4386" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="318" reactiontime="+109" swimtime="00:01:01.03" resultid="3245" heatid="4438" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Chomicka" birthdate="1952-01-01" gender="F" nation="POL" swrid="4302084" athleteid="3238">
              <RESULTS>
                <RESULT eventid="1059" points="113" swimtime="00:01:03.54" resultid="3239" heatid="4268" lane="1" />
                <RESULT eventid="1215" points="154" reactiontime="+77" swimtime="00:01:04.70" resultid="3240" heatid="4312" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Skwarło" birthdate="1939-01-01" gender="M" nation="POL" swrid="4302086" athleteid="3230">
              <RESULTS>
                <RESULT eventid="1076" points="229" reactiontime="+101" swimtime="00:00:52.21" resultid="3231" heatid="4275" lane="5" entrytime="00:00:54.50" />
                <RESULT eventid="1112" points="403" reactiontime="+113" swimtime="00:04:29.23" resultid="3232" heatid="4292" lane="1" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.82" />
                    <SPLIT distance="100" swimtime="00:02:59.52" />
                    <SPLIT distance="150" swimtime="00:04:22.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="225" reactiontime="+104" swimtime="00:01:02.74" resultid="3233" heatid="4320" lane="1" entrytime="00:01:03.30" entrycourse="LCM" />
                <RESULT eventid="1250" points="312" reactiontime="+102" swimtime="00:05:06.37" resultid="3234" heatid="4330" lane="4" entrytime="00:04:52.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.99" />
                    <SPLIT distance="100" swimtime="00:02:27.21" />
                    <SPLIT distance="150" swimtime="00:03:49.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="317" reactiontime="+95" swimtime="00:02:18.47" resultid="3235" heatid="4367" lane="7" entrytime="00:02:20.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="184" reactiontime="+111" swimtime="00:02:32.08" resultid="3236" heatid="4390" lane="8" entrytime="00:02:28.07" entrycourse="LCM" />
                <RESULT eventid="1697" points="384" reactiontime="+98" swimtime="00:00:57.32" resultid="3237" heatid="4443" lane="5" entrytime="00:00:55.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Mysiak" birthdate="1961-01-01" gender="F" nation="POL" swrid="4754669" athleteid="3221">
              <RESULTS>
                <RESULT eventid="1474" points="290" reactiontime="+88" swimtime="00:01:52.56" resultid="3222" heatid="4387" lane="6" entrytime="00:01:40.00" />
                <RESULT eventid="1508" points="269" reactiontime="+99" swimtime="00:03:38.40" resultid="3223" heatid="4396" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                    <SPLIT distance="100" swimtime="00:01:44.11" />
                    <SPLIT distance="150" swimtime="00:02:43.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="307" reactiontime="+89" swimtime="00:03:59.44" resultid="3224" heatid="4430" lane="1" entrytime="00:03:57.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="286" reactiontime="+101" swimtime="00:07:35.10" resultid="3225" heatid="4453" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                    <SPLIT distance="100" swimtime="00:01:42.42" />
                    <SPLIT distance="150" swimtime="00:02:40.16" />
                    <SPLIT distance="200" swimtime="00:03:39.76" />
                    <SPLIT distance="250" swimtime="00:04:39.18" />
                    <SPLIT distance="300" swimtime="00:05:39.35" />
                    <SPLIT distance="350" swimtime="00:06:39.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" swimtime="00:03:27.30" resultid="3246" heatid="4488" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.79" />
                    <SPLIT distance="100" swimtime="00:02:02.80" />
                    <SPLIT distance="150" swimtime="00:02:47.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3226" number="1" />
                    <RELAYPOSITION athleteid="3238" number="2" />
                    <RELAYPOSITION athleteid="3241" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="3230" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1714" reactiontime="+87" swimtime="00:03:21.16" resultid="3247" heatid="4498" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.60" />
                    <SPLIT distance="100" swimtime="00:01:47.98" />
                    <SPLIT distance="150" swimtime="00:02:36.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3241" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3230" number="2" />
                    <RELAYPOSITION athleteid="3226" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3221" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="10414" nation="POL" region="14" clubid="1938" name="Klub Sportowy Mako">
          <CONTACT city="Warszawa" email="ania.plywanie@gmail.com" name="Anna Dąbrowska" phone="601 480 280" />
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Safrończyk" birthdate="1988-05-30" gender="M" nation="POL" swrid="4072743" athleteid="3712">
              <RESULTS>
                <RESULT eventid="1250" points="711" reactiontime="+65" swimtime="00:02:34.65" resultid="3713" heatid="4334" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="150" swimtime="00:01:53.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="761" reactiontime="+62" swimtime="00:01:07.10" resultid="3714" heatid="4371" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="856" reactiontime="+63" swimtime="00:00:29.44" resultid="3715" heatid="4449" lane="5" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Rurak" birthdate="1988-05-09" gender="M" nation="POL" swrid="4072773" athleteid="3710">
              <RESULTS>
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="3711" heatid="4303" lane="4" entrytime="00:08:59.43" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Dąbrowska" birthdate="1987-05-20" gender="F" nation="POL" license="510414600006" swrid="4655165" athleteid="1939">
              <RESULTS>
                <RESULT eventid="1059" points="286" reactiontime="+104" swimtime="00:00:39.44" resultid="1940" heatid="4269" lane="2" entrytime="00:00:39.38" entrycourse="LCM" />
                <RESULT eventid="1094" points="210" reactiontime="+108" swimtime="00:03:57.92" resultid="1941" heatid="4288" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.36" />
                    <SPLIT distance="100" swimtime="00:01:57.41" />
                    <SPLIT distance="150" swimtime="00:03:04.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="147" reactiontime="+113" swimtime="00:00:54.27" resultid="1942" heatid="4312" lane="8" />
                <RESULT eventid="1284" points="237" reactiontime="+112" swimtime="00:01:33.86" resultid="1943" heatid="4336" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="122" reactiontime="+99" swimtime="00:02:04.61" resultid="1944" heatid="4385" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="212" reactiontime="+108" swimtime="00:03:31.15" resultid="1945" heatid="4395" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.19" />
                    <SPLIT distance="100" swimtime="00:01:42.16" />
                    <SPLIT distance="150" swimtime="00:02:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="138" reactiontime="+95" swimtime="00:04:27.43" resultid="1946" heatid="4429" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.87" />
                    <SPLIT distance="150" swimtime="00:03:23.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="200" reactiontime="+109" swimtime="00:07:34.77" resultid="1947" heatid="4455" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.41" />
                    <SPLIT distance="100" swimtime="00:01:48.09" />
                    <SPLIT distance="150" swimtime="00:02:44.85" />
                    <SPLIT distance="200" swimtime="00:03:43.17" />
                    <SPLIT distance="250" swimtime="00:04:42.54" />
                    <SPLIT distance="300" swimtime="00:05:42.30" />
                    <SPLIT distance="350" swimtime="00:06:39.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Rudziński" birthdate="1966-05-10" gender="M" nation="POL" license="510414700010" swrid="4934041" athleteid="1972">
              <RESULTS>
                <RESULT eventid="1250" points="334" reactiontime="+114" swimtime="00:03:37.15" resultid="1973" heatid="4330" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.03" />
                    <SPLIT distance="100" swimtime="00:01:42.51" />
                    <SPLIT distance="150" swimtime="00:02:40.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="218" reactiontime="+104" swimtime="00:03:47.17" resultid="1974" heatid="4355" lane="2" entrytime="00:04:08.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:40.35" />
                    <SPLIT distance="150" swimtime="00:02:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="252" reactiontime="+102" swimtime="00:00:42.05" resultid="1975" heatid="4377" lane="4" />
                <RESULT eventid="1593" points="262" reactiontime="+116" swimtime="00:07:51.42" resultid="1976" heatid="4417" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                    <SPLIT distance="100" swimtime="00:04:05.70" />
                    <SPLIT distance="150" swimtime="00:02:58.38" />
                    <SPLIT distance="200" swimtime="00:06:02.96" />
                    <SPLIT distance="250" swimtime="00:05:02.46" />
                    <SPLIT distance="350" swimtime="00:06:57.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="219" reactiontime="+105" swimtime="00:01:40.50" resultid="1977" heatid="4423" lane="4" entrytime="00:01:43.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="161" reactiontime="+102" swimtime="00:04:18.93" resultid="1978" heatid="4432" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.70" />
                    <SPLIT distance="100" swimtime="00:02:07.80" />
                    <SPLIT distance="150" swimtime="00:03:16.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" license="510414700072" swrid="5506637" athleteid="1965">
              <RESULTS>
                <RESULT eventid="1267" points="229" reactiontime="+73" swimtime="00:00:47.48" resultid="1966" heatid="4318" lane="6" />
                <RESULT eventid="1301" points="224" reactiontime="+95" swimtime="00:01:32.22" resultid="1967" heatid="4342" lane="0" />
                <RESULT eventid="1491" points="178" reactiontime="+86" swimtime="00:01:52.91" resultid="1968" heatid="4389" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="182" reactiontime="+102" swimtime="00:03:38.69" resultid="1969" heatid="4400" lane="0">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="218" reactiontime="+94" swimtime="00:03:54.14" resultid="1970" heatid="4433" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.69" />
                    <SPLIT distance="100" swimtime="00:01:54.94" />
                    <SPLIT distance="150" swimtime="00:02:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="168" reactiontime="+94" swimtime="00:07:55.28" resultid="1971" heatid="4462" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.49" />
                    <SPLIT distance="100" swimtime="00:01:47.68" />
                    <SPLIT distance="150" swimtime="00:02:48.28" />
                    <SPLIT distance="200" swimtime="00:03:50.64" />
                    <SPLIT distance="250" swimtime="00:04:51.44" />
                    <SPLIT distance="300" swimtime="00:05:52.33" />
                    <SPLIT distance="350" swimtime="00:06:55.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" license="510414700009" swrid="4655152" athleteid="1948">
              <RESULTS>
                <RESULT eventid="1076" points="221" reactiontime="+86" swimtime="00:00:40.42" resultid="1949" heatid="4277" lane="9" entrytime="00:00:38.57" entrycourse="LCM" />
                <RESULT eventid="1250" status="DNS" swimtime="00:00:00.00" resultid="1950" heatid="4329" lane="1" />
                <RESULT eventid="1301" points="236" reactiontime="+73" swimtime="00:01:30.62" resultid="1951" heatid="4344" lane="3" entrytime="00:01:33.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="278" reactiontime="+70" swimtime="00:01:43.60" resultid="1952" heatid="4368" lane="0" entrytime="00:01:45.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="193" reactiontime="+73" swimtime="00:03:34.76" resultid="1953" heatid="4400" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:41.37" />
                    <SPLIT distance="100" swimtime="00:01:44.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="309" reactiontime="+73" swimtime="00:00:44.40" resultid="1954" heatid="4444" lane="5" entrytime="00:00:44.46" entrycourse="LCM" />
                <RESULT eventid="1748" points="185" reactiontime="+91" swimtime="00:07:40.87" resultid="1955" heatid="4461" lane="2" entrytime="00:07:15.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.70" />
                    <SPLIT distance="100" swimtime="00:01:49.40" />
                    <SPLIT distance="150" swimtime="00:02:50.65" />
                    <SPLIT distance="200" swimtime="00:03:51.28" />
                    <SPLIT distance="250" swimtime="00:04:50.49" />
                    <SPLIT distance="300" swimtime="00:05:48.49" />
                    <SPLIT distance="350" swimtime="00:06:46.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Domeracki" birthdate="1982-02-27" gender="M" nation="POL" athleteid="3716">
              <RESULTS>
                <RESULT eventid="1197" points="394" reactiontime="+83" swimtime="00:22:22.96" resultid="3717" heatid="4309" lane="0" entrytime="00:21:30.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:04.26" />
                    <SPLIT distance="200" swimtime="00:02:48.67" />
                    <SPLIT distance="250" swimtime="00:03:33.23" />
                    <SPLIT distance="300" swimtime="00:04:18.29" />
                    <SPLIT distance="350" swimtime="00:05:02.81" />
                    <SPLIT distance="400" swimtime="00:05:47.75" />
                    <SPLIT distance="450" swimtime="00:06:32.33" />
                    <SPLIT distance="500" swimtime="00:07:17.12" />
                    <SPLIT distance="550" swimtime="00:08:01.81" />
                    <SPLIT distance="600" swimtime="00:08:47.18" />
                    <SPLIT distance="650" swimtime="00:09:32.49" />
                    <SPLIT distance="700" swimtime="00:10:17.96" />
                    <SPLIT distance="750" swimtime="00:11:03.62" />
                    <SPLIT distance="800" swimtime="00:11:49.38" />
                    <SPLIT distance="850" swimtime="00:12:34.65" />
                    <SPLIT distance="900" swimtime="00:13:20.46" />
                    <SPLIT distance="950" swimtime="00:14:05.57" />
                    <SPLIT distance="1000" swimtime="00:14:51.29" />
                    <SPLIT distance="1050" swimtime="00:15:36.32" />
                    <SPLIT distance="1100" swimtime="00:16:22.07" />
                    <SPLIT distance="1150" swimtime="00:17:07.82" />
                    <SPLIT distance="1200" swimtime="00:17:53.05" />
                    <SPLIT distance="1250" swimtime="00:18:38.17" />
                    <SPLIT distance="1300" swimtime="00:19:23.64" />
                    <SPLIT distance="1350" swimtime="00:20:08.93" />
                    <SPLIT distance="1400" swimtime="00:20:54.35" />
                    <SPLIT distance="1450" swimtime="00:21:38.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michal" lastname="Gugała" birthdate="1979-01-13" gender="M" nation="POL" swrid="4992802" athleteid="3703">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3704" heatid="4279" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="3705" heatid="4305" lane="0" entrytime="00:13:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Timea" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" license="510414600003" swrid="5240601" athleteid="1956">
              <RESULTS>
                <RESULT eventid="1094" points="560" reactiontime="+81" swimtime="00:03:03.24" resultid="1957" heatid="4289" lane="4" entrytime="00:03:04.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:31.93" />
                    <SPLIT distance="150" swimtime="00:02:20.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="507" reactiontime="+90" swimtime="00:12:00.09" resultid="1958" heatid="4302" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                    <SPLIT distance="100" swimtime="00:01:24.86" />
                    <SPLIT distance="150" swimtime="00:02:10.35" />
                    <SPLIT distance="200" swimtime="00:02:56.14" />
                    <SPLIT distance="250" swimtime="00:03:41.73" />
                    <SPLIT distance="300" swimtime="00:04:27.66" />
                    <SPLIT distance="350" swimtime="00:05:13.38" />
                    <SPLIT distance="400" swimtime="00:05:59.63" />
                    <SPLIT distance="450" swimtime="00:06:44.49" />
                    <SPLIT distance="500" swimtime="00:07:29.52" />
                    <SPLIT distance="550" swimtime="00:08:15.11" />
                    <SPLIT distance="600" swimtime="00:09:01.19" />
                    <SPLIT distance="650" swimtime="00:09:46.77" />
                    <SPLIT distance="700" swimtime="00:10:32.38" />
                    <SPLIT distance="750" swimtime="00:11:17.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1233" points="699" reactiontime="+87" swimtime="00:03:12.61" resultid="1959" heatid="4328" lane="1" entrytime="00:03:18.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:34.23" />
                    <SPLIT distance="150" swimtime="00:02:24.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="447" reactiontime="+87" swimtime="00:01:19.00" resultid="1960" heatid="4339" lane="0" entrytime="00:01:18.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="646" reactiontime="+81" swimtime="00:01:27.32" resultid="1961" heatid="4365" lane="7" entrytime="00:01:29.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="496" reactiontime="+85" swimtime="00:02:48.21" resultid="1962" heatid="4395" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:02:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="672" reactiontime="+83" swimtime="00:00:39.03" resultid="1963" heatid="4441" lane="7" entrytime="00:00:39.14" entrycourse="LCM" />
                <RESULT eventid="1731" points="518" reactiontime="+88" swimtime="00:05:49.52" resultid="1964" heatid="4453" lane="4" entrytime="00:05:58.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                    <SPLIT distance="100" swimtime="00:01:23.23" />
                    <SPLIT distance="150" swimtime="00:02:08.08" />
                    <SPLIT distance="200" swimtime="00:02:53.27" />
                    <SPLIT distance="250" swimtime="00:03:36.78" />
                    <SPLIT distance="300" swimtime="00:04:21.45" />
                    <SPLIT distance="350" swimtime="00:05:06.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Ostapczuk" birthdate="1970-07-13" gender="M" nation="POL" athleteid="3706">
              <RESULTS>
                <RESULT eventid="1250" points="313" reactiontime="+101" swimtime="00:03:37.54" resultid="3707" heatid="4331" lane="4" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.85" />
                    <SPLIT distance="100" swimtime="00:01:42.25" />
                    <SPLIT distance="150" swimtime="00:02:39.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="287" reactiontime="+96" swimtime="00:01:22.13" resultid="3708" heatid="4345" lane="9" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="316" reactiontime="+93" swimtime="00:01:37.46" resultid="3709" heatid="4368" lane="6" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Mania" birthdate="1970-03-02" gender="M" nation="POL" swrid="5521445" athleteid="3718">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3719" heatid="4279" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="3720" heatid="4347" lane="8" entrytime="00:01:10.00" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="3721" heatid="4404" lane="8" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1386" points="278" reactiontime="+63" swimtime="00:02:49.87" resultid="1980" heatid="4491" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.22" />
                    <SPLIT distance="100" swimtime="00:01:33.31" />
                    <SPLIT distance="150" swimtime="00:02:16.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1965" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="1948" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="1972" number="3" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3706" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="1981" heatid="4495" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3706" number="1" />
                    <RELAYPOSITION athleteid="1965" number="2" />
                    <RELAYPOSITION athleteid="1972" number="3" />
                    <RELAYPOSITION athleteid="1948" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" points="325" reactiontime="+81" swimtime="00:02:28.81" resultid="1979" heatid="4489" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:15.75" />
                    <SPLIT distance="150" swimtime="00:01:55.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1956" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="1939" number="2" />
                    <RELAYPOSITION athleteid="1948" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3716" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1714" points="284" reactiontime="+84" swimtime="00:02:52.28" resultid="1982" heatid="4499" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.75" />
                    <SPLIT distance="100" swimtime="00:01:28.08" />
                    <SPLIT distance="150" swimtime="00:02:09.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1965" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="1956" number="2" />
                    <RELAYPOSITION athleteid="3706" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="1939" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="3087" name="Kauno Takas">
          <CONTACT email="kaunotakas@gmail.com" name="Romaldas Bickauskas" />
          <ATHLETES>
            <ATHLETE firstname="Vedestas" lastname="Sefleris" birthdate="1972-02-06" gender="M" nation="LTU" swrid="5186190" athleteid="3088">
              <RESULTS>
                <RESULT eventid="1112" points="710" reactiontime="+67" swimtime="00:02:27.04" resultid="3089" heatid="4296" lane="5" entrytime="00:02:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:08.36" />
                    <SPLIT distance="150" swimtime="00:01:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="777" reactiontime="+65" swimtime="00:00:58.89" resultid="3090" heatid="4351" lane="0" entrytime="00:00:58.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1525" points="767" reactiontime="+68" swimtime="00:02:09.58" resultid="3091" heatid="4407" lane="9" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:03.13" />
                    <SPLIT distance="150" swimtime="00:01:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="716" reactiontime="+65" swimtime="00:01:03.97" resultid="3092" heatid="4426" lane="5" entrytime="00:01:03.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1748" points="786" reactiontime="+80" swimtime="00:04:37.32" resultid="3093" heatid="4456" lane="8" entrytime="00:04:38.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="150" swimtime="00:01:40.14" />
                    <SPLIT distance="200" swimtime="00:02:16.03" />
                    <SPLIT distance="250" swimtime="00:02:52.07" />
                    <SPLIT distance="300" swimtime="00:03:28.24" />
                    <SPLIT distance="350" swimtime="00:04:03.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Linas" lastname="Kersevicius" birthdate="1971-06-18" gender="M" nation="LTU" swrid="4199514" athleteid="3094">
              <RESULTS>
                <RESULT eventid="1076" points="562" reactiontime="+83" swimtime="00:00:29.18" resultid="3095" heatid="4280" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1267" points="611" reactiontime="+82" swimtime="00:00:33.68" resultid="3096" heatid="4324" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1663" points="608" reactiontime="+85" swimtime="00:02:38.83" resultid="3097" heatid="4437" lane="0" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:18.42" />
                    <SPLIT distance="150" swimtime="00:01:59.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arlandas" lastname="Juodeska" birthdate="1961-12-26" gender="M" nation="LTU" swrid="4720137" athleteid="3098">
              <RESULTS>
                <RESULT eventid="1267" points="685" reactiontime="+72" swimtime="00:00:34.71" resultid="3099" heatid="4323" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1406" points="475" reactiontime="+81" swimtime="00:01:31.92" resultid="3100" heatid="4369" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="555" reactiontime="+72" swimtime="00:01:20.43" resultid="3101" heatid="4392" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="643" reactiontime="+76" swimtime="00:00:38.00" resultid="3102" heatid="4446" lane="1" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="2133" name="KS Warta Poznań">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Janyga" birthdate="1966-03-27" gender="M" nation="POL" license="100115700346" athleteid="4125">
              <RESULTS>
                <RESULT eventid="1076" points="616" reactiontime="+78" swimtime="00:00:28.73" resultid="4126" heatid="4283" lane="1" entrytime="00:00:27.89" />
                <RESULT eventid="1163" points="531" reactiontime="+86" swimtime="00:11:07.07" resultid="4127" heatid="4304" lane="3" entrytime="00:10:44.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                    <SPLIT distance="150" swimtime="00:01:55.63" />
                    <SPLIT distance="200" swimtime="00:02:36.82" />
                    <SPLIT distance="250" swimtime="00:03:18.85" />
                    <SPLIT distance="300" swimtime="00:04:00.83" />
                    <SPLIT distance="350" swimtime="00:04:42.59" />
                    <SPLIT distance="400" swimtime="00:05:24.45" />
                    <SPLIT distance="450" swimtime="00:06:06.84" />
                    <SPLIT distance="500" swimtime="00:06:50.27" />
                    <SPLIT distance="550" swimtime="00:07:33.54" />
                    <SPLIT distance="600" swimtime="00:08:16.97" />
                    <SPLIT distance="650" swimtime="00:08:59.74" />
                    <SPLIT distance="700" swimtime="00:09:42.84" />
                    <SPLIT distance="750" swimtime="00:10:25.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="607" reactiontime="+85" swimtime="00:00:34.28" resultid="4128" heatid="4324" lane="8" entrytime="00:00:33.16" />
                <RESULT eventid="1491" points="649" reactiontime="+74" swimtime="00:01:13.36" resultid="4129" heatid="4393" lane="5" entrytime="00:01:11.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="643" reactiontime="+91" swimtime="00:02:23.71" resultid="4130" heatid="4405" lane="8" entrytime="00:02:22.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:02:23.71" />
                    <SPLIT distance="150" swimtime="00:01:46.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="581" reactiontime="+83" swimtime="00:02:48.79" resultid="4131" heatid="4436" lane="9" entrytime="00:02:47.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:24.52" />
                    <SPLIT distance="150" swimtime="00:02:08.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Kuca" birthdate="1994-07-23" gender="M" nation="POL" license="100115700396" athleteid="4140">
              <RESULTS>
                <RESULT eventid="1076" points="782" reactiontime="+63" swimtime="00:00:24.20" resultid="4141" heatid="4286" lane="3" entrytime="00:00:24.49" />
                <RESULT eventid="1301" points="803" reactiontime="+78" swimtime="00:00:54.28" resultid="4142" heatid="4352" lane="6" entrytime="00:00:54.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="734" reactiontime="+62" swimtime="00:00:26.28" resultid="4143" heatid="4384" lane="6" entrytime="00:00:26.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Błażej" lastname="Wachowski" birthdate="1980-10-08" gender="M" nation="POL" license="100115700545" athleteid="4165">
              <RESULTS>
                <RESULT eventid="1076" points="516" reactiontime="+81" swimtime="00:00:28.98" resultid="4166" heatid="4283" lane="0" entrytime="00:00:27.90" />
                <RESULT eventid="1163" points="496" reactiontime="+84" swimtime="00:10:51.54" resultid="4167" heatid="4304" lane="5" entrytime="00:10:44.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:15.39" />
                    <SPLIT distance="150" swimtime="00:01:55.51" />
                    <SPLIT distance="200" swimtime="00:02:35.84" />
                    <SPLIT distance="250" swimtime="00:03:16.21" />
                    <SPLIT distance="300" swimtime="00:03:56.59" />
                    <SPLIT distance="350" swimtime="00:04:37.41" />
                    <SPLIT distance="400" swimtime="00:05:18.20" />
                    <SPLIT distance="450" swimtime="00:05:59.33" />
                    <SPLIT distance="500" swimtime="00:06:40.73" />
                    <SPLIT distance="550" swimtime="00:07:22.53" />
                    <SPLIT distance="600" swimtime="00:08:04.54" />
                    <SPLIT distance="650" swimtime="00:08:47.35" />
                    <SPLIT distance="700" swimtime="00:09:29.92" />
                    <SPLIT distance="750" swimtime="00:10:12.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="424" reactiontime="+87" swimtime="00:02:47.06" resultid="4168" heatid="4357" lane="8" entrytime="00:02:44.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:17.30" />
                    <SPLIT distance="150" swimtime="00:02:00.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="510" reactiontime="+90" swimtime="00:02:22.28" resultid="4169" heatid="4405" lane="0" entrytime="00:02:22.20">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="464" reactiontime="+86" swimtime="00:01:12.58" resultid="4170" heatid="4425" lane="1" entrytime="00:01:12.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="513" reactiontime="+94" swimtime="00:05:08.26" resultid="4171" heatid="4458" lane="8" entrytime="00:05:12.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="150" swimtime="00:01:53.82" />
                    <SPLIT distance="200" swimtime="00:02:33.49" />
                    <SPLIT distance="250" swimtime="00:03:13.00" />
                    <SPLIT distance="300" swimtime="00:03:52.41" />
                    <SPLIT distance="350" swimtime="00:04:32.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kotecka" birthdate="1965-05-08" gender="F" nation="POL" license="100115600357" athleteid="4132">
              <RESULTS>
                <RESULT eventid="1146" points="371" swimtime="00:13:33.81" resultid="4133" heatid="4300" lane="8" entrytime="00:13:25.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                    <SPLIT distance="100" swimtime="00:01:32.08" />
                    <SPLIT distance="150" swimtime="00:02:23.08" />
                    <SPLIT distance="200" swimtime="00:03:13.61" />
                    <SPLIT distance="250" swimtime="00:04:04.74" />
                    <SPLIT distance="300" swimtime="00:04:55.85" />
                    <SPLIT distance="350" swimtime="00:05:47.86" />
                    <SPLIT distance="400" swimtime="00:06:39.69" />
                    <SPLIT distance="450" swimtime="00:07:31.09" />
                    <SPLIT distance="500" swimtime="00:08:22.58" />
                    <SPLIT distance="550" swimtime="00:09:14.11" />
                    <SPLIT distance="600" swimtime="00:10:06.29" />
                    <SPLIT distance="650" swimtime="00:10:58.30" />
                    <SPLIT distance="700" swimtime="00:11:50.83" />
                    <SPLIT distance="750" swimtime="00:12:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="264" reactiontime="+118" swimtime="00:00:49.87" resultid="4134" heatid="4314" lane="6" entrytime="00:00:49.37" />
                <RESULT eventid="1284" points="351" reactiontime="+103" swimtime="00:01:27.91" resultid="4135" heatid="4337" lane="4" entrytime="00:01:29.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="300" reactiontime="+113" swimtime="00:01:44.15" resultid="4136" heatid="4388" lane="5" entrytime="00:01:11.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="379" reactiontime="+99" swimtime="00:03:08.33" resultid="4137" heatid="4397" lane="0" entrytime="00:03:09.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="317" reactiontime="+134" swimtime="00:03:42.67" resultid="4138" heatid="4430" lane="6" entrytime="00:03:38.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.30" />
                    <SPLIT distance="100" swimtime="00:01:49.59" />
                    <SPLIT distance="150" swimtime="00:02:47.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="356" reactiontime="+103" swimtime="00:06:40.03" resultid="4139" heatid="4453" lane="7" entrytime="00:06:39.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                    <SPLIT distance="100" swimtime="00:01:32.97" />
                    <SPLIT distance="150" swimtime="00:02:23.63" />
                    <SPLIT distance="200" swimtime="00:03:14.01" />
                    <SPLIT distance="250" swimtime="00:04:05.51" />
                    <SPLIT distance="300" swimtime="00:04:57.07" />
                    <SPLIT distance="350" swimtime="00:05:49.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Osik" birthdate="1976-01-02" gender="M" nation="POL" license="500115700521" athleteid="4150">
              <RESULTS>
                <RESULT eventid="1076" points="562" reactiontime="+81" swimtime="00:00:28.53" resultid="4151" heatid="4283" lane="8" entrytime="00:00:27.89" />
                <RESULT eventid="1197" points="623" reactiontime="+87" swimtime="00:19:29.76" resultid="4152" heatid="4309" lane="7" entrytime="00:19:28.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="150" swimtime="00:01:52.60" />
                    <SPLIT distance="250" swimtime="00:03:10.55" />
                    <SPLIT distance="350" swimtime="00:04:29.83" />
                    <SPLIT distance="400" swimtime="00:06:28.99" />
                    <SPLIT distance="450" swimtime="00:05:49.18" />
                    <SPLIT distance="500" swimtime="00:07:48.21" />
                    <SPLIT distance="550" swimtime="00:07:08.31" />
                    <SPLIT distance="600" swimtime="00:09:07.55" />
                    <SPLIT distance="650" swimtime="00:08:27.39" />
                    <SPLIT distance="700" swimtime="00:10:25.13" />
                    <SPLIT distance="750" swimtime="00:09:45.93" />
                    <SPLIT distance="800" swimtime="00:11:44.03" />
                    <SPLIT distance="850" swimtime="00:11:04.64" />
                    <SPLIT distance="900" swimtime="00:13:01.99" />
                    <SPLIT distance="950" swimtime="00:12:22.66" />
                    <SPLIT distance="1000" swimtime="00:14:19.14" />
                    <SPLIT distance="1050" swimtime="00:13:40.44" />
                    <SPLIT distance="1100" swimtime="00:15:37.65" />
                    <SPLIT distance="1150" swimtime="00:14:58.45" />
                    <SPLIT distance="1200" swimtime="00:18:13.96" />
                    <SPLIT distance="1250" swimtime="00:16:17.18" />
                    <SPLIT distance="1350" swimtime="00:17:35.00" />
                    <SPLIT distance="1450" swimtime="00:18:51.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="555" reactiontime="+71" swimtime="00:00:33.60" resultid="4153" heatid="4324" lane="6" entrytime="00:00:32.10" />
                <RESULT eventid="1491" points="610" reactiontime="+82" swimtime="00:01:10.89" resultid="4154" heatid="4393" lane="6" entrytime="00:01:14.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="647" reactiontime="+85" swimtime="00:02:16.15" resultid="4155" heatid="4405" lane="4" entrytime="00:02:17.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="100" swimtime="00:01:06.05" />
                    <SPLIT distance="150" swimtime="00:01:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="628" reactiontime="+82" swimtime="00:02:33.62" resultid="4156" heatid="4436" lane="1" entrytime="00:02:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:15.05" />
                    <SPLIT distance="150" swimtime="00:01:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="641" reactiontime="+88" swimtime="00:04:51.20" resultid="4157" heatid="4457" lane="2" entrytime="00:04:49.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:09.22" />
                    <SPLIT distance="150" swimtime="00:01:46.13" />
                    <SPLIT distance="200" swimtime="00:02:23.94" />
                    <SPLIT distance="250" swimtime="00:03:00.23" />
                    <SPLIT distance="300" swimtime="00:03:37.25" />
                    <SPLIT distance="350" swimtime="00:04:14.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Majchrzak" birthdate="1983-01-21" gender="M" nation="POL" license="104215700019" athleteid="4144">
              <RESULTS>
                <RESULT eventid="1076" points="530" reactiontime="+75" swimtime="00:00:28.13" resultid="4145" heatid="4283" lane="6" entrytime="00:00:27.50" />
                <RESULT eventid="1301" points="539" reactiontime="+77" swimtime="00:01:02.40" resultid="4146" heatid="4350" lane="1" entrytime="00:00:59.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="556" reactiontime="+77" swimtime="00:00:29.36" resultid="4147" heatid="4382" lane="4" entrytime="00:00:29.12" />
                <RESULT eventid="1525" points="525" reactiontime="+84" swimtime="00:02:19.86" resultid="4148" heatid="4406" lane="7" entrytime="00:02:13.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:44.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="493" reactiontime="+82" swimtime="00:01:07.93" resultid="4149" heatid="4426" lane="1" entrytime="00:01:06.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szymkowiak" birthdate="1980-04-12" gender="M" nation="POL" license="500115700523" athleteid="4158">
              <RESULTS>
                <RESULT eventid="1076" points="654" reactiontime="+67" swimtime="00:00:26.79" resultid="4159" heatid="4285" lane="6" entrytime="00:00:26.32" />
                <RESULT eventid="1112" points="598" reactiontime="+75" swimtime="00:02:35.02" resultid="4160" heatid="4297" lane="0" entrytime="00:02:27.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:01:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1250" points="677" reactiontime="+74" swimtime="00:02:37.85" resultid="4161" heatid="4334" lane="7" entrytime="00:02:39.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:15.08" />
                    <SPLIT distance="150" swimtime="00:01:56.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="799" reactiontime="+72" swimtime="00:01:08.55" resultid="4162" heatid="4371" lane="6" entrytime="00:01:07.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="4163" heatid="4415" lane="3" entrytime="00:05:47.00" />
                <RESULT eventid="1697" points="829" reactiontime="+69" swimtime="00:00:30.70" resultid="4164" heatid="4449" lane="6" entrytime="00:00:30.42" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Wieja" birthdate="1978-09-08" gender="M" nation="POL" license="500115700467" swrid="5331775" athleteid="4172">
              <RESULTS>
                <RESULT eventid="1076" points="665" reactiontime="+68" swimtime="00:00:26.64" resultid="4173" heatid="4284" lane="8" entrytime="00:00:27.08" />
                <RESULT eventid="1112" points="660" reactiontime="+71" swimtime="00:02:30.01" resultid="4174" heatid="4296" lane="2" entrytime="00:02:31.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:56.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="603" reactiontime="+78" swimtime="00:00:32.11" resultid="4175" heatid="4325" lane="9" entrytime="00:00:31.61" />
                <RESULT eventid="1301" points="670" reactiontime="+73" swimtime="00:00:58.53" resultid="4176" heatid="4350" lane="7" entrytime="00:00:59.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="541" reactiontime="+69" swimtime="00:01:11.74" resultid="4177" heatid="4394" lane="9" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="4178" heatid="4415" lane="5" entrytime="00:05:45.12" />
                <RESULT comment="G1" eventid="1663" points="544" reactiontime="+75" swimtime="00:02:36.92" resultid="4179" heatid="4437" lane="1" entrytime="00:02:35.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:01:16.37" />
                    <SPLIT distance="150" swimtime="00:01:57.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="541" reactiontime="+66" swimtime="00:00:35.39" resultid="4180" heatid="4447" lane="0" entrytime="00:00:36.41" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Witt" birthdate="1991-08-11" gender="M" nation="POL" license="500115700645" swrid="5062813" athleteid="4181">
              <RESULTS>
                <RESULT eventid="1076" points="689" reactiontime="+70" swimtime="00:00:25.05" resultid="4182" heatid="4286" lane="5" entrytime="00:00:24.34" />
                <RESULT eventid="1267" points="568" reactiontime="+80" swimtime="00:00:31.36" resultid="4183" heatid="4325" lane="3" entrytime="00:00:29.90" />
                <RESULT eventid="1301" points="694" reactiontime="+74" swimtime="00:00:56.26" resultid="4184" heatid="4351" lane="3" entrytime="00:00:56.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="597" reactiontime="+76" swimtime="00:00:27.62" resultid="4185" heatid="4384" lane="9" entrytime="00:00:27.97" />
                <RESULT eventid="1525" points="597" reactiontime="+75" swimtime="00:02:10.13" resultid="4186" heatid="4407" lane="0" entrytime="00:02:08.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.40" />
                    <SPLIT distance="150" swimtime="00:01:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="569" reactiontime="+74" swimtime="00:01:04.75" resultid="4187" heatid="4426" lane="7" entrytime="00:01:06.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="570" reactiontime="+77" swimtime="00:04:47.23" resultid="4188" heatid="4457" lane="6" entrytime="00:04:49.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="150" swimtime="00:01:46.08" />
                    <SPLIT distance="200" swimtime="00:02:23.27" />
                    <SPLIT distance="250" swimtime="00:03:00.43" />
                    <SPLIT distance="300" swimtime="00:03:37.12" />
                    <SPLIT distance="350" swimtime="00:04:13.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1386" points="750" reactiontime="+61" swimtime="00:01:56.07" resultid="4189" heatid="4493" lane="5" entrytime="00:01:57.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:01.83" />
                    <SPLIT distance="150" swimtime="00:01:27.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4172" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4158" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4140" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="4125" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1386" points="504" reactiontime="+80" swimtime="00:02:08.53" resultid="4190" heatid="4493" lane="2" entrytime="00:02:03.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:40.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4181" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4144" number="2" />
                    <RELAYPOSITION athleteid="4150" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="4165" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1559" points="709" reactiontime="+68" swimtime="00:01:46.45" resultid="4191" heatid="4497" lane="5" entrytime="00:01:44.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                    <SPLIT distance="100" swimtime="00:00:52.87" />
                    <SPLIT distance="150" swimtime="00:01:21.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4172" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4158" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="4125" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4181" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Marcin" gender="M" lastname="Szymkowiak" license="500115700523" type="HEADCOACH" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3678" name="Rydułtowska Akademia Aktywnego Seniora 60+">
          <ATHLETES>
            <ATHLETE firstname="MARIA" lastname="LIPPA" birthdate="1946-01-01" gender="F" nation="POL" swrid="5484413" athleteid="3688">
              <RESULTS>
                <RESULT eventid="1059" points="42" swimtime="00:01:38.39" resultid="3689" heatid="4268" lane="2" entrytime="00:01:32.99" entrycourse="SCM" />
                <RESULT eventid="1215" points="67" reactiontime="+167" swimtime="00:01:38.54" resultid="3690" heatid="4313" lane="3" entrytime="00:01:38.15" entrycourse="SCM" />
                <RESULT eventid="1284" points="64" swimtime="00:03:13.12" resultid="3691" heatid="4337" lane="0" entrytime="00:03:09.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="71" reactiontime="+173" swimtime="00:03:34.52" resultid="3692" heatid="4387" lane="9" entrytime="00:03:26.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="84" swimtime="00:06:38.43" resultid="3693" heatid="4395" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:32.45" />
                    <SPLIT distance="100" swimtime="00:03:13.81" />
                    <SPLIT distance="150" swimtime="00:04:56.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="97" swimtime="00:13:30.64" resultid="3694" heatid="4455" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.72" />
                    <SPLIT distance="100" swimtime="00:03:08.86" />
                    <SPLIT distance="150" swimtime="00:04:52.91" />
                    <SPLIT distance="200" swimtime="00:06:34.53" />
                    <SPLIT distance="250" swimtime="00:08:19.55" />
                    <SPLIT distance="300" swimtime="00:10:07.74" />
                    <SPLIT distance="350" swimtime="00:11:49.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="197" reactiontime="+194" swimtime="00:05:38.34" resultid="3695" heatid="4428" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.94" />
                    <SPLIT distance="100" swimtime="00:03:41.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="CIECIOR" birthdate="1953-01-01" gender="M" nation="POL" swrid="4934027" athleteid="3679">
              <RESULTS>
                <RESULT eventid="1112" points="295" reactiontime="+91" swimtime="00:03:38.06" resultid="3680" heatid="4293" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                    <SPLIT distance="100" swimtime="00:01:43.31" />
                    <SPLIT distance="150" swimtime="00:02:49.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1197" points="369" reactiontime="+89" swimtime="00:27:16.09" resultid="3681" heatid="4310" lane="1" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                    <SPLIT distance="100" swimtime="00:01:38.26" />
                    <SPLIT distance="150" swimtime="00:02:32.42" />
                    <SPLIT distance="200" swimtime="00:03:27.05" />
                    <SPLIT distance="250" swimtime="00:04:21.73" />
                    <SPLIT distance="300" swimtime="00:05:16.57" />
                    <SPLIT distance="350" swimtime="00:06:11.69" />
                    <SPLIT distance="400" swimtime="00:07:06.62" />
                    <SPLIT distance="450" swimtime="00:08:01.92" />
                    <SPLIT distance="500" swimtime="00:08:56.97" />
                    <SPLIT distance="550" swimtime="00:09:52.15" />
                    <SPLIT distance="600" swimtime="00:10:47.47" />
                    <SPLIT distance="650" swimtime="00:11:42.47" />
                    <SPLIT distance="700" swimtime="00:12:36.39" />
                    <SPLIT distance="750" swimtime="00:13:31.58" />
                    <SPLIT distance="800" swimtime="00:14:26.81" />
                    <SPLIT distance="850" swimtime="00:15:21.97" />
                    <SPLIT distance="900" swimtime="00:16:16.23" />
                    <SPLIT distance="950" swimtime="00:17:11.30" />
                    <SPLIT distance="1000" swimtime="00:18:06.28" />
                    <SPLIT distance="1050" swimtime="00:19:01.38" />
                    <SPLIT distance="1100" swimtime="00:19:56.71" />
                    <SPLIT distance="1150" swimtime="00:20:52.03" />
                    <SPLIT distance="1200" swimtime="00:21:46.78" />
                    <SPLIT distance="1250" swimtime="00:22:41.91" />
                    <SPLIT distance="1300" swimtime="00:23:37.52" />
                    <SPLIT distance="1350" swimtime="00:24:33.23" />
                    <SPLIT distance="1400" swimtime="00:25:28.62" />
                    <SPLIT distance="1450" swimtime="00:26:23.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="226" reactiontime="+82" swimtime="00:04:11.86" resultid="3682" heatid="4355" lane="6" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.31" />
                    <SPLIT distance="100" swimtime="00:02:01.21" />
                    <SPLIT distance="150" swimtime="00:03:06.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="376" reactiontime="+93" swimtime="00:00:42.90" resultid="3683" heatid="4322" lane="0" entrytime="00:00:40.65" entrycourse="SCM" />
                <RESULT eventid="1457" points="340" reactiontime="+85" swimtime="00:00:40.65" resultid="3684" heatid="4379" lane="6" entrytime="00:00:41.21" entrycourse="SCM" />
                <RESULT eventid="1593" points="265" reactiontime="+92" swimtime="00:08:07.77" resultid="3685" heatid="4416" lane="7" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.62" />
                    <SPLIT distance="100" swimtime="00:02:00.95" />
                    <SPLIT distance="150" swimtime="00:03:03.29" />
                    <SPLIT distance="200" swimtime="00:04:05.26" />
                    <SPLIT distance="250" swimtime="00:05:14.10" />
                    <SPLIT distance="300" swimtime="00:06:22.60" />
                    <SPLIT distance="350" swimtime="00:07:15.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="222" reactiontime="+87" swimtime="00:01:48.65" resultid="3686" heatid="4423" lane="6" entrytime="00:01:49.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="325" reactiontime="+104" swimtime="00:03:48.53" resultid="3687" heatid="4434" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.17" />
                    <SPLIT distance="100" swimtime="00:01:49.00" />
                    <SPLIT distance="150" swimtime="00:02:49.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="WŁADYSŁAW" lastname="SZUREK" birthdate="1940-01-01" gender="M" nation="POL" swrid="5450542" athleteid="3696">
              <RESULTS>
                <RESULT eventid="1076" points="46" swimtime="00:01:29.52" resultid="3697" heatid="4275" lane="6" entrytime="00:01:17.05" entrycourse="SCM" />
                <RESULT eventid="1267" points="34" reactiontime="+115" swimtime="00:01:57.95" resultid="3698" heatid="4319" lane="4" entrytime="00:01:38.29" entrycourse="SCM" />
                <RESULT eventid="1301" points="50" swimtime="00:03:15.00" resultid="3699" heatid="4343" lane="5" entrytime="00:02:45.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="31" reactiontime="+105" swimtime="00:04:34.26" resultid="3700" heatid="4390" lane="9" entrytime="00:03:34.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:04.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="46" swimtime="00:07:27.78" resultid="3701" heatid="4400" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.04" />
                    <SPLIT distance="100" swimtime="00:03:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="36" reactiontime="+103" swimtime="00:09:50.44" resultid="3702" heatid="4432" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:03.91" />
                    <SPLIT distance="150" swimtime="00:07:10.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="113/14" nation="POL" clubid="3258" name="Fundacja HASTEN">
          <CONTACT email="hasten@hasten.pl" name="Bochyńska Sonia" />
          <ATHLETES>
            <ATHLETE firstname="Natalia" lastname="Pawlaczek" birthdate="1993-04-01" gender="F" nation="POL" athleteid="3259">
              <RESULTS>
                <RESULT eventid="1059" points="804" reactiontime="+77" swimtime="00:00:27.34" resultid="3260" heatid="4272" lane="3" entrytime="00:00:27.50" />
                <RESULT eventid="1284" points="842" reactiontime="+78" swimtime="00:01:00.31" resultid="3261" heatid="4340" lane="4" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="704" reactiontime="+76" swimtime="00:00:29.59" resultid="3262" heatid="4375" lane="5" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Węgier" birthdate="1996-02-01" gender="F" nation="POL" swrid="4228268" athleteid="3271">
              <RESULTS>
                <RESULT eventid="1215" points="496" reactiontime="+73" swimtime="00:00:35.86" resultid="3272" heatid="4316" lane="9" entrytime="00:00:36.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Karpińska" birthdate="1991-07-26" gender="F" nation="POL" athleteid="3267">
              <RESULTS>
                <RESULT eventid="1059" points="677" reactiontime="+71" swimtime="00:00:29.31" resultid="3268" heatid="4272" lane="9" entrytime="00:00:29.99" />
                <RESULT eventid="1284" points="623" reactiontime="+80" swimtime="00:01:04.69" resultid="3269" heatid="4340" lane="2" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="661" reactiontime="+82" swimtime="00:00:31.54" resultid="3270" heatid="4375" lane="8" entrytime="00:00:31.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sonia" lastname="Bochyńska" birthdate="1990-06-10" gender="F" nation="POL" swrid="4061587" athleteid="3263">
              <RESULTS>
                <RESULT eventid="1059" points="587" reactiontime="+78" swimtime="00:00:30.74" resultid="3264" heatid="4272" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1215" points="616" reactiontime="+70" swimtime="00:00:33.58" resultid="3265" heatid="4316" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1440" points="667" reactiontime="+74" swimtime="00:00:31.45" resultid="3266" heatid="4375" lane="7" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1369" points="701" reactiontime="+68" swimtime="00:02:15.16" resultid="3273" heatid="4490" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="150" swimtime="00:01:45.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3271" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3259" number="2" />
                    <RELAYPOSITION athleteid="3267" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3263" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1542" points="819" reactiontime="+78" swimtime="00:01:57.89" resultid="3274" heatid="4494" lane="4" entrytime="00:01:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="100" swimtime="00:00:59.00" />
                    <SPLIT distance="150" swimtime="00:01:30.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3267" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3263" number="2" />
                    <RELAYPOSITION athleteid="3271" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3259" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" clubid="2687" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501370222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Ślężyński" birthdate="1931-04-27" gender="M" nation="POL" license="100611700315" swrid="4992723" athleteid="2688">
              <RESULTS>
                <RESULT eventid="1076" points="236" reactiontime="+115" swimtime="00:01:05.92" resultid="2689" heatid="4275" lane="2" entrytime="00:01:25.66" />
                <RESULT eventid="1250" points="260" reactiontime="+100" swimtime="00:07:20.64" resultid="2691" heatid="4330" lane="3" entrytime="00:07:45.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:43.95" />
                    <SPLIT distance="100" swimtime="00:03:38.08" />
                    <SPLIT distance="150" swimtime="00:05:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="98" reactiontime="+90" swimtime="00:03:32.03" resultid="2692" heatid="4343" lane="3" entrytime="00:03:15.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="204" reactiontime="+86" swimtime="00:03:32.65" resultid="2693" heatid="4367" lane="8" entrytime="00:03:35.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:41.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="153" swimtime="00:06:39.54" resultid="2694" heatid="4401" lane="7" entrytime="00:06:36.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.00" />
                    <SPLIT distance="150" swimtime="00:05:07.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="162" reactiontime="+98" swimtime="00:01:32.95" resultid="2695" heatid="4443" lane="6" entrytime="00:01:45.57" />
                <RESULT eventid="1748" points="165" reactiontime="+113" swimtime="00:13:57.32" resultid="2696" heatid="4462" lane="3" entrytime="00:15:05.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.16" />
                    <SPLIT distance="100" swimtime="00:03:24.91" />
                    <SPLIT distance="150" swimtime="00:05:14.85" />
                    <SPLIT distance="200" swimtime="00:07:04.06" />
                    <SPLIT distance="250" swimtime="00:08:53.20" />
                    <SPLIT distance="300" swimtime="00:10:38.46" />
                    <SPLIT distance="350" swimtime="00:12:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="89" swimtime="00:34:18.14" resultid="2697" heatid="4306" lane="8" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:43.56" />
                    <SPLIT distance="100" swimtime="00:03:58.93" />
                    <SPLIT distance="150" swimtime="00:06:04.90" />
                    <SPLIT distance="200" swimtime="00:08:14.89" />
                    <SPLIT distance="250" swimtime="00:10:22.91" />
                    <SPLIT distance="300" swimtime="00:12:36.84" />
                    <SPLIT distance="350" swimtime="00:14:53.39" />
                    <SPLIT distance="400" swimtime="00:17:08.57" />
                    <SPLIT distance="450" swimtime="00:19:20.34" />
                    <SPLIT distance="500" swimtime="00:21:32.30" />
                    <SPLIT distance="550" swimtime="00:23:50.56" />
                    <SPLIT distance="600" swimtime="00:26:08.66" />
                    <SPLIT distance="650" swimtime="00:28:34.54" />
                    <SPLIT distance="700" swimtime="00:30:44.01" />
                    <SPLIT distance="750" swimtime="00:32:42.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2810" name="MASTERS Zdzieszowice">
          <CONTACT email="masters.zdzieszowice@gmail.com" name="jajuga" phone="505127695" />
          <ATHLETES>
            <ATHLETE firstname="Dorota" lastname="Woźniak" birthdate="1973-09-18" gender="F" nation="POL" swrid="4992846" athleteid="2811">
              <RESULTS>
                <RESULT eventid="1215" points="438" reactiontime="+78" swimtime="00:00:40.85" resultid="2812" heatid="4315" lane="6" entrytime="00:00:38.11" />
                <RESULT eventid="1335" points="367" reactiontime="+102" swimtime="00:03:21.62" resultid="2813" heatid="4354" lane="2" entrytime="00:03:00.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                    <SPLIT distance="150" swimtime="00:02:27.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="425" reactiontime="+97" swimtime="00:00:37.78" resultid="2814" heatid="4374" lane="6" entrytime="00:00:37.34" />
                <RESULT eventid="1576" points="454" reactiontime="+96" swimtime="00:06:48.35" resultid="2815" heatid="4412" lane="2" entrytime="00:06:34.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:31.70" />
                    <SPLIT distance="150" swimtime="00:02:25.07" />
                    <SPLIT distance="200" swimtime="00:03:16.53" />
                    <SPLIT distance="250" swimtime="00:04:13.93" />
                    <SPLIT distance="300" swimtime="00:05:13.64" />
                    <SPLIT distance="350" swimtime="00:06:01.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="425" reactiontime="+90" swimtime="00:01:26.43" resultid="2816" heatid="4420" lane="4" entrytime="00:01:23.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="424" reactiontime="+83" swimtime="00:03:11.75" resultid="2817" heatid="4431" lane="2" entrytime="00:03:00.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                    <SPLIT distance="100" swimtime="00:01:33.68" />
                    <SPLIT distance="150" swimtime="00:02:23.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04514" nation="POL" clubid="3148" name="UKS 307 Warszawa-Mokotów">
          <CONTACT email="uks307warszawa@gmail.com" name="Ilczyszyn" />
          <ATHLETES>
            <ATHLETE firstname="Damian" lastname="Ziółkowski" birthdate="1978-02-03" gender="M" nation="POL" license="104514700202" athleteid="3149">
              <RESULTS>
                <RESULT eventid="1457" points="439" reactiontime="+80" swimtime="00:00:32.98" resultid="3150" heatid="4380" lane="3" entrytime="00:00:34.17" />
                <RESULT eventid="1629" points="257" reactiontime="+79" swimtime="00:01:28.34" resultid="3151" heatid="4424" lane="1" entrytime="00:01:30.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3356" name="Masters Białystok">
          <CONTACT city="Białystok" email="ajeje@poczta.onet.pl" name="Twarowski Andrzej" phone="+48600361168" state="PODLA" street="Pułaskiego 133/6" zip="15-337" />
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Twarowski" birthdate="1965-05-24" gender="M" nation="POL" athleteid="3357">
              <RESULTS>
                <RESULT eventid="1197" points="286" reactiontime="+98" swimtime="00:26:21.93" resultid="3358" heatid="4310" lane="2" entrytime="00:26:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.63" />
                    <SPLIT distance="100" swimtime="00:01:36.21" />
                    <SPLIT distance="150" swimtime="00:02:29.53" />
                    <SPLIT distance="200" swimtime="00:03:21.73" />
                    <SPLIT distance="250" swimtime="00:04:15.79" />
                    <SPLIT distance="300" swimtime="00:05:08.01" />
                    <SPLIT distance="350" swimtime="00:06:02.39" />
                    <SPLIT distance="400" swimtime="00:06:55.19" />
                    <SPLIT distance="450" swimtime="00:07:49.47" />
                    <SPLIT distance="500" swimtime="00:08:41.62" />
                    <SPLIT distance="550" swimtime="00:09:33.71" />
                    <SPLIT distance="600" swimtime="00:10:26.66" />
                    <SPLIT distance="650" swimtime="00:11:19.64" />
                    <SPLIT distance="700" swimtime="00:12:12.63" />
                    <SPLIT distance="750" swimtime="00:13:06.19" />
                    <SPLIT distance="800" swimtime="00:13:59.49" />
                    <SPLIT distance="850" swimtime="00:14:52.45" />
                    <SPLIT distance="900" swimtime="00:15:46.40" />
                    <SPLIT distance="950" swimtime="00:16:39.12" />
                    <SPLIT distance="1000" swimtime="00:17:32.41" />
                    <SPLIT distance="1050" swimtime="00:18:26.03" />
                    <SPLIT distance="1100" swimtime="00:19:20.44" />
                    <SPLIT distance="1150" swimtime="00:20:13.23" />
                    <SPLIT distance="1200" swimtime="00:21:06.72" />
                    <SPLIT distance="1250" swimtime="00:22:00.33" />
                    <SPLIT distance="1300" swimtime="00:22:54.23" />
                    <SPLIT distance="1350" swimtime="00:23:47.19" />
                    <SPLIT distance="1400" swimtime="00:24:40.06" />
                    <SPLIT distance="1450" swimtime="00:25:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="426" reactiontime="+77" swimtime="00:00:38.57" resultid="3359" heatid="4322" lane="2" entrytime="00:00:39.00" entrycourse="LCM" />
                <RESULT eventid="1352" points="179" reactiontime="+98" swimtime="00:04:02.58" resultid="3360" heatid="4355" lane="4" entrytime="00:03:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.69" />
                    <SPLIT distance="100" swimtime="00:01:54.51" />
                    <SPLIT distance="150" swimtime="00:03:00.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="354" reactiontime="+73" swimtime="00:01:29.80" resultid="3361" heatid="4391" lane="4" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="268" reactiontime="+101" swimtime="00:07:47.95" resultid="3362" heatid="4416" lane="8" entrytime="00:07:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.56" />
                    <SPLIT distance="100" swimtime="00:01:57.24" />
                    <SPLIT distance="150" swimtime="00:02:56.96" />
                    <SPLIT distance="200" swimtime="00:03:57.51" />
                    <SPLIT distance="250" swimtime="00:05:01.06" />
                    <SPLIT distance="300" swimtime="00:06:04.07" />
                    <SPLIT distance="350" swimtime="00:06:58.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="310" reactiontime="+70" swimtime="00:03:28.17" resultid="3363" heatid="4434" lane="4" entrytime="00:03:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="100" swimtime="00:01:43.98" />
                    <SPLIT distance="150" swimtime="00:02:37.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="3364" heatid="4461" lane="4" entrytime="00:06:40.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01713" nation="POL" region="13" clubid="1807" name="Stowarzyszenie Pływackie Masters Olsztyn">
          <CONTACT name="Goździejewska" />
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Koźlikowski" birthdate="1961-09-09" gender="M" nation="POL" license="501713700011" swrid="4992727" athleteid="1885">
              <RESULTS>
                <RESULT eventid="1112" points="432" reactiontime="+99" swimtime="00:03:07.78" resultid="1886" heatid="4291" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="100" swimtime="00:01:33.77" />
                    <SPLIT distance="150" swimtime="00:02:25.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="449" reactiontime="+102" swimtime="00:12:24.09" resultid="1887" heatid="4307" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:26.47" />
                    <SPLIT distance="150" swimtime="00:02:13.41" />
                    <SPLIT distance="200" swimtime="00:03:00.67" />
                    <SPLIT distance="250" swimtime="00:03:48.44" />
                    <SPLIT distance="300" swimtime="00:04:36.34" />
                    <SPLIT distance="350" swimtime="00:05:24.21" />
                    <SPLIT distance="400" swimtime="00:06:12.48" />
                    <SPLIT distance="450" swimtime="00:06:59.87" />
                    <SPLIT distance="500" swimtime="00:07:47.51" />
                    <SPLIT distance="550" swimtime="00:08:34.50" />
                    <SPLIT distance="600" swimtime="00:09:21.41" />
                    <SPLIT distance="650" swimtime="00:10:08.12" />
                    <SPLIT distance="700" swimtime="00:10:54.90" />
                    <SPLIT distance="750" swimtime="00:11:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="488" reactiontime="+103" swimtime="00:03:23.47" resultid="1888" heatid="4329" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                    <SPLIT distance="100" swimtime="00:01:35.84" />
                    <SPLIT distance="150" swimtime="00:02:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="416" reactiontime="+105" swimtime="00:06:52.91" resultid="1889" heatid="4416" lane="3" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                    <SPLIT distance="100" swimtime="00:01:41.04" />
                    <SPLIT distance="150" swimtime="00:02:38.88" />
                    <SPLIT distance="200" swimtime="00:03:36.22" />
                    <SPLIT distance="250" swimtime="00:04:29.57" />
                    <SPLIT distance="300" swimtime="00:05:23.84" />
                    <SPLIT distance="350" swimtime="00:06:08.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="464" reactiontime="+101" swimtime="00:05:57.71" resultid="1890" heatid="4462" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                    <SPLIT distance="100" swimtime="00:01:23.93" />
                    <SPLIT distance="150" swimtime="00:02:08.86" />
                    <SPLIT distance="200" swimtime="00:02:54.54" />
                    <SPLIT distance="250" swimtime="00:03:40.53" />
                    <SPLIT distance="300" swimtime="00:04:26.61" />
                    <SPLIT distance="350" swimtime="00:05:12.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="4239" heatid="4403" lane="0" entrytime="00:02:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Mówiński" birthdate="1969-09-01" gender="M" nation="POL" license="501713700007" swrid="4992726" athleteid="1913">
              <RESULTS>
                <RESULT eventid="1352" points="336" reactiontime="+91" swimtime="00:03:11.82" resultid="1914" heatid="4355" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                    <SPLIT distance="100" swimtime="00:01:29.96" />
                    <SPLIT distance="150" swimtime="00:02:21.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="395" reactiontime="+85" swimtime="00:02:41.73" resultid="1915" heatid="4400" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                    <SPLIT distance="150" swimtime="00:02:00.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="410" reactiontime="+96" swimtime="00:05:44.37" resultid="1916" heatid="4462" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                    <SPLIT distance="150" swimtime="00:02:05.00" />
                    <SPLIT distance="200" swimtime="00:02:49.67" />
                    <SPLIT distance="250" swimtime="00:03:33.92" />
                    <SPLIT distance="300" swimtime="00:04:18.18" />
                    <SPLIT distance="350" swimtime="00:05:02.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Grabowski" birthdate="1989-02-10" gender="M" nation="POL" swrid="5230712" athleteid="2771">
              <RESULTS>
                <RESULT eventid="1076" points="552" reactiontime="+76" swimtime="00:00:26.98" resultid="2772" heatid="4285" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="1301" points="500" reactiontime="+81" swimtime="00:01:02.75" resultid="2773" heatid="4350" lane="9" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="420" reactiontime="+75" swimtime="00:00:31.07" resultid="2774" heatid="4382" lane="2" entrytime="00:00:29.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kozikowski" birthdate="1980-03-13" gender="M" nation="POL" license="501713700027" swrid="4992728" athleteid="1878">
              <RESULTS>
                <RESULT eventid="1112" status="DNS" swimtime="00:00:00.00" resultid="1879" heatid="4291" lane="7" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="1880" heatid="4307" lane="4" />
                <RESULT eventid="1250" status="DNS" swimtime="00:00:00.00" resultid="1881" heatid="4334" lane="1" entrytime="00:02:40.37" entrycourse="SCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="1882" heatid="4371" lane="8" entrytime="00:01:13.06" entrycourse="SCM" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="1883" heatid="4400" lane="3" />
                <RESULT eventid="1697" status="DNS" swimtime="00:00:00.00" resultid="1884" heatid="4448" lane="4" entrytime="00:00:33.19" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oriana" lastname="Kowalińska" birthdate="1993-03-19" gender="F" nation="POL" swrid="4086694" athleteid="4102">
              <RESULTS>
                <RESULT eventid="1094" points="714" reactiontime="+83" swimtime="00:02:37.41" resultid="4103" heatid="4290" lane="3" entrytime="00:02:31.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                    <SPLIT distance="150" swimtime="00:02:01.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="565" reactiontime="+72" swimtime="00:10:36.04" resultid="4104" heatid="4300" lane="5" entrytime="00:09:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="150" swimtime="00:01:55.68" />
                    <SPLIT distance="250" swimtime="00:03:15.84" />
                    <SPLIT distance="350" swimtime="00:04:36.53" />
                    <SPLIT distance="450" swimtime="00:05:57.21" />
                    <SPLIT distance="550" swimtime="00:07:17.95" />
                    <SPLIT distance="650" swimtime="00:08:38.37" />
                    <SPLIT distance="750" swimtime="00:09:57.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1335" points="685" reactiontime="+83" swimtime="00:02:33.16" resultid="4105" heatid="4354" lane="5" entrytime="00:02:30.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="602" reactiontime="+85" swimtime="00:00:31.17" resultid="4106" heatid="4375" lane="2" entrytime="00:00:30.89" />
                <RESULT eventid="1576" points="698" reactiontime="+76" swimtime="00:05:41.26" resultid="4107" heatid="4412" lane="5" entrytime="00:05:29.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:02:01.68" />
                    <SPLIT distance="200" swimtime="00:02:46.97" />
                    <SPLIT distance="250" swimtime="00:03:36.41" />
                    <SPLIT distance="300" swimtime="00:04:25.67" />
                    <SPLIT distance="350" swimtime="00:05:04.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="686" reactiontime="+85" swimtime="00:01:08.03" resultid="4108" heatid="4421" lane="6" entrytime="00:01:10.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="610" reactiontime="+71" swimtime="00:05:04.92" resultid="4109" heatid="4452" lane="5" entrytime="00:04:58.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:12.52" />
                    <SPLIT distance="150" swimtime="00:01:50.88" />
                    <SPLIT distance="200" swimtime="00:02:29.87" />
                    <SPLIT distance="250" swimtime="00:03:08.59" />
                    <SPLIT distance="300" swimtime="00:03:48.25" />
                    <SPLIT distance="350" swimtime="00:04:27.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Dąbrowski" birthdate="1974-01-14" gender="M" nation="POL" license="501713700022" swrid="5355776" athleteid="1899">
              <RESULTS>
                <RESULT eventid="1163" points="432" reactiontime="+94" swimtime="00:11:28.68" resultid="1900" heatid="4306" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:01:23.07" />
                    <SPLIT distance="150" swimtime="00:02:06.42" />
                    <SPLIT distance="200" swimtime="00:02:50.05" />
                    <SPLIT distance="250" swimtime="00:03:33.26" />
                    <SPLIT distance="300" swimtime="00:04:16.51" />
                    <SPLIT distance="350" swimtime="00:04:58.87" />
                    <SPLIT distance="400" swimtime="00:05:42.08" />
                    <SPLIT distance="450" swimtime="00:06:25.07" />
                    <SPLIT distance="500" swimtime="00:07:07.93" />
                    <SPLIT distance="550" swimtime="00:07:51.28" />
                    <SPLIT distance="600" swimtime="00:08:35.13" />
                    <SPLIT distance="650" swimtime="00:09:18.73" />
                    <SPLIT distance="700" swimtime="00:10:02.55" />
                    <SPLIT distance="750" swimtime="00:10:46.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="433" reactiontime="+77" swimtime="00:00:36.51" resultid="1901" heatid="4319" lane="3" />
                <RESULT eventid="1301" points="475" reactiontime="+79" swimtime="00:01:06.97" resultid="1902" heatid="4342" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="424" reactiontime="+75" swimtime="00:01:20.03" resultid="1903" heatid="4393" lane="2" entrytime="00:01:14.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="440" reactiontime="+87" swimtime="00:02:34.85" resultid="1904" heatid="4399" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:01:57.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="375" reactiontime="+84" swimtime="00:03:02.38" resultid="1905" heatid="4433" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:29.60" />
                    <SPLIT distance="150" swimtime="00:02:16.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="456" reactiontime="+82" swimtime="00:05:26.16" resultid="1906" heatid="4459" lane="4" entrytime="00:05:18.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:17.51" />
                    <SPLIT distance="150" swimtime="00:01:58.71" />
                    <SPLIT distance="200" swimtime="00:02:40.50" />
                    <SPLIT distance="250" swimtime="00:03:22.32" />
                    <SPLIT distance="300" swimtime="00:04:04.12" />
                    <SPLIT distance="350" swimtime="00:04:46.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Góralska" birthdate="1977-12-05" gender="F" nation="POL" athleteid="2760">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="2761" heatid="4269" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1146" status="DNS" swimtime="00:00:00.00" resultid="2762" heatid="4301" lane="4" entrytime="00:14:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jowita" lastname="Kucharska" birthdate="1980-02-15" gender="F" nation="POL" swrid="4313184" athleteid="4110">
              <RESULTS>
                <RESULT eventid="1646" points="324" reactiontime="+86" swimtime="00:03:28.51" resultid="4111" heatid="4430" lane="5" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                    <SPLIT distance="100" swimtime="00:01:41.96" />
                    <SPLIT distance="150" swimtime="00:02:37.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Drzewicka" birthdate="1976-10-26" gender="F" nation="POL" license="501713600017" swrid="5282851" athleteid="1825">
              <RESULTS>
                <RESULT eventid="1059" points="429" reactiontime="+84" swimtime="00:00:35.26" resultid="1826" heatid="4270" lane="2" entrytime="00:00:34.87" entrycourse="SCM" />
                <RESULT eventid="1215" points="542" reactiontime="+84" swimtime="00:00:38.04" resultid="1827" heatid="4316" lane="0" entrytime="00:00:36.36" entrycourse="SCM" />
                <RESULT eventid="1284" points="354" reactiontime="+90" swimtime="00:01:21.15" resultid="1828" heatid="4336" lane="8" />
                <RESULT eventid="1474" points="511" reactiontime="+72" swimtime="00:01:23.88" resultid="1829" heatid="4386" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Trzeszczkowski" birthdate="1980-09-13" gender="M" nation="POL" license="501713700021" swrid="5268961" athleteid="1907">
              <RESULTS>
                <RESULT eventid="1197" points="341" swimtime="00:23:30.10" resultid="1908" heatid="4311" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:14.39" />
                    <SPLIT distance="200" swimtime="00:03:02.26" />
                    <SPLIT distance="250" swimtime="00:03:50.08" />
                    <SPLIT distance="300" swimtime="00:04:37.50" />
                    <SPLIT distance="350" swimtime="00:05:24.79" />
                    <SPLIT distance="400" swimtime="00:06:12.19" />
                    <SPLIT distance="450" swimtime="00:06:59.56" />
                    <SPLIT distance="500" swimtime="00:07:46.88" />
                    <SPLIT distance="550" swimtime="00:08:34.97" />
                    <SPLIT distance="600" swimtime="00:09:23.25" />
                    <SPLIT distance="650" swimtime="00:10:11.20" />
                    <SPLIT distance="700" swimtime="00:10:59.24" />
                    <SPLIT distance="750" swimtime="00:11:46.85" />
                    <SPLIT distance="800" swimtime="00:12:34.49" />
                    <SPLIT distance="850" swimtime="00:13:22.02" />
                    <SPLIT distance="900" swimtime="00:14:10.19" />
                    <SPLIT distance="950" swimtime="00:14:57.79" />
                    <SPLIT distance="1000" swimtime="00:15:45.85" />
                    <SPLIT distance="1050" swimtime="00:16:33.58" />
                    <SPLIT distance="1100" swimtime="00:17:21.52" />
                    <SPLIT distance="1150" swimtime="00:18:09.01" />
                    <SPLIT distance="1200" swimtime="00:18:55.88" />
                    <SPLIT distance="1250" swimtime="00:19:42.63" />
                    <SPLIT distance="1300" swimtime="00:20:28.51" />
                    <SPLIT distance="1350" swimtime="00:21:14.83" />
                    <SPLIT distance="1400" swimtime="00:22:01.40" />
                    <SPLIT distance="1450" swimtime="00:22:46.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mieszko" lastname="Palmi-Kukiełko" birthdate="1993-09-15" gender="M" nation="POL" license="101713700006" swrid="4073437" athleteid="1869">
              <RESULTS>
                <RESULT eventid="1112" points="710" reactiontime="+72" swimtime="00:02:18.56" resultid="1870" heatid="4297" lane="5" entrytime="00:02:12.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                    <SPLIT distance="150" swimtime="00:01:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1197" points="646" reactiontime="+73" swimtime="00:18:46.48" resultid="1871" heatid="4309" lane="6" entrytime="00:17:45.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:06.40" />
                    <SPLIT distance="150" swimtime="00:01:42.84" />
                    <SPLIT distance="200" swimtime="00:02:19.92" />
                    <SPLIT distance="250" swimtime="00:02:57.22" />
                    <SPLIT distance="300" swimtime="00:03:35.18" />
                    <SPLIT distance="350" swimtime="00:04:13.05" />
                    <SPLIT distance="400" swimtime="00:04:51.42" />
                    <SPLIT distance="450" swimtime="00:05:29.86" />
                    <SPLIT distance="500" swimtime="00:06:08.09" />
                    <SPLIT distance="550" swimtime="00:06:46.24" />
                    <SPLIT distance="600" swimtime="00:07:24.17" />
                    <SPLIT distance="650" swimtime="00:08:01.62" />
                    <SPLIT distance="700" swimtime="00:08:38.91" />
                    <SPLIT distance="750" swimtime="00:09:16.43" />
                    <SPLIT distance="800" swimtime="00:09:54.32" />
                    <SPLIT distance="850" swimtime="00:10:31.82" />
                    <SPLIT distance="900" swimtime="00:11:09.87" />
                    <SPLIT distance="950" swimtime="00:11:47.69" />
                    <SPLIT distance="1000" swimtime="00:12:25.67" />
                    <SPLIT distance="1050" swimtime="00:13:03.73" />
                    <SPLIT distance="1100" swimtime="00:13:41.91" />
                    <SPLIT distance="1150" swimtime="00:14:20.30" />
                    <SPLIT distance="1200" swimtime="00:14:58.67" />
                    <SPLIT distance="1250" swimtime="00:15:37.03" />
                    <SPLIT distance="1300" swimtime="00:16:15.46" />
                    <SPLIT distance="1350" swimtime="00:16:53.84" />
                    <SPLIT distance="1400" swimtime="00:17:32.26" />
                    <SPLIT distance="1450" swimtime="00:18:09.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="678" reactiontime="+76" swimtime="00:00:57.43" resultid="1872" heatid="4352" lane="2" entrytime="00:00:54.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="616" reactiontime="+73" swimtime="00:02:22.19" resultid="1873" heatid="4357" lane="6" entrytime="00:02:27.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                    <SPLIT distance="150" swimtime="00:01:43.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="723" reactiontime="+74" swimtime="00:00:26.42" resultid="1874" heatid="4384" lane="3" entrytime="00:00:26.40" />
                <RESULT eventid="1593" points="732" reactiontime="+73" swimtime="00:04:59.59" resultid="1875" heatid="4414" lane="4" entrytime="00:04:49.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                    <SPLIT distance="100" swimtime="00:01:04.51" />
                    <SPLIT distance="150" swimtime="00:01:44.34" />
                    <SPLIT distance="200" swimtime="00:02:24.01" />
                    <SPLIT distance="250" swimtime="00:03:07.19" />
                    <SPLIT distance="300" swimtime="00:03:50.54" />
                    <SPLIT distance="350" swimtime="00:04:25.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="489" reactiontime="+81" swimtime="00:01:07.40" resultid="1876" heatid="4427" lane="5" entrytime="00:00:57.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="508" reactiontime="+76" swimtime="00:02:33.83" resultid="1877" heatid="4437" lane="5" entrytime="00:02:12.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:13.89" />
                    <SPLIT distance="150" swimtime="00:01:54.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Łagowska" birthdate="1982-06-07" gender="F" nation="POL" license="501713600008" athleteid="1808">
              <RESULTS>
                <RESULT eventid="1059" points="355" reactiontime="+87" swimtime="00:00:37.35" resultid="1809" heatid="4267" lane="1" />
                <RESULT eventid="1215" points="230" reactiontime="+101" swimtime="00:00:48.35" resultid="1810" heatid="4313" lane="9" />
                <RESULT eventid="1284" points="317" reactiontime="+88" swimtime="00:01:25.15" resultid="1811" heatid="4335" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="1812" heatid="4385" lane="5" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="1813" heatid="4395" lane="3" />
                <RESULT eventid="1646" points="237" reactiontime="+88" swimtime="00:03:51.38" resultid="1814" heatid="4429" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.39" />
                    <SPLIT distance="100" swimtime="00:01:48.75" />
                    <SPLIT distance="150" swimtime="00:02:51.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="259" reactiontime="+66" swimtime="00:06:52.65" resultid="1815" heatid="4454" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                    <SPLIT distance="100" swimtime="00:01:33.15" />
                    <SPLIT distance="150" swimtime="00:02:27.89" />
                    <SPLIT distance="200" swimtime="00:03:20.34" />
                    <SPLIT distance="250" swimtime="00:04:15.06" />
                    <SPLIT distance="300" swimtime="00:05:09.77" />
                    <SPLIT distance="350" swimtime="00:06:03.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Gregorowicz" birthdate="1974-10-30" gender="M" nation="POL" license="101713700002" swrid="4992729" athleteid="1844">
              <RESULTS>
                <RESULT eventid="1076" points="704" reactiontime="+71" swimtime="00:00:26.47" resultid="1845" heatid="4282" lane="8" entrytime="00:00:28.30" entrycourse="SCM" />
                <RESULT eventid="1163" points="707" reactiontime="+74" swimtime="00:09:44.53" resultid="1846" heatid="4303" lane="6" entrytime="00:09:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:09.12" />
                    <SPLIT distance="150" swimtime="00:01:45.65" />
                    <SPLIT distance="200" swimtime="00:02:22.38" />
                    <SPLIT distance="250" swimtime="00:02:59.36" />
                    <SPLIT distance="300" swimtime="00:03:36.36" />
                    <SPLIT distance="350" swimtime="00:04:13.24" />
                    <SPLIT distance="400" swimtime="00:04:50.11" />
                    <SPLIT distance="450" swimtime="00:05:27.26" />
                    <SPLIT distance="500" swimtime="00:06:04.48" />
                    <SPLIT distance="550" swimtime="00:06:41.95" />
                    <SPLIT distance="600" swimtime="00:07:19.15" />
                    <SPLIT distance="650" swimtime="00:07:56.36" />
                    <SPLIT distance="700" swimtime="00:08:32.99" />
                    <SPLIT distance="750" swimtime="00:09:09.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="667" reactiontime="+75" swimtime="00:02:25.25" resultid="1847" heatid="4357" lane="3" entrytime="00:02:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:10.06" />
                    <SPLIT distance="150" swimtime="00:01:48.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="721" reactiontime="+70" swimtime="00:00:28.15" resultid="1848" heatid="4377" lane="0" />
                <RESULT eventid="1593" points="707" reactiontime="+75" swimtime="00:05:18.56" resultid="1849" heatid="4414" lane="7" entrytime="00:05:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:09.69" />
                    <SPLIT distance="150" swimtime="00:01:55.75" />
                    <SPLIT distance="200" swimtime="00:02:39.10" />
                    <SPLIT distance="250" swimtime="00:03:24.39" />
                    <SPLIT distance="300" swimtime="00:04:08.43" />
                    <SPLIT distance="350" swimtime="00:04:44.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="776" reactiontime="+71" swimtime="00:01:01.87" resultid="1850" heatid="4427" lane="1" entrytime="00:01:01.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="723" reactiontime="+73" swimtime="00:04:39.79" resultid="1851" heatid="4456" lane="1" entrytime="00:04:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="150" swimtime="00:01:41.97" />
                    <SPLIT distance="200" swimtime="00:02:17.67" />
                    <SPLIT distance="250" swimtime="00:02:53.23" />
                    <SPLIT distance="300" swimtime="00:03:28.97" />
                    <SPLIT distance="350" swimtime="00:04:04.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Lemańczyk" birthdate="1977-10-01" gender="M" nation="POL" license="501713700050" athleteid="1837">
              <RESULTS>
                <RESULT eventid="1076" points="272" reactiontime="+82" swimtime="00:00:36.33" resultid="1838" heatid="4275" lane="0" />
                <RESULT eventid="1250" points="313" reactiontime="+90" swimtime="00:03:25.37" resultid="1839" heatid="4330" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                    <SPLIT distance="100" swimtime="00:01:40.50" />
                    <SPLIT distance="150" swimtime="00:02:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="261" reactiontime="+76" swimtime="00:01:21.74" resultid="1840" heatid="4342" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="343" reactiontime="+90" swimtime="00:01:32.55" resultid="1841" heatid="4367" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="312" reactiontime="+85" swimtime="00:02:53.65" resultid="1842" heatid="4400" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:21.33" />
                    <SPLIT distance="150" swimtime="00:02:06.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="293" reactiontime="+92" swimtime="00:06:17.81" resultid="1843" heatid="4463" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:01:26.96" />
                    <SPLIT distance="150" swimtime="00:02:15.10" />
                    <SPLIT distance="200" swimtime="00:03:05.07" />
                    <SPLIT distance="250" swimtime="00:03:54.02" />
                    <SPLIT distance="300" swimtime="00:04:42.55" />
                    <SPLIT distance="350" swimtime="00:05:30.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Gozdan" birthdate="1968-08-16" gender="M" nation="POL" license="501713700009" swrid="5230704" athleteid="1830">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="1831" heatid="4273" lane="4" />
                <RESULT eventid="1250" points="308" reactiontime="+84" swimtime="00:03:38.71" resultid="1832" heatid="4329" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                    <SPLIT distance="100" swimtime="00:01:36.74" />
                    <SPLIT distance="150" swimtime="00:02:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="296" reactiontime="+89" swimtime="00:01:21.25" resultid="1833" heatid="4343" lane="6" />
                <RESULT eventid="1406" points="329" reactiontime="+86" swimtime="00:01:36.20" resultid="1834" heatid="4366" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="243" reactiontime="+97" swimtime="00:03:09.98" resultid="1835" heatid="4399" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="100" swimtime="00:01:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="363" reactiontime="+92" swimtime="00:00:42.29" resultid="1836" heatid="4443" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Goździejewska" birthdate="1967-03-18" gender="F" nation="POL" license="501713600014" swrid="4313183" athleteid="1816">
              <RESULTS>
                <RESULT eventid="1059" points="522" reactiontime="+65" swimtime="00:00:35.14" resultid="1817" heatid="4270" lane="8" entrytime="00:00:35.06" entrycourse="SCM" />
                <RESULT eventid="1233" points="493" reactiontime="+87" swimtime="00:03:46.43" resultid="1819" heatid="4326" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.83" />
                    <SPLIT distance="100" swimtime="00:01:49.02" />
                    <SPLIT distance="150" swimtime="00:02:47.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="490" swimtime="00:01:18.67" resultid="1820" heatid="4337" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="503" swimtime="00:02:51.37" resultid="1821" heatid="4396" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                    <SPLIT distance="100" swimtime="00:01:23.43" />
                    <SPLIT distance="150" swimtime="00:02:08.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1576" points="353" swimtime="00:07:36.36" resultid="1822" heatid="4413" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.98" />
                    <SPLIT distance="100" swimtime="00:02:07.69" />
                    <SPLIT distance="150" swimtime="00:03:05.53" />
                    <SPLIT distance="200" swimtime="00:04:04.00" />
                    <SPLIT distance="250" swimtime="00:05:03.17" />
                    <SPLIT distance="300" swimtime="00:06:02.69" />
                    <SPLIT distance="350" swimtime="00:06:50.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="310" reactiontime="+102" swimtime="00:03:44.38" resultid="1823" heatid="4430" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                    <SPLIT distance="100" swimtime="00:01:47.84" />
                    <SPLIT distance="150" swimtime="00:02:46.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1731" points="452" swimtime="00:06:09.27" resultid="1824" heatid="4452" lane="9" entrytime="00:05:56.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:28.37" />
                    <SPLIT distance="150" swimtime="00:02:15.45" />
                    <SPLIT distance="200" swimtime="00:03:02.84" />
                    <SPLIT distance="250" swimtime="00:03:50.07" />
                    <SPLIT distance="300" swimtime="00:04:36.78" />
                    <SPLIT distance="350" swimtime="00:05:23.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="498" reactiontime="+86" swimtime="00:12:17.50" resultid="4091" heatid="4300" lane="6" entrytime="00:11:59.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:23.72" />
                    <SPLIT distance="150" swimtime="00:02:09.36" />
                    <SPLIT distance="200" swimtime="00:02:55.03" />
                    <SPLIT distance="250" swimtime="00:03:41.10" />
                    <SPLIT distance="300" swimtime="00:04:26.90" />
                    <SPLIT distance="350" swimtime="00:05:13.53" />
                    <SPLIT distance="400" swimtime="00:06:00.39" />
                    <SPLIT distance="450" swimtime="00:06:48.09" />
                    <SPLIT distance="500" swimtime="00:07:35.02" />
                    <SPLIT distance="550" swimtime="00:08:23.02" />
                    <SPLIT distance="600" swimtime="00:09:09.70" />
                    <SPLIT distance="650" swimtime="00:09:57.33" />
                    <SPLIT distance="700" swimtime="00:10:44.35" />
                    <SPLIT distance="750" swimtime="00:11:32.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Łuczak" birthdate="1978-03-18" gender="M" nation="POL" license="501713700016" swrid="5416815" athleteid="1909">
              <RESULTS>
                <RESULT eventid="1250" points="391" reactiontime="+69" swimtime="00:03:09.48" resultid="1910" heatid="4333" lane="7" entrytime="00:02:57.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:01:31.49" />
                    <SPLIT distance="150" swimtime="00:02:21.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="450" reactiontime="+67" swimtime="00:01:22.97" resultid="1911" heatid="4369" lane="5" entrytime="00:01:20.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="508" reactiontime="+75" swimtime="00:00:36.15" resultid="1912" heatid="4448" lane="0" entrytime="00:00:34.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Matusiak vel Matuszewski" birthdate="1974-06-25" gender="M" nation="POL" license="501713700004" athleteid="1852">
              <RESULTS>
                <RESULT eventid="1076" points="329" reactiontime="+84" swimtime="00:00:34.13" resultid="1853" heatid="4273" lane="7" />
                <RESULT eventid="1267" points="270" reactiontime="+70" swimtime="00:00:42.75" resultid="1855" heatid="4318" lane="3" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="1856" heatid="4343" lane="1" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="1857" heatid="4376" lane="5" />
                <RESULT eventid="1525" points="339" reactiontime="+81" swimtime="00:02:48.80" resultid="1858" heatid="4400" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:19.97" />
                    <SPLIT distance="150" swimtime="00:02:03.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="1859" heatid="4463" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Konopacki" birthdate="1978-04-01" gender="M" nation="POL" license="501713700019" swrid="5282843" athleteid="1860">
              <RESULTS>
                <RESULT eventid="1076" points="586" reactiontime="+80" swimtime="00:00:27.78" resultid="1861" heatid="4275" lane="9" />
                <RESULT eventid="1197" points="566" reactiontime="+71" swimtime="00:19:50.54" resultid="1862" heatid="4309" lane="2" entrytime="00:19:03.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                    <SPLIT distance="200" swimtime="00:02:32.96" />
                    <SPLIT distance="250" swimtime="00:03:12.64" />
                    <SPLIT distance="300" swimtime="00:03:52.81" />
                    <SPLIT distance="350" swimtime="00:04:33.50" />
                    <SPLIT distance="400" swimtime="00:05:13.85" />
                    <SPLIT distance="450" swimtime="00:05:54.57" />
                    <SPLIT distance="500" swimtime="00:06:34.71" />
                    <SPLIT distance="550" swimtime="00:07:15.04" />
                    <SPLIT distance="600" swimtime="00:07:54.68" />
                    <SPLIT distance="650" swimtime="00:08:34.87" />
                    <SPLIT distance="700" swimtime="00:09:14.53" />
                    <SPLIT distance="750" swimtime="00:09:54.55" />
                    <SPLIT distance="800" swimtime="00:10:34.22" />
                    <SPLIT distance="850" swimtime="00:11:14.51" />
                    <SPLIT distance="900" swimtime="00:11:54.60" />
                    <SPLIT distance="950" swimtime="00:12:34.62" />
                    <SPLIT distance="1000" swimtime="00:13:14.77" />
                    <SPLIT distance="1050" swimtime="00:13:54.59" />
                    <SPLIT distance="1100" swimtime="00:14:34.59" />
                    <SPLIT distance="1150" swimtime="00:15:14.68" />
                    <SPLIT distance="1200" swimtime="00:15:54.66" />
                    <SPLIT distance="1250" swimtime="00:16:35.07" />
                    <SPLIT distance="1300" swimtime="00:17:14.49" />
                    <SPLIT distance="1350" swimtime="00:17:54.10" />
                    <SPLIT distance="1400" swimtime="00:18:33.79" />
                    <SPLIT distance="1450" swimtime="00:19:12.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="511" reactiontime="+73" swimtime="00:00:33.93" resultid="1863" heatid="4324" lane="4" entrytime="00:00:31.94" entrycourse="SCM" />
                <RESULT eventid="1301" points="556" reactiontime="+69" swimtime="00:01:02.27" resultid="1864" heatid="4341" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="585" reactiontime="+61" swimtime="00:02:15.88" resultid="1865" heatid="4406" lane="1" entrytime="00:02:14.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                    <SPLIT distance="150" swimtime="00:01:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="555" reactiontime="+69" swimtime="00:05:44.27" resultid="1866" heatid="4417" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                    <SPLIT distance="100" swimtime="00:01:23.61" />
                    <SPLIT distance="150" swimtime="00:02:08.18" />
                    <SPLIT distance="200" swimtime="00:02:52.55" />
                    <SPLIT distance="250" swimtime="00:03:43.24" />
                    <SPLIT distance="300" swimtime="00:04:32.37" />
                    <SPLIT distance="350" swimtime="00:05:08.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="464" reactiontime="+77" swimtime="00:02:45.43" resultid="1867" heatid="4437" lane="8" entrytime="00:02:35.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:02:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="566" reactiontime="+72" swimtime="00:04:58.30" resultid="1868" heatid="4457" lane="3" entrytime="00:04:48.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:10.52" />
                    <SPLIT distance="150" swimtime="00:01:48.50" />
                    <SPLIT distance="200" swimtime="00:02:26.99" />
                    <SPLIT distance="250" swimtime="00:03:05.18" />
                    <SPLIT distance="300" swimtime="00:03:44.09" />
                    <SPLIT distance="350" swimtime="00:04:22.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kieres" birthdate="1984-06-13" gender="M" nation="POL" license="101713700001" swrid="5282844" athleteid="1891">
              <RESULTS>
                <RESULT eventid="1112" status="DNS" swimtime="00:00:00.00" resultid="1892" heatid="4291" lane="1" />
                <RESULT eventid="1250" points="383" reactiontime="+75" swimtime="00:03:13.13" resultid="1893" heatid="4332" lane="3" entrytime="00:03:01.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="100" swimtime="00:01:29.30" />
                    <SPLIT distance="150" swimtime="00:02:20.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="274" reactiontime="+82" swimtime="00:03:08.68" resultid="1894" heatid="4356" lane="4" entrytime="00:02:55.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:20.64" />
                    <SPLIT distance="150" swimtime="00:02:13.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="339" reactiontime="+72" swimtime="00:01:29.53" resultid="1895" heatid="4367" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="333" reactiontime="+73" swimtime="00:00:34.82" resultid="1896" heatid="4378" lane="0" />
                <RESULT eventid="1629" points="355" reactiontime="+71" swimtime="00:01:15.79" resultid="1897" heatid="4424" lane="4" entrytime="00:01:15.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="326" reactiontime="+79" swimtime="00:00:41.35" resultid="1898" heatid="4446" lane="2" entrytime="00:00:37.29" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1386" points="531" reactiontime="+68" swimtime="00:02:06.37" resultid="1920" heatid="4493" lane="6" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:10.51" />
                    <SPLIT distance="150" swimtime="00:01:39.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1869" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="1837" number="2" />
                    <RELAYPOSITION athleteid="1844" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="2771" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="1924" heatid="4497" lane="7" entrytime="00:01:49.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1869" number="1" />
                    <RELAYPOSITION athleteid="1844" number="2" />
                    <RELAYPOSITION athleteid="1878" number="3" />
                    <RELAYPOSITION athleteid="2771" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1386" points="483" reactiontime="+73" swimtime="00:02:14.41" resultid="1921" heatid="4492" lane="4" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:46.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1899" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="1909" number="2" />
                    <RELAYPOSITION athleteid="1891" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="1860" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" points="507" reactiontime="+77" swimtime="00:01:59.07" resultid="1925" heatid="4496" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="100" swimtime="00:00:59.67" />
                    <SPLIT distance="150" swimtime="00:01:26.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1860" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="1909" number="2" />
                    <RELAYPOSITION athleteid="1899" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="1891" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1386" points="365" reactiontime="+66" swimtime="00:02:35.07" resultid="1922" heatid="4492" lane="3" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                    <SPLIT distance="100" swimtime="00:01:23.92" />
                    <SPLIT distance="150" swimtime="00:02:01.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1852" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="1830" number="2" />
                    <RELAYPOSITION athleteid="1913" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="1885" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" points="383" reactiontime="+99" swimtime="00:02:15.31" resultid="1926" heatid="4496" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:07.75" />
                    <SPLIT distance="150" swimtime="00:01:41.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1885" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="1913" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="1852" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="1837" number="4" reactiontime="-10" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1369" points="488" swimtime="00:02:38.42" resultid="1919" heatid="4490" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="150" swimtime="00:01:59.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1825" number="1" />
                    <RELAYPOSITION athleteid="1816" number="2" />
                    <RELAYPOSITION athleteid="4102" number="3" />
                    <RELAYPOSITION athleteid="1808" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1542" status="DNS" swimtime="00:00:00.00" resultid="1923" heatid="4494" lane="3" entrytime="00:02:18.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4102" number="1" />
                    <RELAYPOSITION athleteid="1825" number="2" />
                    <RELAYPOSITION athleteid="4110" number="3" />
                    <RELAYPOSITION athleteid="1808" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" points="583" reactiontime="+75" swimtime="00:01:59.90" resultid="1917" heatid="4489" lane="6" entrytime="00:01:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.27" />
                    <SPLIT distance="100" swimtime="00:00:55.00" />
                    <SPLIT distance="150" swimtime="00:01:25.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1869" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="1844" number="2" reactiontime="+15" />
                    <RELAYPOSITION athleteid="4102" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="1825" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1714" points="592" reactiontime="+84" swimtime="00:02:11.91" resultid="1927" heatid="4499" lane="3" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="150" swimtime="00:01:44.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1825" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="1869" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="4102" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="1844" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1129" points="466" reactiontime="+80" swimtime="00:02:11.91" resultid="1918" heatid="4489" lane="2" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                    <SPLIT distance="100" swimtime="00:00:57.77" />
                    <SPLIT distance="150" swimtime="00:01:34.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1899" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="1860" number="2" />
                    <RELAYPOSITION athleteid="1816" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="1808" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1714" points="460" reactiontime="+66" swimtime="00:02:26.74" resultid="1928" heatid="4498" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:22.33" />
                    <SPLIT distance="150" swimtime="00:01:52.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1860" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="1816" number="2" />
                    <RELAYPOSITION athleteid="2771" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4110" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3449" name="RMKS Rybnik">
          <CONTACT email="aniaduda0511@tlen.pl" name="Duda Anna" phone="792666159" />
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Duda" birthdate="1981-04-15" gender="F" nation="POL" athleteid="3450">
              <RESULTS>
                <RESULT eventid="1059" points="762" reactiontime="+75" swimtime="00:00:28.95" resultid="3451" heatid="4272" lane="1" entrytime="00:00:28.80" />
                <RESULT eventid="1094" points="629" reactiontime="+86" swimtime="00:02:49.31" resultid="3452" heatid="4290" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:18.81" />
                    <SPLIT distance="150" swimtime="00:02:11.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="499" reactiontime="+72" swimtime="00:00:37.35" resultid="3453" heatid="4315" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1284" points="677" reactiontime="+80" swimtime="00:01:06.09" resultid="3454" heatid="4340" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1440" points="798" reactiontime="+71" swimtime="00:00:30.58" resultid="3455" heatid="4375" lane="3" entrytime="00:00:29.80" />
                <RESULT eventid="1474" points="427" reactiontime="+68" swimtime="00:01:25.92" resultid="3456" heatid="4388" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" status="DNS" swimtime="00:00:00.00" resultid="3457" heatid="4441" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12914" nation="POL" region="14" clubid="2642" name="Water Squad">
          <CONTACT email="agnieszka.kaczmarek85@gmail.com" name="Kaczmarek Agnieszka" phone="531799855" />
          <ATHLETES>
            <ATHLETE firstname="Karolina" lastname="Szyszkowska" birthdate="1996-11-05" gender="F" nation="POL" athleteid="2789">
              <RESULTS>
                <RESULT eventid="1059" points="704" reactiontime="+84" swimtime="00:00:28.57" resultid="2790" heatid="4272" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="1233" points="744" reactiontime="+88" swimtime="00:02:51.60" resultid="2791" heatid="4328" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:22.91" />
                    <SPLIT distance="150" swimtime="00:02:06.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="726" reactiontime="+86" swimtime="00:01:18.51" resultid="2792" heatid="4365" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="706" reactiontime="+81" swimtime="00:00:35.48" resultid="2793" heatid="4441" lane="4" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kulisz" birthdate="1977-06-16" gender="M" nation="POL" license="512914700002" swrid="5416809" athleteid="2649">
              <RESULTS>
                <RESULT eventid="1076" points="441" reactiontime="+79" swimtime="00:00:30.93" resultid="2650" heatid="4279" lane="6" entrytime="00:00:31.48" entrycourse="LCM" />
                <RESULT eventid="1301" points="428" reactiontime="+78" swimtime="00:01:09.31" resultid="2651" heatid="4346" lane="3" entrytime="00:01:12.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="438" reactiontime="+88" swimtime="00:00:33.23" resultid="2652" heatid="4377" lane="8" />
                <RESULT eventid="1525" points="413" reactiontime="+81" swimtime="00:02:38.12" resultid="2653" heatid="4403" lane="7" entrytime="00:02:40.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                    <SPLIT distance="150" swimtime="00:01:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="363" reactiontime="+86" swimtime="00:00:40.97" resultid="2654" heatid="4443" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Korpetta" birthdate="1959-12-27" gender="M" nation="POL" license="112914700013" swrid="4754654" athleteid="2655">
              <RESULTS>
                <RESULT eventid="1076" points="363" reactiontime="+99" swimtime="00:00:35.36" resultid="2656" heatid="4274" lane="9" />
                <RESULT eventid="1163" points="370" reactiontime="+99" swimtime="00:13:13.40" resultid="2657" heatid="4307" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                    <SPLIT distance="100" swimtime="00:01:29.42" />
                    <SPLIT distance="150" swimtime="00:02:19.25" />
                    <SPLIT distance="200" swimtime="00:03:10.80" />
                    <SPLIT distance="250" swimtime="00:04:02.48" />
                    <SPLIT distance="300" swimtime="00:04:55.15" />
                    <SPLIT distance="350" swimtime="00:05:47.55" />
                    <SPLIT distance="400" swimtime="00:06:39.40" />
                    <SPLIT distance="450" swimtime="00:07:30.27" />
                    <SPLIT distance="500" swimtime="00:08:22.03" />
                    <SPLIT distance="550" swimtime="00:09:12.84" />
                    <SPLIT distance="600" swimtime="00:10:04.00" />
                    <SPLIT distance="650" swimtime="00:10:53.98" />
                    <SPLIT distance="700" swimtime="00:11:43.76" />
                    <SPLIT distance="750" swimtime="00:12:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="331" reactiontime="+71" swimtime="00:00:44.24" resultid="2658" heatid="4318" lane="4" />
                <RESULT eventid="1301" points="391" reactiontime="+100" swimtime="00:01:19.01" resultid="2659" heatid="4342" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="2660" heatid="4399" lane="5" />
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="2661" heatid="4418" lane="5" />
                <RESULT eventid="1663" points="355" reactiontime="+69" swimtime="00:03:26.45" resultid="2662" heatid="4432" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                    <SPLIT distance="100" swimtime="00:01:39.46" />
                    <SPLIT distance="150" swimtime="00:02:34.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="381" reactiontime="+102" swimtime="00:06:21.79" resultid="2663" heatid="4462" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:28.19" />
                    <SPLIT distance="150" swimtime="00:02:17.68" />
                    <SPLIT distance="200" swimtime="00:03:07.42" />
                    <SPLIT distance="250" swimtime="00:05:37.50" />
                    <SPLIT distance="300" swimtime="00:06:21.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Markowski" birthdate="1976-01-04" gender="M" nation="POL" license="512914700011" swrid="5471789" athleteid="2669">
              <RESULTS>
                <RESULT eventid="1112" points="525" reactiontime="+79" swimtime="00:02:41.27" resultid="2670" heatid="4291" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:15.67" />
                    <SPLIT distance="150" swimtime="00:02:02.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="543" reactiontime="+81" swimtime="00:00:30.94" resultid="2671" heatid="4381" lane="7" entrytime="00:00:31.47" entrycourse="LCM" />
                <RESULT eventid="1491" points="502" reactiontime="+88" swimtime="00:01:15.67" resultid="2672" heatid="4393" lane="8" entrytime="00:01:16.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="558" reactiontime="+68" swimtime="00:01:09.07" resultid="2673" heatid="4426" lane="9" entrytime="00:01:08.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="502" reactiontime="+62" swimtime="00:02:45.54" resultid="2674" heatid="4436" lane="0" entrytime="00:02:46.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:20.99" />
                    <SPLIT distance="150" swimtime="00:02:03.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kośmider" birthdate="1966-03-01" gender="M" nation="POL" swrid="4992964" athleteid="2802">
              <RESULTS>
                <RESULT eventid="1076" points="502" reactiontime="+72" swimtime="00:00:30.77" resultid="2803" heatid="4281" lane="0" entrytime="00:00:29.50" />
                <RESULT eventid="1163" points="515" reactiontime="+76" swimtime="00:11:13.81" resultid="2804" heatid="4304" lane="8" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                    <SPLIT distance="100" swimtime="00:01:20.39" />
                    <SPLIT distance="150" swimtime="00:02:02.30" />
                    <SPLIT distance="200" swimtime="00:02:44.72" />
                    <SPLIT distance="250" swimtime="00:03:27.53" />
                    <SPLIT distance="300" swimtime="00:04:10.62" />
                    <SPLIT distance="350" swimtime="00:04:53.07" />
                    <SPLIT distance="400" swimtime="00:05:35.96" />
                    <SPLIT distance="450" swimtime="00:06:18.03" />
                    <SPLIT distance="500" swimtime="00:07:00.20" />
                    <SPLIT distance="550" swimtime="00:07:42.14" />
                    <SPLIT distance="600" swimtime="00:08:24.59" />
                    <SPLIT distance="650" swimtime="00:09:07.30" />
                    <SPLIT distance="700" swimtime="00:09:49.96" />
                    <SPLIT distance="750" swimtime="00:10:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="511" reactiontime="+72" swimtime="00:03:08.44" resultid="2805" heatid="4332" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:28.67" />
                    <SPLIT distance="150" swimtime="00:02:16.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="477" reactiontime="+78" swimtime="00:01:26.60" resultid="2806" heatid="4370" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="520" reactiontime="+81" swimtime="00:06:15.37" resultid="2807" heatid="4415" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                    <SPLIT distance="100" swimtime="00:01:34.79" />
                    <SPLIT distance="150" swimtime="00:02:26.44" />
                    <SPLIT distance="200" swimtime="00:03:13.47" />
                    <SPLIT distance="250" swimtime="00:04:02.72" />
                    <SPLIT distance="300" swimtime="00:04:52.99" />
                    <SPLIT distance="350" swimtime="00:05:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="527" reactiontime="+75" swimtime="00:00:37.17" resultid="2808" heatid="4446" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1748" points="530" reactiontime="+81" swimtime="00:05:24.41" resultid="2809" heatid="4457" lane="9" entrytime="00:05:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:01:57.56" />
                    <SPLIT distance="200" swimtime="00:02:39.51" />
                    <SPLIT distance="250" swimtime="00:03:20.58" />
                    <SPLIT distance="300" swimtime="00:04:02.37" />
                    <SPLIT distance="350" swimtime="00:04:44.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Dolińska" birthdate="1990-07-06" gender="F" nation="POL" license="512914600056" swrid="4251116" athleteid="2643">
              <RESULTS>
                <RESULT eventid="1059" points="466" reactiontime="+89" swimtime="00:00:33.19" resultid="2644" heatid="4268" lane="9" />
                <RESULT eventid="1215" points="252" reactiontime="+84" swimtime="00:00:45.26" resultid="2645" heatid="4312" lane="6" />
                <RESULT eventid="1284" points="394" reactiontime="+102" swimtime="00:01:15.36" resultid="2646" heatid="4335" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="248" reactiontime="+98" swimtime="00:01:38.37" resultid="2647" heatid="4386" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="364" reactiontime="+112" swimtime="00:02:51.32" resultid="2648" heatid="4395" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="100" swimtime="00:01:23.04" />
                    <SPLIT distance="150" swimtime="00:02:08.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Żemier" birthdate="1982-11-09" gender="M" nation="POL" athleteid="2780">
              <RESULTS>
                <RESULT eventid="1076" points="679" reactiontime="+79" swimtime="00:00:26.45" resultid="2781" heatid="4285" lane="9" entrytime="00:00:26.65" />
                <RESULT eventid="1112" points="737" reactiontime="+75" swimtime="00:02:24.63" resultid="2782" heatid="4297" lane="7" entrytime="00:02:21.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                    <SPLIT distance="100" swimtime="00:01:06.86" />
                    <SPLIT distance="150" swimtime="00:01:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="758" reactiontime="+66" swimtime="00:00:29.76" resultid="2783" heatid="4325" lane="5" entrytime="00:00:29.81" />
                <RESULT eventid="1301" points="685" reactiontime="+76" swimtime="00:00:58.09" resultid="2784" heatid="4351" lane="7" entrytime="00:00:57.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="706" reactiontime="+77" swimtime="00:00:28.15" resultid="2785" heatid="4383" lane="2" entrytime="00:00:28.81" />
                <RESULT eventid="1491" points="736" reactiontime="+66" swimtime="00:01:04.75" resultid="2786" heatid="4394" lane="5" entrytime="00:01:03.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="691" reactiontime="+76" swimtime="00:01:03.54" resultid="2787" heatid="4427" lane="9" entrytime="00:01:02.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="649" reactiontime="+64" swimtime="00:02:27.93" resultid="2788" heatid="4437" lane="3" entrytime="00:02:21.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:10.30" />
                    <SPLIT distance="150" swimtime="00:01:49.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Brożyna" birthdate="1980-04-28" gender="M" nation="POL" license="512914700006" swrid="5312396" athleteid="2675">
              <RESULTS>
                <RESULT eventid="1112" points="499" reactiontime="+91" swimtime="00:02:44.74" resultid="2676" heatid="4292" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                    <SPLIT distance="150" swimtime="00:02:06.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="469" reactiontime="+65" swimtime="00:00:34.91" resultid="2677" heatid="4323" lane="0" entrytime="00:00:35.40" entrycourse="LCM" />
                <RESULT eventid="1491" points="469" reactiontime="+71" swimtime="00:01:15.21" resultid="2678" heatid="4393" lane="1" entrytime="00:01:16.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="473" reactiontime="+85" swimtime="00:06:03.22" resultid="2679" heatid="4418" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:01:29.57" />
                    <SPLIT distance="150" swimtime="00:02:13.61" />
                    <SPLIT distance="200" swimtime="00:02:57.07" />
                    <SPLIT distance="250" swimtime="00:03:48.70" />
                    <SPLIT distance="300" swimtime="00:04:40.68" />
                    <SPLIT distance="350" swimtime="00:05:22.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="464" reactiontime="+70" swimtime="00:02:45.43" resultid="2680" heatid="4436" lane="7" entrytime="00:02:41.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:22.26" />
                    <SPLIT distance="150" swimtime="00:02:05.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="450" reactiontime="+89" swimtime="00:05:22.07" resultid="2681" heatid="4463" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:14.84" />
                    <SPLIT distance="150" swimtime="00:01:55.82" />
                    <SPLIT distance="200" swimtime="00:02:36.81" />
                    <SPLIT distance="250" swimtime="00:03:18.70" />
                    <SPLIT distance="300" swimtime="00:04:00.60" />
                    <SPLIT distance="350" swimtime="00:04:42.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Romuald" lastname="Kozłowski" birthdate="1966-08-13" gender="M" nation="POL" license="512914700012" swrid="5425564" athleteid="2664">
              <RESULTS>
                <RESULT eventid="1076" points="621" reactiontime="+79" swimtime="00:00:28.66" resultid="2665" heatid="4273" lane="6" />
                <RESULT eventid="1250" points="493" reactiontime="+88" swimtime="00:03:10.68" resultid="2666" heatid="4329" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:01:25.02" />
                    <SPLIT distance="150" swimtime="00:02:16.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="586" reactiontime="+85" swimtime="00:01:20.85" resultid="2667" heatid="4370" lane="2" entrytime="00:01:17.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="617" reactiontime="+82" swimtime="00:00:35.27" resultid="2668" heatid="4447" lane="5" entrytime="00:00:34.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Fluder" birthdate="1986-03-01" gender="M" nation="POL" athleteid="2794">
              <RESULTS>
                <RESULT eventid="1076" points="641" reactiontime="+71" swimtime="00:00:26.40" resultid="2795" heatid="4286" lane="0" entrytime="00:00:25.99" />
                <RESULT eventid="1197" points="657" reactiontime="+83" swimtime="00:18:24.42" resultid="2796" heatid="4309" lane="4" entrytime="00:17:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:06.45" />
                    <SPLIT distance="150" swimtime="00:01:42.86" />
                    <SPLIT distance="200" swimtime="00:02:19.46" />
                    <SPLIT distance="250" swimtime="00:02:55.78" />
                    <SPLIT distance="300" swimtime="00:03:32.61" />
                    <SPLIT distance="350" swimtime="00:04:09.31" />
                    <SPLIT distance="400" swimtime="00:04:46.27" />
                    <SPLIT distance="450" swimtime="00:05:23.18" />
                    <SPLIT distance="500" swimtime="00:06:00.04" />
                    <SPLIT distance="550" swimtime="00:07:51.24" />
                    <SPLIT distance="600" swimtime="00:07:13.91" />
                    <SPLIT distance="650" swimtime="00:09:05.37" />
                    <SPLIT distance="700" swimtime="00:08:28.25" />
                    <SPLIT distance="750" swimtime="00:10:20.52" />
                    <SPLIT distance="800" swimtime="00:09:42.93" />
                    <SPLIT distance="850" swimtime="00:11:35.17" />
                    <SPLIT distance="900" swimtime="00:10:57.79" />
                    <SPLIT distance="950" swimtime="00:12:50.28" />
                    <SPLIT distance="1000" swimtime="00:12:12.70" />
                    <SPLIT distance="1050" swimtime="00:14:06.12" />
                    <SPLIT distance="1100" swimtime="00:15:58.68" />
                    <SPLIT distance="1150" swimtime="00:15:21.16" />
                    <SPLIT distance="1200" swimtime="00:18:24.42" />
                    <SPLIT distance="1250" swimtime="00:16:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="711" reactiontime="+77" swimtime="00:00:56.90" resultid="2797" heatid="4352" lane="7" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="594" reactiontime="+76" swimtime="00:00:28.72" resultid="2798" heatid="4383" lane="6" entrytime="00:00:28.70" />
                <RESULT eventid="1525" points="695" reactiontime="+85" swimtime="00:02:07.39" resultid="2799" heatid="4407" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:02.01" />
                    <SPLIT distance="150" swimtime="00:01:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="546" reactiontime="+86" swimtime="00:01:05.65" resultid="2800" heatid="4427" lane="0" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="732" reactiontime="+88" swimtime="00:04:32.86" resultid="2801" heatid="4456" lane="5" entrytime="00:04:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:05.12" />
                    <SPLIT distance="150" swimtime="00:01:40.13" />
                    <SPLIT distance="200" swimtime="00:02:15.09" />
                    <SPLIT distance="250" swimtime="00:02:49.26" />
                    <SPLIT distance="300" swimtime="00:03:24.32" />
                    <SPLIT distance="350" swimtime="00:03:59.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arkadiusz" lastname="Aptewicz" birthdate="1993-12-20" gender="M" nation="POL" athleteid="2775">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1197" points="837" reactiontime="+67" swimtime="00:17:13.46" resultid="2776" heatid="4309" lane="3" entrytime="00:17:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="100" swimtime="00:01:03.59" />
                    <SPLIT distance="150" swimtime="00:01:38.53" />
                    <SPLIT distance="200" swimtime="00:02:13.27" />
                    <SPLIT distance="250" swimtime="00:02:47.91" />
                    <SPLIT distance="300" swimtime="00:03:22.41" />
                    <SPLIT distance="350" swimtime="00:03:57.04" />
                    <SPLIT distance="400" swimtime="00:04:31.32" />
                    <SPLIT distance="450" swimtime="00:05:05.86" />
                    <SPLIT distance="500" swimtime="00:05:40.28" />
                    <SPLIT distance="550" swimtime="00:06:14.88" />
                    <SPLIT distance="600" swimtime="00:06:49.20" />
                    <SPLIT distance="650" swimtime="00:07:23.91" />
                    <SPLIT distance="700" swimtime="00:07:58.49" />
                    <SPLIT distance="750" swimtime="00:08:33.04" />
                    <SPLIT distance="800" swimtime="00:09:07.91" />
                    <SPLIT distance="850" swimtime="00:09:42.97" />
                    <SPLIT distance="900" swimtime="00:10:17.71" />
                    <SPLIT distance="950" swimtime="00:10:52.58" />
                    <SPLIT distance="1000" swimtime="00:11:27.38" />
                    <SPLIT distance="1050" swimtime="00:12:02.28" />
                    <SPLIT distance="1100" swimtime="00:12:37.29" />
                    <SPLIT distance="1150" swimtime="00:13:12.01" />
                    <SPLIT distance="1200" swimtime="00:13:47.03" />
                    <SPLIT distance="1250" swimtime="00:14:21.92" />
                    <SPLIT distance="1300" swimtime="00:14:56.95" />
                    <SPLIT distance="1350" swimtime="00:15:31.89" />
                    <SPLIT distance="1400" swimtime="00:16:06.47" />
                    <SPLIT distance="1450" swimtime="00:16:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="667" reactiontime="+68" swimtime="00:02:30.82" resultid="2777" heatid="4334" lane="4" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:51.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="758" reactiontime="+70" swimtime="00:04:56.24" resultid="2778" heatid="4414" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:06.71" />
                    <SPLIT distance="150" swimtime="00:01:49.11" />
                    <SPLIT distance="200" swimtime="00:02:29.49" />
                    <SPLIT distance="250" swimtime="00:03:09.40" />
                    <SPLIT distance="300" swimtime="00:03:50.18" />
                    <SPLIT distance="350" swimtime="00:04:24.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="823" reactiontime="+64" swimtime="00:04:17.17" resultid="2779" heatid="4456" lane="4" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                    <SPLIT distance="100" swimtime="00:01:00.32" />
                    <SPLIT distance="150" swimtime="00:01:33.03" />
                    <SPLIT distance="200" swimtime="00:02:05.96" />
                    <SPLIT distance="250" swimtime="00:02:38.72" />
                    <SPLIT distance="300" swimtime="00:03:11.78" />
                    <SPLIT distance="350" swimtime="00:03:45.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1386" points="716" reactiontime="+69" swimtime="00:01:57.87" resultid="5044" heatid="4491" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="100" swimtime="00:01:04.94" />
                    <SPLIT distance="150" swimtime="00:01:32.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2780" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2664" number="2" />
                    <RELAYPOSITION athleteid="2794" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="2775" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1559" points="704" reactiontime="+77" swimtime="00:01:46.72" resultid="5047" heatid="4495" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.97" />
                    <SPLIT distance="100" swimtime="00:00:54.48" />
                    <SPLIT distance="150" swimtime="00:01:21.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2780" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2664" number="2" />
                    <RELAYPOSITION athleteid="2794" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="2775" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M">
              <RESULTS>
                <RESULT eventid="1559" points="471" reactiontime="+76" swimtime="00:02:06.27" resultid="5046" heatid="4495" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:00:59.86" />
                    <SPLIT distance="150" swimtime="00:01:30.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2675" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2802" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="2669" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="2655" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Water Squad 2">
              <RESULTS>
                <RESULT eventid="1386" points="492" reactiontime="+76" swimtime="00:02:20.37" resultid="5045" heatid="4492" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:11.62" />
                    <SPLIT distance="150" swimtime="00:01:45.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2675" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2802" number="2" />
                    <RELAYPOSITION athleteid="2649" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="2655" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X">
              <RESULTS>
                <RESULT eventid="1129" points="684" reactiontime="+91" swimtime="00:01:53.67" resultid="5038" heatid="4488" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:00.62" />
                    <SPLIT distance="150" swimtime="00:01:25.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2643" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="2789" number="2" />
                    <RELAYPOSITION athleteid="2775" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="2780" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3103" name="Masters Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos" phone="604184311" />
          <ATHLETES>
            <ATHLETE firstname="Przemysław" lastname="Michniewski" birthdate="1983-04-11" gender="M" nation="POL" license="503605700012" athleteid="3133">
              <RESULTS>
                <RESULT eventid="1076" points="564" reactiontime="+81" swimtime="00:00:27.55" resultid="3134" heatid="4282" lane="6" entrytime="00:00:28.10" />
                <RESULT eventid="1112" points="475" reactiontime="+76" swimtime="00:02:41.09" resultid="3135" heatid="4294" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:15.39" />
                    <SPLIT distance="150" swimtime="00:02:01.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="529" reactiontime="+84" swimtime="00:02:53.44" resultid="3136" heatid="4333" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="100" swimtime="00:01:22.20" />
                    <SPLIT distance="150" swimtime="00:02:08.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="527" reactiontime="+84" swimtime="00:01:17.26" resultid="3137" heatid="4370" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="551" reactiontime="+80" swimtime="00:00:34.73" resultid="3138" heatid="4447" lane="6" entrytime="00:00:35.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Olejarczyk" birthdate="1979-06-12" gender="M" nation="POL" license="503605700007" swrid="4992959" athleteid="3126">
              <RESULTS>
                <RESULT eventid="1076" points="600" reactiontime="+77" swimtime="00:00:27.56" resultid="3127" heatid="4284" lane="2" entrytime="00:00:27.00" />
                <RESULT eventid="1301" points="591" reactiontime="+77" swimtime="00:01:01.04" resultid="3128" heatid="4349" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" status="DNS" swimtime="00:00:00.00" resultid="3129" heatid="4356" lane="5" entrytime="00:03:00.00" />
                <RESULT eventid="1457" points="606" reactiontime="+73" swimtime="00:00:29.62" resultid="3130" heatid="4383" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1525" points="468" reactiontime="+81" swimtime="00:02:26.33" resultid="3131" heatid="4404" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:01:48.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="544" reactiontime="+74" swimtime="00:01:08.81" resultid="3132" heatid="4426" lane="0" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Babuchowski" birthdate="1984-06-08" gender="M" nation="POL" license="503605700040" athleteid="3117">
              <RESULTS>
                <RESULT eventid="1301" points="742" reactiontime="+69" swimtime="00:00:56.08" resultid="3118" heatid="4351" lane="4" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="795" reactiontime="+69" swimtime="00:00:26.06" resultid="3119" heatid="4384" lane="5" entrytime="00:00:26.00" />
                <RESULT eventid="1629" points="664" reactiontime="+72" swimtime="00:01:01.49" resultid="3120" heatid="4427" lane="7" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Adamska" birthdate="1984-09-25" gender="F" nation="POL" license="503605600036" athleteid="3109">
              <RESULTS>
                <RESULT eventid="1059" points="454" reactiontime="+61" swimtime="00:00:33.80" resultid="3110" heatid="4270" lane="5" entrytime="00:00:34.00" />
                <RESULT comment="Z3/G8" eventid="1094" status="DSQ" swimtime="00:00:00.00" resultid="3111" heatid="4287" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:03:27.28" />
                    <SPLIT distance="150" swimtime="00:02:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="341" reactiontime="+84" swimtime="00:00:40.96" resultid="3112" heatid="4315" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1284" points="421" reactiontime="+78" swimtime="00:01:17.53" resultid="3113" heatid="4339" lane="8" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="382" swimtime="00:00:37.86" resultid="3114" heatid="4374" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1508" points="323" reactiontime="+82" swimtime="00:03:03.56" resultid="3115" heatid="4396" lane="0">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="279" reactiontime="+76" swimtime="00:01:35.58" resultid="3116" heatid="4420" lane="2" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Frąckowiak" birthdate="1978-06-28" gender="M" nation="POL" license="503605700020" athleteid="3139">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3140" heatid="4282" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="3141" heatid="4348" lane="7" entrytime="00:01:05.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="3142" heatid="4381" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1697" status="DNS" swimtime="00:00:00.00" resultid="3143" heatid="4445" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Kurstak-Jagiełło" birthdate="1981-06-30" gender="F" nation="POL" license="503605600022" athleteid="3121">
              <RESULTS>
                <RESULT eventid="1059" points="679" reactiontime="+75" swimtime="00:00:30.08" resultid="3122" heatid="4266" lane="5" />
                <RESULT eventid="1284" points="649" reactiontime="+79" swimtime="00:01:07.04" resultid="3123" heatid="4335" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="577" reactiontime="+81" swimtime="00:02:35.27" resultid="3124" heatid="4395" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:56.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="432" reactiontime="+82" swimtime="00:00:42.94" resultid="3125" heatid="4438" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Woźniak" birthdate="1981-08-25" gender="M" nation="POL" license="503605700034" athleteid="3104">
              <RESULTS>
                <RESULT eventid="1267" status="DNS" swimtime="00:00:00.00" resultid="3105" heatid="4325" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="3106" heatid="4378" lane="9" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3107" heatid="4394" lane="6" entrytime="00:01:07.00" />
                <RESULT eventid="1663" status="DNS" swimtime="00:00:00.00" resultid="3108" heatid="4437" lane="2" entrytime="00:02:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1386" status="DNS" swimtime="00:00:00.00" resultid="3145" heatid="4493" lane="1" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3104" number="1" />
                    <RELAYPOSITION athleteid="3133" number="2" />
                    <RELAYPOSITION athleteid="3126" number="3" />
                    <RELAYPOSITION athleteid="3117" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="3146" heatid="4497" lane="3" entrytime="00:01:48.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3104" number="1" />
                    <RELAYPOSITION athleteid="3133" number="2" />
                    <RELAYPOSITION athleteid="3126" number="3" />
                    <RELAYPOSITION athleteid="3117" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1129" points="626" reactiontime="+85" swimtime="00:01:59.56" resultid="3144" heatid="4489" lane="3" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:01.74" />
                    <SPLIT distance="150" swimtime="00:01:31.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3109" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="3126" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="3121" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3133" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1714" points="577" reactiontime="+77" swimtime="00:02:16.04" resultid="3147" heatid="4499" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:16.78" />
                    <SPLIT distance="150" swimtime="00:01:46.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3109" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3133" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3126" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3121" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="04303" nation="POL" region="03" clubid="2202" name="Masters Avia Świdnik">
          <CONTACT city="Świdnik" email="tom.sitkowski@interia.pl" name="Sitkowski" phone="517487426" state="LUBEL" street="Modrzewiowa  10/13" zip="21-040" />
          <ATHLETES>
            <ATHLETE firstname="Cezary" lastname="Lipiński" birthdate="1972-04-11" gender="M" nation="POL" license="104303700002" swrid="5449345" athleteid="2208">
              <RESULTS>
                <RESULT eventid="1076" points="546" reactiontime="+70" swimtime="00:00:29.46" resultid="2209" heatid="4280" lane="5" entrytime="00:00:29.94" entrycourse="LCM" />
                <RESULT eventid="1163" points="510" reactiontime="+76" swimtime="00:11:09.54" resultid="2210" heatid="4305" lane="4" entrytime="00:11:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                    <SPLIT distance="150" swimtime="00:01:58.25" />
                    <SPLIT distance="200" swimtime="00:02:39.76" />
                    <SPLIT distance="250" swimtime="00:03:21.99" />
                    <SPLIT distance="300" swimtime="00:04:03.88" />
                    <SPLIT distance="350" swimtime="00:04:45.68" />
                    <SPLIT distance="400" swimtime="00:05:28.62" />
                    <SPLIT distance="450" swimtime="00:06:10.25" />
                    <SPLIT distance="500" swimtime="00:06:52.91" />
                    <SPLIT distance="550" swimtime="00:07:35.25" />
                    <SPLIT distance="600" swimtime="00:08:18.02" />
                    <SPLIT distance="650" swimtime="00:09:01.27" />
                    <SPLIT distance="700" swimtime="00:09:44.29" />
                    <SPLIT distance="750" swimtime="00:10:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="560" reactiontime="+77" swimtime="00:01:05.69" resultid="2211" heatid="4347" lane="6" entrytime="00:01:08.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="443" reactiontime="+81" swimtime="00:00:33.96" resultid="2212" heatid="4380" lane="4" entrytime="00:00:33.96" entrycourse="LCM" />
                <RESULT eventid="1525" points="496" reactiontime="+69" swimtime="00:02:29.81" resultid="2213" heatid="4403" lane="5" entrytime="00:02:30.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:12.08" />
                    <SPLIT distance="150" swimtime="00:01:51.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="534" reactiontime="+66" swimtime="00:05:15.53" resultid="2214" heatid="4459" lane="6" entrytime="00:05:22.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="150" swimtime="00:01:53.70" />
                    <SPLIT distance="200" swimtime="00:02:34.34" />
                    <SPLIT distance="300" swimtime="00:03:53.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Lipiec" birthdate="1973-03-19" gender="F" nation="POL" license="504303600010" athleteid="2203">
              <RESULTS>
                <RESULT eventid="1059" points="400" reactiontime="+95" swimtime="00:00:36.09" resultid="2204" heatid="4270" lane="1" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1284" points="365" reactiontime="+93" swimtime="00:01:20.32" resultid="2205" heatid="4339" lane="2" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="2206" heatid="4395" lane="0" />
                <RESULT eventid="1680" points="328" reactiontime="+92" swimtime="00:00:48.65" resultid="2207" heatid="4440" lane="6" entrytime="00:00:45.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Zielonka" birthdate="1986-05-26" gender="M" nation="POL" license="104303700006" swrid="4061691" athleteid="2224">
              <RESULTS>
                <RESULT eventid="1076" points="632" reactiontime="+71" swimtime="00:00:26.52" resultid="2225" heatid="4285" lane="3" entrytime="00:00:26.21" entrycourse="LCM" />
                <RESULT eventid="1163" points="518" reactiontime="+71" swimtime="00:10:20.61" resultid="2226" heatid="4303" lane="2" entrytime="00:09:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:08.15" />
                    <SPLIT distance="150" swimtime="00:01:45.10" />
                    <SPLIT distance="200" swimtime="00:02:22.69" />
                    <SPLIT distance="250" swimtime="00:03:01.09" />
                    <SPLIT distance="300" swimtime="00:03:40.22" />
                    <SPLIT distance="350" swimtime="00:04:19.49" />
                    <SPLIT distance="400" swimtime="00:04:59.10" />
                    <SPLIT distance="450" swimtime="00:05:38.86" />
                    <SPLIT distance="500" swimtime="00:06:19.09" />
                    <SPLIT distance="550" swimtime="00:06:59.64" />
                    <SPLIT distance="600" swimtime="00:07:40.22" />
                    <SPLIT distance="650" swimtime="00:08:20.95" />
                    <SPLIT distance="700" swimtime="00:09:01.39" />
                    <SPLIT distance="750" swimtime="00:09:41.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="695" reactiontime="+70" swimtime="00:00:57.33" resultid="2227" heatid="4351" lane="2" entrytime="00:00:57.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="601" reactiontime="+69" swimtime="00:00:28.60" resultid="2228" heatid="4384" lane="0" entrytime="00:00:27.88" entrycourse="LCM" />
                <RESULT eventid="1525" points="660" reactiontime="+69" swimtime="00:02:09.61" resultid="2229" heatid="4407" lane="1" entrytime="00:02:07.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:03.62" />
                    <SPLIT distance="150" swimtime="00:01:36.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" status="DNS" swimtime="00:00:00.00" resultid="2230" heatid="4426" lane="2" entrytime="00:01:04.82" entrycourse="LCM" />
                <RESULT eventid="1748" points="644" reactiontime="+76" swimtime="00:04:44.76" resultid="2231" heatid="4456" lane="7" entrytime="00:04:37.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:41.99" />
                    <SPLIT distance="200" swimtime="00:02:18.34" />
                    <SPLIT distance="250" swimtime="00:02:54.81" />
                    <SPLIT distance="300" swimtime="00:03:31.99" />
                    <SPLIT distance="350" swimtime="00:04:08.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Mazur" birthdate="1995-03-13" gender="M" nation="POL" license="104303700009" swrid="4195380" athleteid="2215">
              <RESULTS>
                <RESULT eventid="1076" points="678" reactiontime="+61" swimtime="00:00:25.38" resultid="2216" heatid="4286" lane="7" entrytime="00:00:25.24" entrycourse="LCM" />
                <RESULT eventid="1301" points="753" reactiontime="+70" swimtime="00:00:55.45" resultid="2217" heatid="4352" lane="8" entrytime="00:00:55.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="696" reactiontime="+67" swimtime="00:00:26.76" resultid="2218" heatid="4384" lane="8" entrytime="00:00:27.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Sitkowski" birthdate="1974-10-05" gender="M" nation="POL" license="504303700001" swrid="5439542" athleteid="2219">
              <RESULTS>
                <RESULT eventid="1076" points="586" reactiontime="+78" swimtime="00:00:28.14" resultid="2220" heatid="4281" lane="5" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1267" points="572" reactiontime="+70" swimtime="00:00:33.28" resultid="2221" heatid="4323" lane="3" entrytime="00:00:34.43" entrycourse="LCM" />
                <RESULT eventid="1491" points="529" reactiontime="+64" swimtime="00:01:14.34" resultid="2222" heatid="4393" lane="0" entrytime="00:01:17.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="431" reactiontime="+76" swimtime="00:02:54.22" resultid="2223" heatid="4435" lane="4" entrytime="00:02:53.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                    <SPLIT distance="150" swimtime="00:02:11.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1386" points="641" reactiontime="+80" swimtime="00:02:02.34" resultid="3828" heatid="4493" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:06.77" />
                    <SPLIT distance="150" swimtime="00:01:33.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2219" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2224" number="2" />
                    <RELAYPOSITION athleteid="2215" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2208" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="S1" eventid="1559" status="DSQ" swimtime="00:00:00.00" resultid="3829" heatid="4497" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.93" />
                    <SPLIT distance="100" swimtime="00:00:54.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2215" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2208" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2219" number="3" reactiontime="+55" status="DSQ" />
                    <RELAYPOSITION athleteid="2224" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" clubid="3495" name="Uks Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Płaneta" birthdate="1974-09-12" gender="M" nation="POL" license="500408700210" athleteid="3505">
              <RESULTS>
                <RESULT eventid="1076" points="428" reactiontime="+80" swimtime="00:00:31.25" resultid="3506" heatid="4279" lane="3" entrytime="00:00:31.30" />
                <RESULT eventid="1163" points="391" reactiontime="+86" swimtime="00:11:52.33" resultid="3507" heatid="4305" lane="8" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                    <SPLIT distance="100" swimtime="00:01:22.03" />
                    <SPLIT distance="150" swimtime="00:02:05.40" />
                    <SPLIT distance="200" swimtime="00:02:49.19" />
                    <SPLIT distance="250" swimtime="00:03:33.59" />
                    <SPLIT distance="300" swimtime="00:04:18.27" />
                    <SPLIT distance="350" swimtime="00:05:02.81" />
                    <SPLIT distance="400" swimtime="00:05:48.50" />
                    <SPLIT distance="450" swimtime="00:06:33.60" />
                    <SPLIT distance="500" swimtime="00:07:19.05" />
                    <SPLIT distance="550" swimtime="00:08:04.34" />
                    <SPLIT distance="600" swimtime="00:08:50.63" />
                    <SPLIT distance="650" swimtime="00:09:36.32" />
                    <SPLIT distance="700" swimtime="00:10:22.84" />
                    <SPLIT distance="750" swimtime="00:11:09.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="367" reactiontime="+101" swimtime="00:00:38.58" resultid="3508" heatid="4322" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1352" points="235" reactiontime="+84" swimtime="00:03:25.75" resultid="3509" heatid="4356" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                    <SPLIT distance="100" swimtime="00:01:36.02" />
                    <SPLIT distance="150" swimtime="00:02:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="317" reactiontime="+91" swimtime="00:01:28.18" resultid="3510" heatid="4392" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="377" reactiontime="+80" swimtime="00:02:43.05" resultid="3511" heatid="4403" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:20.52" />
                    <SPLIT distance="150" swimtime="00:02:03.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1663" points="324" reactiontime="+80" swimtime="00:03:11.47" resultid="3512" heatid="4434" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                    <SPLIT distance="100" swimtime="00:01:33.89" />
                    <SPLIT distance="150" swimtime="00:02:23.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" status="DNS" swimtime="00:00:00.00" resultid="3513" heatid="4459" lane="0" entrytime="00:05:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Janus" birthdate="1987-10-02" gender="F" nation="POL" athleteid="3496">
              <RESULTS>
                <RESULT eventid="1059" points="650" reactiontime="+75" swimtime="00:00:29.99" resultid="3497" heatid="4271" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1094" points="529" reactiontime="+91" swimtime="00:02:54.95" resultid="3498" heatid="4290" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:22.63" />
                    <SPLIT distance="150" swimtime="00:02:15.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="483" reactiontime="+76" swimtime="00:00:36.48" resultid="3499" heatid="4316" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1284" points="649" reactiontime="+85" swimtime="00:01:07.10" resultid="3500" heatid="4339" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="474" reactiontime="+84" swimtime="00:01:32.80" resultid="3501" heatid="4365" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="437" reactiontime="+77" swimtime="00:01:21.38" resultid="3502" heatid="4388" lane="1" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1646" points="439" reactiontime="+64" swimtime="00:03:01.83" resultid="3503" heatid="4431" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="493" reactiontime="+84" swimtime="00:00:41.35" resultid="3504" heatid="4440" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Ślęczka" birthdate="1974-10-23" gender="M" nation="POL" license="500408700205" athleteid="3514">
              <RESULTS>
                <RESULT eventid="1076" points="613" reactiontime="+84" swimtime="00:00:27.73" resultid="3515" heatid="4279" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1112" points="560" reactiontime="+84" swimtime="00:02:37.86" resultid="3516" heatid="4295" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:02:02.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="606" reactiontime="+73" swimtime="00:01:01.73" resultid="3517" heatid="4347" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="604" reactiontime="+76" swimtime="00:01:16.61" resultid="3518" heatid="4369" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="616" reactiontime="+77" swimtime="00:02:18.42" resultid="3519" heatid="4405" lane="3" entrytime="00:02:18.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="150" swimtime="00:01:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="565" reactiontime="+85" swimtime="00:00:35.35" resultid="3520" heatid="4446" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1748" points="539" reactiontime="+81" swimtime="00:05:08.59" resultid="3521" heatid="4458" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:13.90" />
                    <SPLIT distance="150" swimtime="00:01:53.43" />
                    <SPLIT distance="200" swimtime="00:02:33.72" />
                    <SPLIT distance="250" swimtime="00:03:14.25" />
                    <SPLIT distance="300" swimtime="00:03:54.78" />
                    <SPLIT distance="350" swimtime="00:04:32.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="2716" name="Pamirsti">
          <CONTACT name="Eimantas" />
          <ATHLETES>
            <ATHLETE firstname="Eimantas" lastname="Milius" birthdate="1996-07-22" gender="M" nation="LTU" athleteid="2717">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1112" points="919" reactiontime="+62" swimtime="00:02:07.13" resultid="2718" heatid="4297" lane="4" entrytime="00:02:05.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                    <SPLIT distance="100" swimtime="00:00:59.28" />
                    <SPLIT distance="150" swimtime="00:01:36.45" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1491" points="872" reactiontime="+61" swimtime="00:00:57.66" resultid="2719" heatid="4394" lane="4" entrytime="00:00:56.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1663" points="909" reactiontime="+57" swimtime="00:02:06.73" resultid="2720" heatid="4437" lane="4" entrytime="00:02:04.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:01.24" />
                    <SPLIT distance="150" swimtime="00:01:34.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gantas" lastname="Grigalionis" birthdate="2001-10-13" gender="M" nation="LTU" athleteid="2721">
              <RESULTS>
                <RESULT eventid="1112" reactiontime="+62" swimtime="00:02:12.31" resultid="2722" heatid="4297" lane="3" entrytime="00:02:12.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                    <SPLIT distance="100" swimtime="00:01:01.63" />
                    <SPLIT distance="150" swimtime="00:01:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" reactiontime="+57" swimtime="00:00:53.11" resultid="2723" heatid="4352" lane="5" entrytime="00:00:53.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" reactiontime="+62" swimtime="00:00:58.20" resultid="2724" heatid="4427" lane="3" entrytime="00:00:58.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3584" name="5 Styl Akademia Zajawki">
          <CONTACT city="Warszawa" name="Pawel Korzeniowski" phone="509249354" />
          <ATHLETES>
            <ATHLETE firstname="Pawel" lastname="Korzeniowski" birthdate="1985-07-09" gender="M" nation="POL" swrid="4042751" athleteid="3602">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1301" points="948" reactiontime="+75" swimtime="00:00:51.69" resultid="3603" heatid="4352" lane="4" entrytime="00:00:49.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters, Wynik lepszy od Rekordu Europy w kat. masters" eventid="1457" points="967" reactiontime="+68" swimtime="00:00:24.41" resultid="3604" heatid="4384" lane="4" entrytime="00:00:23.70" entrycourse="LCM" />
                <RESULT comment="Rekord Polski w kat.masters" eventid="1525" points="907" reactiontime="+74" swimtime="00:01:56.59" resultid="3605" heatid="4407" lane="4" entrytime="00:01:50.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.20" />
                    <SPLIT distance="100" swimtime="00:00:56.60" />
                    <SPLIT distance="150" swimtime="00:01:26.96" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1629" points="985" reactiontime="+71" swimtime="00:00:53.93" resultid="3606" heatid="4427" lane="4" entrytime="00:00:51.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Kozyra" birthdate="1959-12-25" gender="M" nation="POL" athleteid="3635">
              <RESULTS>
                <RESULT eventid="1076" points="364" reactiontime="+106" swimtime="00:00:35.35" resultid="3636" heatid="4277" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1112" points="248" reactiontime="+103" swimtime="00:03:45.92" resultid="3637" heatid="4292" lane="3" entrytime="00:04:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                    <SPLIT distance="100" swimtime="00:01:45.08" />
                    <SPLIT distance="150" swimtime="00:02:56.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="46" swimtime="00:01:17.32" resultid="3638" heatid="4378" lane="5" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Kulik" birthdate="1981-04-10" gender="M" nation="POL" athleteid="3622">
              <RESULTS>
                <RESULT eventid="1076" points="388" reactiontime="+79" swimtime="00:00:31.89" resultid="3623" heatid="4280" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1267" points="241" reactiontime="+92" swimtime="00:00:43.57" resultid="3624" heatid="4322" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1301" points="362" reactiontime="+81" swimtime="00:01:11.85" resultid="3625" heatid="4346" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="322" reactiontime="+80" swimtime="00:00:36.58" resultid="3626" heatid="4379" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1697" points="271" reactiontime="+76" swimtime="00:00:44.55" resultid="3627" heatid="4444" lane="6" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michal" lastname="Barnasiuk" birthdate="1992-02-04" gender="M" nation="POL" swrid="4273597" athleteid="3595">
              <RESULTS>
                <RESULT eventid="1112" points="613" reactiontime="+70" swimtime="00:02:23.84" resultid="3596" heatid="4296" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:50.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="671" reactiontime="+74" swimtime="00:02:37.71" resultid="3597" heatid="4334" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:14.58" />
                    <SPLIT distance="150" swimtime="00:01:56.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="626" reactiontime="+68" swimtime="00:01:11.61" resultid="3598" heatid="4371" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="598" reactiontime="+64" swimtime="00:05:09.64" resultid="3599" heatid="4414" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:09.47" />
                    <SPLIT distance="150" swimtime="00:01:52.74" />
                    <SPLIT distance="200" swimtime="00:02:35.37" />
                    <SPLIT distance="250" swimtime="00:03:16.81" />
                    <SPLIT distance="300" swimtime="00:03:59.59" />
                    <SPLIT distance="350" swimtime="00:04:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="554" reactiontime="+67" swimtime="00:01:05.32" resultid="3600" heatid="4425" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="629" reactiontime="+67" swimtime="00:00:32.62" resultid="3601" heatid="4448" lane="3" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Broniszewski" birthdate="1980-09-26" gender="M" nation="POL" athleteid="3585">
              <RESULTS>
                <RESULT eventid="1076" points="320" reactiontime="+84" swimtime="00:00:33.99" resultid="3586" heatid="4278" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1301" points="275" reactiontime="+87" swimtime="00:01:18.75" resultid="3587" heatid="4345" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="243" reactiontime="+88" swimtime="00:03:02.12" resultid="3588" heatid="4402" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="100" swimtime="00:01:23.70" />
                    <SPLIT distance="150" swimtime="00:02:12.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafal" lastname="Wziatek" birthdate="1988-01-14" gender="M" nation="POL" athleteid="3607">
              <RESULTS>
                <RESULT eventid="1197" points="248" reactiontime="+96" swimtime="00:24:34.32" resultid="3608" heatid="4309" lane="8" entrytime="00:20:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:19.61" />
                    <SPLIT distance="150" swimtime="00:02:04.99" />
                    <SPLIT distance="200" swimtime="00:02:51.82" />
                    <SPLIT distance="250" swimtime="00:03:40.01" />
                    <SPLIT distance="300" swimtime="00:04:28.53" />
                    <SPLIT distance="350" swimtime="00:05:18.01" />
                    <SPLIT distance="400" swimtime="00:06:07.54" />
                    <SPLIT distance="450" swimtime="00:06:57.31" />
                    <SPLIT distance="500" swimtime="00:07:46.96" />
                    <SPLIT distance="550" swimtime="00:08:36.92" />
                    <SPLIT distance="600" swimtime="00:09:26.32" />
                    <SPLIT distance="650" swimtime="00:10:16.35" />
                    <SPLIT distance="700" swimtime="00:11:06.67" />
                    <SPLIT distance="750" swimtime="00:11:57.04" />
                    <SPLIT distance="800" swimtime="00:12:47.91" />
                    <SPLIT distance="850" swimtime="00:13:38.58" />
                    <SPLIT distance="900" swimtime="00:14:28.98" />
                    <SPLIT distance="950" swimtime="00:15:19.43" />
                    <SPLIT distance="1000" swimtime="00:16:10.37" />
                    <SPLIT distance="1050" swimtime="00:17:01.50" />
                    <SPLIT distance="1100" swimtime="00:17:52.81" />
                    <SPLIT distance="1150" swimtime="00:18:44.28" />
                    <SPLIT distance="1200" swimtime="00:19:34.90" />
                    <SPLIT distance="1250" swimtime="00:20:24.97" />
                    <SPLIT distance="1300" swimtime="00:21:15.60" />
                    <SPLIT distance="1350" swimtime="00:22:05.76" />
                    <SPLIT distance="1400" swimtime="00:22:56.11" />
                    <SPLIT distance="1450" swimtime="00:23:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="334" reactiontime="+75" swimtime="00:01:11.76" resultid="3609" heatid="4345" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="302" reactiontime="+82" swimtime="00:02:43.33" resultid="3610" heatid="4402" lane="3" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:15.69" />
                    <SPLIT distance="150" swimtime="00:02:00.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Kantor" birthdate="1976-07-20" gender="F" nation="POL" athleteid="3628">
              <RESULTS>
                <RESULT eventid="1146" points="290" swimtime="00:13:53.41" resultid="3629" heatid="4301" lane="5" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                    <SPLIT distance="150" swimtime="00:02:17.81" />
                    <SPLIT distance="250" swimtime="00:05:37.47" />
                    <SPLIT distance="350" swimtime="00:07:18.34" />
                    <SPLIT distance="450" swimtime="00:08:59.63" />
                    <SPLIT distance="550" swimtime="00:10:40.24" />
                    <SPLIT distance="650" swimtime="00:12:20.63" />
                    <SPLIT distance="700" swimtime="00:13:07.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="266" reactiontime="+88" swimtime="00:00:48.22" resultid="3630" heatid="4314" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1284" points="336" reactiontime="+77" swimtime="00:01:22.58" resultid="3631" heatid="4338" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="394" reactiontime="+82" swimtime="00:02:57.41" resultid="3632" heatid="4397" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:25.96" />
                    <SPLIT distance="150" swimtime="00:02:13.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="329" reactiontime="+80" swimtime="00:00:48.62" resultid="3633" heatid="4440" lane="0" entrytime="00:00:50.00" />
                <RESULT eventid="1731" points="352" reactiontime="+44" swimtime="00:06:25.15" resultid="3634" heatid="4453" lane="8" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                    <SPLIT distance="150" swimtime="00:02:20.01" />
                    <SPLIT distance="200" swimtime="00:03:10.42" />
                    <SPLIT distance="250" swimtime="00:05:40.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Niedzwiadek" birthdate="1993-10-18" gender="M" nation="POL" athleteid="3589">
              <RESULTS>
                <RESULT eventid="1076" points="397" reactiontime="+75" swimtime="00:00:30.34" resultid="3590" heatid="4280" lane="1" entrytime="00:00:30.01" />
                <RESULT eventid="1163" points="487" reactiontime="+85" swimtime="00:10:41.58" resultid="3591" heatid="4303" lane="8" entrytime="00:10:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:13.54" />
                    <SPLIT distance="150" swimtime="00:01:53.44" />
                    <SPLIT distance="200" swimtime="00:02:32.90" />
                    <SPLIT distance="250" swimtime="00:03:13.44" />
                    <SPLIT distance="300" swimtime="00:03:53.69" />
                    <SPLIT distance="350" swimtime="00:04:34.81" />
                    <SPLIT distance="400" swimtime="00:05:15.69" />
                    <SPLIT distance="450" swimtime="00:05:56.14" />
                    <SPLIT distance="500" swimtime="00:06:36.69" />
                    <SPLIT distance="550" swimtime="00:07:17.41" />
                    <SPLIT distance="600" swimtime="00:07:58.25" />
                    <SPLIT distance="650" swimtime="00:08:39.32" />
                    <SPLIT distance="700" swimtime="00:09:20.87" />
                    <SPLIT distance="750" swimtime="00:10:01.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="450" reactiontime="+81" swimtime="00:01:05.84" resultid="3592" heatid="4347" lane="3" entrytime="00:01:07.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="469" reactiontime="+80" swimtime="00:02:22.52" resultid="3593" heatid="4404" lane="7" entrytime="00:02:27.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="150" swimtime="00:01:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1748" points="493" reactiontime="+86" swimtime="00:05:05.03" resultid="3594" heatid="4457" lane="8" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                    <SPLIT distance="150" swimtime="00:01:49.71" />
                    <SPLIT distance="200" swimtime="00:02:28.60" />
                    <SPLIT distance="250" swimtime="00:03:07.45" />
                    <SPLIT distance="300" swimtime="00:03:46.95" />
                    <SPLIT distance="350" swimtime="00:04:26.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michal" lastname="Butscher" birthdate="1975-01-18" gender="M" nation="POL" athleteid="3620">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3621" heatid="4278" lane="6" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Łatkowska" birthdate="1965-06-10" gender="F" nation="POL" athleteid="3611">
              <RESULTS>
                <RESULT eventid="1094" points="257" reactiontime="+84" swimtime="00:03:58.24" resultid="3612" heatid="4288" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.75" />
                    <SPLIT distance="100" swimtime="00:01:54.14" />
                    <SPLIT distance="150" swimtime="00:03:00.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="271" reactiontime="+86" swimtime="00:28:44.18" resultid="3613" heatid="4308" lane="6" entrytime="00:29:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.32" />
                    <SPLIT distance="100" swimtime="00:01:42.70" />
                    <SPLIT distance="150" swimtime="00:02:38.66" />
                    <SPLIT distance="200" swimtime="00:03:35.75" />
                    <SPLIT distance="250" swimtime="00:04:32.22" />
                    <SPLIT distance="300" swimtime="00:05:30.26" />
                    <SPLIT distance="350" swimtime="00:06:28.17" />
                    <SPLIT distance="400" swimtime="00:07:27.47" />
                    <SPLIT distance="450" swimtime="00:08:24.81" />
                    <SPLIT distance="500" swimtime="00:09:24.94" />
                    <SPLIT distance="550" swimtime="00:10:21.40" />
                    <SPLIT distance="600" swimtime="00:11:21.04" />
                    <SPLIT distance="650" swimtime="00:12:18.76" />
                    <SPLIT distance="700" swimtime="00:13:17.55" />
                    <SPLIT distance="750" swimtime="00:14:14.28" />
                    <SPLIT distance="800" swimtime="00:15:14.49" />
                    <SPLIT distance="850" swimtime="00:16:10.86" />
                    <SPLIT distance="900" swimtime="00:17:09.52" />
                    <SPLIT distance="950" swimtime="00:18:07.06" />
                    <SPLIT distance="1000" swimtime="00:19:06.67" />
                    <SPLIT distance="1050" swimtime="00:20:03.98" />
                    <SPLIT distance="1100" swimtime="00:21:03.81" />
                    <SPLIT distance="1150" swimtime="00:22:02.16" />
                    <SPLIT distance="1200" swimtime="00:23:01.05" />
                    <SPLIT distance="1250" swimtime="00:23:59.38" />
                    <SPLIT distance="1300" swimtime="00:24:58.12" />
                    <SPLIT distance="1350" swimtime="00:25:56.37" />
                    <SPLIT distance="1400" swimtime="00:26:54.45" />
                    <SPLIT distance="1450" swimtime="00:27:50.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="224" reactiontime="+86" swimtime="00:00:52.68" resultid="3614" heatid="4314" lane="7" entrytime="00:00:52.06" />
                <RESULT eventid="1284" points="271" reactiontime="+86" swimtime="00:01:35.89" resultid="3615" heatid="4337" lane="3" entrytime="00:01:37.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="172" swimtime="00:00:54.90" resultid="3616" heatid="4373" lane="7" entrytime="00:00:52.00" />
                <RESULT eventid="1508" points="279" reactiontime="+87" swimtime="00:03:28.66" resultid="3617" heatid="4396" lane="5" entrytime="00:03:29.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:41.74" />
                    <SPLIT distance="150" swimtime="00:02:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1680" points="270" reactiontime="+90" swimtime="00:00:55.60" resultid="3618" heatid="4439" lane="6" entrytime="00:01:00.00" />
                <RESULT eventid="1731" status="DNS" swimtime="00:00:00.00" resultid="3619" heatid="4454" lane="6" entrytime="00:07:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski w kat.masters" eventid="1559" points="564" reactiontime="+75" swimtime="00:01:52.35" resultid="4246" heatid="4496" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.85" />
                    <SPLIT distance="100" swimtime="00:00:51.02" />
                    <SPLIT distance="150" swimtime="00:01:20.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3602" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3595" number="2" />
                    <RELAYPOSITION athleteid="3589" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3622" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1386" points="506" reactiontime="+72" swimtime="00:02:08.40" resultid="4247" heatid="4491" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="100" swimtime="00:01:10.17" />
                    <SPLIT distance="150" swimtime="00:01:38.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3602" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="3585" number="2" />
                    <RELAYPOSITION athleteid="3595" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3589" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1714" points="434" reactiontime="+69" swimtime="00:02:29.53" resultid="4248" heatid="4498" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                    <SPLIT distance="150" swimtime="00:01:51.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3602" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3611" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="3595" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3628" number="4" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KS PIETRAS" nation="POL" clubid="2698" name="Klub Sportowy Pietraszyn">
          <CONTACT city="Pietraszyn" email="adip45@poczta.onet.pl" name="Piechula" phone="606114286" state="SLĄSK" street="Wesoła" zip="47-470" />
          <ATHLETES>
            <ATHLETE firstname="Adolf" lastname="Piechula" birthdate="1957-04-11" gender="M" nation="POL" swrid="4992724" athleteid="2699">
              <RESULTS>
                <RESULT eventid="1112" points="392" reactiontime="+98" swimtime="00:03:18.35" resultid="2700" heatid="4293" lane="2" entrytime="00:03:34.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                    <SPLIT distance="100" swimtime="00:01:33.13" />
                    <SPLIT distance="150" swimtime="00:02:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="411" reactiontime="+93" swimtime="00:03:37.34" resultid="2701" heatid="4331" lane="5" entrytime="00:03:45.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:40.30" />
                    <SPLIT distance="150" swimtime="00:02:39.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="324" reactiontime="+102" swimtime="00:03:43.36" resultid="2702" heatid="4356" lane="0" entrytime="00:03:35.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.39" />
                    <SPLIT distance="100" swimtime="00:01:45.24" />
                    <SPLIT distance="150" swimtime="00:02:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="473" reactiontime="+97" swimtime="00:01:35.98" resultid="2703" heatid="4368" lane="2" entrytime="00:01:38.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="364" reactiontime="+95" swimtime="00:07:18.72" resultid="2704" heatid="4416" lane="4" entrytime="00:06:54.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.88" />
                    <SPLIT distance="100" swimtime="00:01:45.89" />
                    <SPLIT distance="150" swimtime="00:02:42.86" />
                    <SPLIT distance="200" swimtime="00:03:39.22" />
                    <SPLIT distance="250" swimtime="00:04:39.10" />
                    <SPLIT distance="300" swimtime="00:05:39.29" />
                    <SPLIT distance="350" swimtime="00:06:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1629" points="288" reactiontime="+93" swimtime="00:01:39.73" resultid="2705" heatid="4424" lane="0" entrytime="00:01:36.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1697" points="466" reactiontime="+88" swimtime="00:00:42.94" resultid="2706" heatid="4444" lane="7" entrytime="00:00:46.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3739" name="SOPOT MASTERS">
          <ATHLETES>
            <ATHLETE firstname="DARIUSZ" lastname="GORBACZOW" birthdate="1958-01-01" gender="M" nation="POL" athleteid="3738" />
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SiKReT Gliwice" version="11.39204">
    <CONTACT name="Swimrankings" street="Weltpoststrasse 5" city="Bern" zip="3015" country="CH" phone="+41 99 999 99 99" fax="+41 99 999 99 99" email="sales@swimrankings.net" internet="http://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Gliwice" name="Mistrzostwa Polski w Pływaniu Masters" course="SCM" hostclub="SiKReT Gliwice" hostclub.url="http://www.sikret-plywanie.pl" nation="POL" organizer="Samorząd Miasta Gliwice, MZUK Gliwice, PZP,SLOZP,SiKReT Gliwice" result.url="http://www.megatiming.pl" timing="AUTOMATIC">
      <AGEDATE value="2015-11-15" type="YEAR" />
      <POOL name="Olimpijczyk Gliwice" lanemax="9" />
      <POINTTABLE pointtableid="3008" name="FINA Point Scoring" version="2015" />
      <CONTACT email="wisniowicz@interia.pl" name="Wojciech Wiśniowicz" phone="500193225" />
      <FEES>
        <FEE currency="PLN" type="ATHLETE" value="10000" />
        <FEE currency="PLN" type="LATEENTRY.INDIVIDUAL" value="15000" />
      </FEES>
      <SESSIONS>
        <SESSION date="2015-11-13" daytime="15:45" name="BLOK I" number="1" warmupfrom="14:30">
          <EVENTS>
            <EVENT eventid="1130" daytime="18:00" gender="X" number="5" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1182" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7523" />
                    <RANKING order="2" place="-1" resultid="7069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7903" />
                    <RANKING order="2" place="2" resultid="3623" />
                    <RANKING order="3" place="3" resultid="2554" />
                    <RANKING order="4" place="4" resultid="5952" />
                    <RANKING order="5" place="5" resultid="2869" />
                    <RANKING order="6" place="6" resultid="6297" />
                    <RANKING order="7" place="7" resultid="7065" />
                    <RANKING order="8" place="8" resultid="8599" />
                    <RANKING order="9" place="9" resultid="2752" />
                    <RANKING order="10" place="-1" resultid="4803" />
                    <RANKING order="11" place="-1" resultid="5742" />
                    <RANKING order="12" place="-1" resultid="5745" />
                    <RANKING order="13" place="-1" resultid="5828" />
                    <RANKING order="14" place="-1" resultid="7525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7393" />
                    <RANKING order="2" place="2" resultid="4293" />
                    <RANKING order="3" place="3" resultid="6306" />
                    <RANKING order="4" place="4" resultid="6912" />
                    <RANKING order="5" place="5" resultid="6296" />
                    <RANKING order="6" place="6" resultid="6033" />
                    <RANKING order="7" place="7" resultid="5827" />
                    <RANKING order="8" place="8" resultid="5599" />
                    <RANKING order="9" place="9" resultid="4929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7395" />
                    <RANKING order="2" place="2" resultid="3241" />
                    <RANKING order="3" place="3" resultid="6911" />
                    <RANKING order="4" place="4" resultid="2361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3625" />
                    <RANKING order="2" place="2" resultid="6416" />
                    <RANKING order="3" place="3" resultid="7397" />
                    <RANKING order="4" place="4" resultid="2357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6415" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8932" daytime="18:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8933" daytime="18:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8934" daytime="18:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8935" daytime="18:15" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="16:15" gender="M" number="2" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5873" />
                    <RANKING order="2" place="2" resultid="6903" />
                    <RANKING order="3" place="3" resultid="5631" />
                    <RANKING order="4" place="4" resultid="5540" />
                    <RANKING order="5" place="5" resultid="2857" />
                    <RANKING order="6" place="6" resultid="5531" />
                    <RANKING order="7" place="7" resultid="2118" />
                    <RANKING order="8" place="8" resultid="3253" />
                    <RANKING order="9" place="-1" resultid="4148" />
                    <RANKING order="10" place="-1" resultid="6182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5974" />
                    <RANKING order="2" place="2" resultid="2091" />
                    <RANKING order="3" place="3" resultid="2137" />
                    <RANKING order="4" place="4" resultid="5103" />
                    <RANKING order="5" place="5" resultid="3613" />
                    <RANKING order="6" place="6" resultid="4835" />
                    <RANKING order="7" place="7" resultid="4716" />
                    <RANKING order="8" place="8" resultid="4709" />
                    <RANKING order="9" place="9" resultid="3492" />
                    <RANKING order="10" place="10" resultid="4704" />
                    <RANKING order="11" place="11" resultid="2789" />
                    <RANKING order="12" place="12" resultid="7038" />
                    <RANKING order="13" place="13" resultid="2070" />
                    <RANKING order="14" place="14" resultid="7141" />
                    <RANKING order="15" place="15" resultid="1921" />
                    <RANKING order="16" place="16" resultid="1932" />
                    <RANKING order="17" place="17" resultid="4616" />
                    <RANKING order="18" place="-1" resultid="5071" />
                    <RANKING order="19" place="-1" resultid="5925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3711" />
                    <RANKING order="2" place="2" resultid="7188" />
                    <RANKING order="3" place="3" resultid="2085" />
                    <RANKING order="4" place="4" resultid="7237" />
                    <RANKING order="5" place="5" resultid="7172" />
                    <RANKING order="6" place="6" resultid="5116" />
                    <RANKING order="7" place="7" resultid="2472" />
                    <RANKING order="8" place="8" resultid="7181" />
                    <RANKING order="9" place="9" resultid="6888" />
                    <RANKING order="10" place="10" resultid="4713" />
                    <RANKING order="11" place="11" resultid="2844" />
                    <RANKING order="12" place="12" resultid="5896" />
                    <RANKING order="13" place="13" resultid="5920" />
                    <RANKING order="14" place="14" resultid="3717" />
                    <RANKING order="15" place="15" resultid="5585" />
                    <RANKING order="16" place="16" resultid="4763" />
                    <RANKING order="17" place="17" resultid="4951" />
                    <RANKING order="18" place="18" resultid="2745" />
                    <RANKING order="19" place="19" resultid="4200" />
                    <RANKING order="20" place="20" resultid="3209" />
                    <RANKING order="21" place="21" resultid="2539" />
                    <RANKING order="22" place="22" resultid="7059" />
                    <RANKING order="23" place="23" resultid="4884" />
                    <RANKING order="24" place="24" resultid="6158" />
                    <RANKING order="25" place="25" resultid="2725" />
                    <RANKING order="26" place="26" resultid="2548" />
                    <RANKING order="27" place="-1" resultid="2142" />
                    <RANKING order="28" place="-1" resultid="3370" />
                    <RANKING order="29" place="-1" resultid="4778" />
                    <RANKING order="30" place="-1" resultid="5979" />
                    <RANKING order="31" place="-1" resultid="7356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1771" />
                    <RANKING order="2" place="2" resultid="5942" />
                    <RANKING order="3" place="3" resultid="3598" />
                    <RANKING order="4" place="4" resultid="2804" />
                    <RANKING order="5" place="5" resultid="5914" />
                    <RANKING order="6" place="6" resultid="3699" />
                    <RANKING order="7" place="6" resultid="6258" />
                    <RANKING order="8" place="8" resultid="3756" />
                    <RANKING order="9" place="9" resultid="3687" />
                    <RANKING order="10" place="10" resultid="3976" />
                    <RANKING order="11" place="11" resultid="6273" />
                    <RANKING order="12" place="12" resultid="4940" />
                    <RANKING order="13" place="13" resultid="3729" />
                    <RANKING order="14" place="14" resultid="3695" />
                    <RANKING order="15" place="15" resultid="3741" />
                    <RANKING order="16" place="16" resultid="4863" />
                    <RANKING order="17" place="17" resultid="3877" />
                    <RANKING order="18" place="18" resultid="3725" />
                    <RANKING order="19" place="19" resultid="3736" />
                    <RANKING order="20" place="20" resultid="3940" />
                    <RANKING order="21" place="21" resultid="7298" />
                    <RANKING order="22" place="22" resultid="2395" />
                    <RANKING order="23" place="23" resultid="2100" />
                    <RANKING order="24" place="24" resultid="4770" />
                    <RANKING order="25" place="25" resultid="1924" />
                    <RANKING order="26" place="-1" resultid="3705" />
                    <RANKING order="27" place="-1" resultid="4009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2700" />
                    <RANKING order="2" place="2" resultid="6220" />
                    <RANKING order="3" place="3" resultid="2667" />
                    <RANKING order="4" place="4" resultid="4280" />
                    <RANKING order="5" place="5" resultid="4687" />
                    <RANKING order="6" place="6" resultid="3215" />
                    <RANKING order="7" place="7" resultid="4230" />
                    <RANKING order="8" place="8" resultid="3935" />
                    <RANKING order="9" place="9" resultid="3554" />
                    <RANKING order="10" place="10" resultid="5999" />
                    <RANKING order="11" place="11" resultid="4275" />
                    <RANKING order="12" place="12" resultid="3902" />
                    <RANKING order="13" place="13" resultid="2425" />
                    <RANKING order="14" place="14" resultid="7248" />
                    <RANKING order="15" place="15" resultid="1893" />
                    <RANKING order="16" place="16" resultid="5963" />
                    <RANKING order="17" place="17" resultid="7047" />
                    <RANKING order="18" place="18" resultid="4238" />
                    <RANKING order="19" place="19" resultid="4758" />
                    <RANKING order="20" place="20" resultid="2422" />
                    <RANKING order="21" place="21" resultid="2158" />
                    <RANKING order="22" place="22" resultid="2811" />
                    <RANKING order="23" place="23" resultid="6229" />
                    <RANKING order="24" place="24" resultid="3225" />
                    <RANKING order="25" place="25" resultid="3237" />
                    <RANKING order="26" place="26" resultid="2042" />
                    <RANKING order="27" place="-1" resultid="2263" />
                    <RANKING order="28" place="-1" resultid="4269" />
                    <RANKING order="29" place="-1" resultid="4784" />
                    <RANKING order="30" place="-1" resultid="4946" />
                    <RANKING order="31" place="-1" resultid="5711" />
                    <RANKING order="32" place="-1" resultid="5729" />
                    <RANKING order="33" place="-1" resultid="5799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3915" />
                    <RANKING order="2" place="2" resultid="4827" />
                    <RANKING order="3" place="3" resultid="4819" />
                    <RANKING order="4" place="4" resultid="4071" />
                    <RANKING order="5" place="5" resultid="3177" />
                    <RANKING order="6" place="6" resultid="2795" />
                    <RANKING order="7" place="7" resultid="6132" />
                    <RANKING order="8" place="8" resultid="2052" />
                    <RANKING order="9" place="9" resultid="5815" />
                    <RANKING order="10" place="10" resultid="2944" />
                    <RANKING order="11" place="11" resultid="2007" />
                    <RANKING order="12" place="12" resultid="4925" />
                    <RANKING order="13" place="13" resultid="6289" />
                    <RANKING order="14" place="14" resultid="2960" />
                    <RANKING order="15" place="15" resultid="3895" />
                    <RANKING order="16" place="16" resultid="2414" />
                    <RANKING order="17" place="17" resultid="7353" />
                    <RANKING order="18" place="18" resultid="5546" />
                    <RANKING order="19" place="19" resultid="9195" />
                    <RANKING order="20" place="-1" resultid="6333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3884" />
                    <RANKING order="2" place="2" resultid="6898" />
                    <RANKING order="3" place="3" resultid="7105" />
                    <RANKING order="4" place="4" resultid="2044" />
                    <RANKING order="5" place="5" resultid="6150" />
                    <RANKING order="6" place="6" resultid="7303" />
                    <RANKING order="7" place="7" resultid="3390" />
                    <RANKING order="8" place="8" resultid="3231" />
                    <RANKING order="9" place="9" resultid="3579" />
                    <RANKING order="10" place="10" resultid="5678" />
                    <RANKING order="11" place="-1" resultid="3584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3790" />
                    <RANKING order="2" place="2" resultid="5097" />
                    <RANKING order="3" place="3" resultid="6266" />
                    <RANKING order="4" place="4" resultid="5883" />
                    <RANKING order="5" place="5" resultid="2691" />
                    <RANKING order="6" place="6" resultid="6375" />
                    <RANKING order="7" place="7" resultid="2563" />
                    <RANKING order="8" place="8" resultid="7112" />
                    <RANKING order="9" place="9" resultid="4304" />
                    <RANKING order="10" place="10" resultid="4613" />
                    <RANKING order="11" place="11" resultid="7341" />
                    <RANKING order="12" place="12" resultid="2604" />
                    <RANKING order="13" place="13" resultid="3218" />
                    <RANKING order="14" place="14" resultid="7325" />
                    <RANKING order="15" place="15" resultid="2321" />
                    <RANKING order="16" place="16" resultid="3870" />
                    <RANKING order="17" place="17" resultid="2570" />
                    <RANKING order="18" place="18" resultid="2299" />
                    <RANKING order="19" place="19" resultid="7387" />
                    <RANKING order="20" place="-1" resultid="3500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2182" />
                    <RANKING order="2" place="2" resultid="1888" />
                    <RANKING order="3" place="3" resultid="3143" />
                    <RANKING order="4" place="4" resultid="2632" />
                    <RANKING order="5" place="5" resultid="3009" />
                    <RANKING order="6" place="6" resultid="5706" />
                    <RANKING order="7" place="7" resultid="5854" />
                    <RANKING order="8" place="8" resultid="2060" />
                    <RANKING order="9" place="9" resultid="1905" />
                    <RANKING order="10" place="10" resultid="4652" />
                    <RANKING order="11" place="11" resultid="2285" />
                    <RANKING order="12" place="12" resultid="2818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3509" />
                    <RANKING order="2" place="2" resultid="1912" />
                    <RANKING order="3" place="3" resultid="7280" />
                    <RANKING order="4" place="4" resultid="6398" />
                    <RANKING order="5" place="5" resultid="2622" />
                    <RANKING order="6" place="6" resultid="6359" />
                    <RANKING order="7" place="7" resultid="2306" />
                    <RANKING order="8" place="8" resultid="2272" />
                    <RANKING order="9" place="-1" resultid="3815" />
                    <RANKING order="10" place="-1" resultid="2478" />
                    <RANKING order="11" place="-1" resultid="3487" />
                    <RANKING order="12" place="-1" resultid="6932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1784" />
                    <RANKING order="2" place="2" resultid="3840" />
                    <RANKING order="3" place="3" resultid="4644" />
                    <RANKING order="4" place="4" resultid="3361" />
                    <RANKING order="5" place="5" resultid="2952" />
                    <RANKING order="6" place="6" resultid="1879" />
                    <RANKING order="7" place="7" resultid="3325" />
                    <RANKING order="8" place="8" resultid="1990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7097" />
                    <RANKING order="2" place="2" resultid="2992" />
                    <RANKING order="3" place="3" resultid="2494" />
                    <RANKING order="4" place="4" resultid="7334" />
                    <RANKING order="5" place="5" resultid="5847" />
                    <RANKING order="6" place="6" resultid="1956" />
                    <RANKING order="7" place="7" resultid="3824" />
                    <RANKING order="8" place="8" resultid="2499" />
                    <RANKING order="9" place="9" resultid="1983" />
                    <RANKING order="10" place="10" resultid="2293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5734" />
                    <RANKING order="2" place="2" resultid="5753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8894" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8895" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8896" daytime="16:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8897" daytime="16:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8898" daytime="16:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8899" daytime="16:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8900" daytime="16:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8901" daytime="16:30" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8902" daytime="16:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8903" daytime="16:30" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="8904" daytime="16:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="8905" daytime="16:35" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="8906" daytime="16:35" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="8907" daytime="16:35" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="8908" daytime="16:40" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="8909" daytime="16:40" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="8910" daytime="16:40" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="8911" daytime="16:40" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="8912" daytime="16:45" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="8913" daytime="16:45" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="8914" daytime="16:45" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="8915" daytime="16:45" number="22" order="22" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="17:15" gender="M" number="4" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1114" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2257" />
                    <RANKING order="2" place="2" resultid="6904" />
                    <RANKING order="3" place="3" resultid="5632" />
                    <RANKING order="4" place="4" resultid="1801" />
                    <RANKING order="5" place="5" resultid="5077" />
                    <RANKING order="6" place="6" resultid="3356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3593" />
                    <RANKING order="2" place="2" resultid="2092" />
                    <RANKING order="3" place="3" resultid="5104" />
                    <RANKING order="4" place="4" resultid="4877" />
                    <RANKING order="5" place="5" resultid="2850" />
                    <RANKING order="6" place="6" resultid="4215" />
                    <RANKING order="7" place="7" resultid="3167" />
                    <RANKING order="8" place="8" resultid="3493" />
                    <RANKING order="9" place="9" resultid="3849" />
                    <RANKING order="10" place="10" resultid="7142" />
                    <RANKING order="11" place="11" resultid="7024" />
                    <RANKING order="12" place="12" resultid="7039" />
                    <RANKING order="13" place="13" resultid="2128" />
                    <RANKING order="14" place="-1" resultid="2071" />
                    <RANKING order="15" place="-1" resultid="4169" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7091" />
                    <RANKING order="2" place="2" resultid="7189" />
                    <RANKING order="3" place="3" resultid="7173" />
                    <RANKING order="4" place="4" resultid="5897" />
                    <RANKING order="5" place="5" resultid="3856" />
                    <RANKING order="6" place="6" resultid="3718" />
                    <RANKING order="7" place="7" resultid="2540" />
                    <RANKING order="8" place="8" resultid="4885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6879" />
                    <RANKING order="2" place="2" resultid="6259" />
                    <RANKING order="3" place="3" resultid="3910" />
                    <RANKING order="4" place="4" resultid="2153" />
                    <RANKING order="5" place="5" resultid="4894" />
                    <RANKING order="6" place="6" resultid="2658" />
                    <RANKING order="7" place="7" resultid="2650" />
                    <RANKING order="8" place="8" resultid="7381" />
                    <RANKING order="9" place="9" resultid="3730" />
                    <RANKING order="10" place="10" resultid="3941" />
                    <RANKING order="11" place="11" resultid="2684" />
                    <RANKING order="12" place="12" resultid="5808" />
                    <RANKING order="13" place="-1" resultid="2396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2701" />
                    <RANKING order="2" place="2" resultid="4955" />
                    <RANKING order="3" place="3" resultid="6221" />
                    <RANKING order="4" place="4" resultid="2668" />
                    <RANKING order="5" place="5" resultid="4281" />
                    <RANKING order="6" place="6" resultid="4231" />
                    <RANKING order="7" place="7" resultid="3781" />
                    <RANKING order="8" place="8" resultid="2264" />
                    <RANKING order="9" place="9" resultid="3555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3916" />
                    <RANKING order="2" place="2" resultid="3833" />
                    <RANKING order="3" place="3" resultid="4820" />
                    <RANKING order="4" place="4" resultid="3178" />
                    <RANKING order="5" place="5" resultid="4076" />
                    <RANKING order="6" place="6" resultid="4621" />
                    <RANKING order="7" place="7" resultid="2460" />
                    <RANKING order="8" place="8" resultid="2008" />
                    <RANKING order="9" place="-1" resultid="3351" />
                    <RANKING order="10" place="-1" resultid="4828" />
                    <RANKING order="11" place="-1" resultid="5816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2045" />
                    <RANKING order="2" place="2" resultid="3391" />
                    <RANKING order="3" place="3" resultid="4806" />
                    <RANKING order="4" place="4" resultid="6861" />
                    <RANKING order="5" place="5" resultid="6236" />
                    <RANKING order="6" place="6" resultid="5929" />
                    <RANKING order="7" place="7" resultid="6831" />
                    <RANKING order="8" place="8" resultid="3585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2692" />
                    <RANKING order="2" place="2" resultid="3501" />
                    <RANKING order="3" place="3" resultid="5862" />
                    <RANKING order="4" place="4" resultid="2405" />
                    <RANKING order="5" place="5" resultid="4666" />
                    <RANKING order="6" place="6" resultid="3477" />
                    <RANKING order="7" place="7" resultid="2584" />
                    <RANKING order="8" place="8" resultid="7326" />
                    <RANKING order="9" place="-1" resultid="3153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3964" />
                    <RANKING order="2" place="2" resultid="2183" />
                    <RANKING order="3" place="3" resultid="2937" />
                    <RANKING order="4" place="4" resultid="4658" />
                    <RANKING order="5" place="5" resultid="1965" />
                    <RANKING order="6" place="6" resultid="1906" />
                    <RANKING order="7" place="7" resultid="2576" />
                    <RANKING order="8" place="8" resultid="1974" />
                    <RANKING order="9" place="9" resultid="3144" />
                    <RANKING order="10" place="-1" resultid="2524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2676" />
                    <RANKING order="2" place="2" resultid="1927" />
                    <RANKING order="3" place="3" resultid="3510" />
                    <RANKING order="4" place="4" resultid="3020" />
                    <RANKING order="5" place="5" resultid="7281" />
                    <RANKING order="6" place="6" resultid="2485" />
                    <RANKING order="7" place="-1" resultid="2273" />
                    <RANKING order="8" place="-1" resultid="5697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1785" />
                    <RANKING order="2" place="2" resultid="4645" />
                    <RANKING order="3" place="3" resultid="1880" />
                    <RANKING order="4" place="-1" resultid="2313" />
                    <RANKING order="5" place="-1" resultid="7261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6381" />
                    <RANKING order="2" place="2" resultid="2993" />
                    <RANKING order="3" place="3" resultid="1957" />
                    <RANKING order="4" place="4" resultid="3825" />
                    <RANKING order="5" place="-1" resultid="7098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1127" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1129" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8921" daytime="17:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8922" daytime="17:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8923" daytime="17:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8924" daytime="17:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8925" daytime="17:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8926" daytime="17:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8927" daytime="17:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8928" daytime="17:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8929" daytime="17:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8930" daytime="17:55" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="8931" daytime="18:00" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="19:20" gender="M" number="7" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1166" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1802" />
                    <RANKING order="2" place="-1" resultid="4149" />
                    <RANKING order="3" place="-1" resultid="5078" />
                    <RANKING order="4" place="-1" resultid="2258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4157" />
                    <RANKING order="2" place="2" resultid="3168" />
                    <RANKING order="3" place="3" resultid="2200" />
                    <RANKING order="4" place="4" resultid="2129" />
                    <RANKING order="5" place="-1" resultid="2790" />
                    <RANKING order="6" place="-1" resultid="4908" />
                    <RANKING order="7" place="-1" resultid="4164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3857" />
                    <RANKING order="2" place="2" resultid="2746" />
                    <RANKING order="3" place="-1" resultid="7357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6880" />
                    <RANKING order="2" place="2" resultid="3878" />
                    <RANKING order="3" place="3" resultid="3977" />
                    <RANKING order="4" place="4" resultid="5718" />
                    <RANKING order="5" place="5" resultid="3742" />
                    <RANKING order="6" place="6" resultid="3911" />
                    <RANKING order="7" place="7" resultid="2039" />
                    <RANKING order="8" place="8" resultid="6274" />
                    <RANKING order="9" place="9" resultid="2106" />
                    <RANKING order="10" place="10" resultid="5809" />
                    <RANKING order="11" place="-1" resultid="2659" />
                    <RANKING order="12" place="-1" resultid="3688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3782" />
                    <RANKING order="2" place="2" resultid="7317" />
                    <RANKING order="3" place="3" resultid="3666" />
                    <RANKING order="4" place="4" resultid="2208" />
                    <RANKING order="5" place="5" resultid="7249" />
                    <RANKING order="6" place="6" resultid="4977" />
                    <RANKING order="7" place="7" resultid="6005" />
                    <RANKING order="8" place="8" resultid="1894" />
                    <RANKING order="9" place="9" resultid="4239" />
                    <RANKING order="10" place="10" resultid="2159" />
                    <RANKING order="11" place="-1" resultid="3903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2053" />
                    <RANKING order="2" place="2" resultid="2796" />
                    <RANKING order="3" place="3" resultid="6855" />
                    <RANKING order="4" place="4" resultid="7354" />
                    <RANKING order="5" place="5" resultid="9194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8880" />
                    <RANKING order="2" place="2" resultid="5930" />
                    <RANKING order="3" place="3" resultid="3341" />
                    <RANKING order="4" place="4" resultid="6849" />
                    <RANKING order="5" place="-1" resultid="3383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6267" />
                    <RANKING order="2" place="2" resultid="2406" />
                    <RANKING order="3" place="3" resultid="4305" />
                    <RANKING order="4" place="4" resultid="3478" />
                    <RANKING order="5" place="5" resultid="2605" />
                    <RANKING order="6" place="6" resultid="7342" />
                    <RANKING order="7" place="7" resultid="3871" />
                    <RANKING order="8" place="8" resultid="2611" />
                    <RANKING order="9" place="9" resultid="3989" />
                    <RANKING order="10" place="10" resultid="2322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5645" />
                    <RANKING order="2" place="2" resultid="3010" />
                    <RANKING order="3" place="3" resultid="1966" />
                    <RANKING order="4" place="4" resultid="2061" />
                    <RANKING order="5" place="5" resultid="2385" />
                    <RANKING order="6" place="6" resultid="1975" />
                    <RANKING order="7" place="7" resultid="2589" />
                    <RANKING order="8" place="-1" resultid="2819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3816" />
                    <RANKING order="2" place="2" resultid="1913" />
                    <RANKING order="3" place="3" resultid="1944" />
                    <RANKING order="4" place="4" resultid="2623" />
                    <RANKING order="5" place="5" resultid="6933" />
                    <RANKING order="6" place="6" resultid="3609" />
                    <RANKING order="7" place="-1" resultid="2486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3362" />
                    <RANKING order="2" place="2" resultid="3841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7225" />
                    <RANKING order="2" place="2" resultid="7335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1180" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1181" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8940" daytime="19:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8941" daytime="20:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8942" daytime="20:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8943" daytime="21:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8944" daytime="21:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8945" daytime="22:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8946" daytime="22:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8947" daytime="22:50" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="16:50" gender="F" number="3" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2781" />
                    <RANKING order="2" place="2" resultid="5624" />
                    <RANKING order="3" place="3" resultid="7017" />
                    <RANKING order="4" place="4" resultid="1811" />
                    <RANKING order="5" place="5" resultid="7031" />
                    <RANKING order="6" place="-1" resultid="2836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3345" />
                    <RANKING order="2" place="2" resultid="4842" />
                    <RANKING order="3" place="3" resultid="6242" />
                    <RANKING order="4" place="4" resultid="7010" />
                    <RANKING order="5" place="5" resultid="2507" />
                    <RANKING order="6" place="6" resultid="5618" />
                    <RANKING order="7" place="7" resultid="5778" />
                    <RANKING order="8" place="-1" resultid="7003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3984" />
                    <RANKING order="2" place="2" resultid="2761" />
                    <RANKING order="3" place="3" resultid="2516" />
                    <RANKING order="4" place="4" resultid="4698" />
                    <RANKING order="5" place="5" resultid="6186" />
                    <RANKING order="6" place="6" resultid="4970" />
                    <RANKING order="7" place="7" resultid="5553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4254" />
                    <RANKING order="2" place="2" resultid="6250" />
                    <RANKING order="3" place="3" resultid="4752" />
                    <RANKING order="4" place="4" resultid="2734" />
                    <RANKING order="5" place="5" resultid="5560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3540" />
                    <RANKING order="2" place="2" resultid="4903" />
                    <RANKING order="3" place="3" resultid="6010" />
                    <RANKING order="4" place="4" resultid="2443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7347" />
                    <RANKING order="2" place="2" resultid="2642" />
                    <RANKING order="3" place="3" resultid="6281" />
                    <RANKING order="4" place="4" resultid="2452" />
                    <RANKING order="5" place="5" resultid="5592" />
                    <RANKING order="6" place="-1" resultid="5668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="1104" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3465" />
                    <RANKING order="2" place="2" resultid="5792" />
                    <RANKING order="3" place="3" resultid="2240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3001" />
                    <RANKING order="2" place="2" resultid="3617" />
                    <RANKING order="3" place="3" resultid="3029" />
                    <RANKING order="4" place="4" resultid="1818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5568" />
                    <RANKING order="2" place="2" resultid="7290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1108" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1110" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1111" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1112" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8916" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8917" daytime="17:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8918" daytime="17:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8919" daytime="17:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8920" daytime="17:15" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1062" daytime="16:00" gender="F" number="1" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5623" />
                    <RANKING order="2" place="2" resultid="7133" />
                    <RANKING order="3" place="3" resultid="2780" />
                    <RANKING order="4" place="4" resultid="7052" />
                    <RANKING order="5" place="5" resultid="5762" />
                    <RANKING order="6" place="6" resultid="4183" />
                    <RANKING order="7" place="7" resultid="1810" />
                    <RANKING order="8" place="8" resultid="7016" />
                    <RANKING order="9" place="9" resultid="7030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4722" />
                    <RANKING order="2" place="2" resultid="4870" />
                    <RANKING order="3" place="3" resultid="7127" />
                    <RANKING order="4" place="4" resultid="1938" />
                    <RANKING order="5" place="5" resultid="5909" />
                    <RANKING order="6" place="6" resultid="3376" />
                    <RANKING order="7" place="7" resultid="5968" />
                    <RANKING order="8" place="8" resultid="2078" />
                    <RANKING order="9" place="9" resultid="7165" />
                    <RANKING order="10" place="10" resultid="6138" />
                    <RANKING order="11" place="11" resultid="6029" />
                    <RANKING order="12" place="-1" resultid="3572" />
                    <RANKING order="13" place="-1" resultid="7157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3983" />
                    <RANKING order="2" place="2" resultid="3440" />
                    <RANKING order="3" place="3" resultid="4697" />
                    <RANKING order="4" place="4" resultid="4962" />
                    <RANKING order="5" place="5" resultid="3865" />
                    <RANKING order="6" place="6" resultid="5904" />
                    <RANKING order="7" place="7" resultid="4812" />
                    <RANKING order="8" place="8" resultid="3681" />
                    <RANKING order="9" place="9" resultid="3748" />
                    <RANKING order="10" place="-1" resultid="4015" />
                    <RANKING order="11" place="-1" resultid="4790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2531" />
                    <RANKING order="2" place="2" resultid="6194" />
                    <RANKING order="3" place="3" resultid="4751" />
                    <RANKING order="4" place="4" resultid="4262" />
                    <RANKING order="5" place="5" resultid="6249" />
                    <RANKING order="6" place="6" resultid="2733" />
                    <RANKING order="7" place="7" resultid="4253" />
                    <RANKING order="8" place="8" resultid="4850" />
                    <RANKING order="9" place="9" resultid="3202" />
                    <RANKING order="10" place="10" resultid="4900" />
                    <RANKING order="11" place="-1" resultid="6294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3547" />
                    <RANKING order="2" place="2" resultid="3923" />
                    <RANKING order="3" place="3" resultid="3140" />
                    <RANKING order="4" place="4" resultid="7254" />
                    <RANKING order="5" place="5" resultid="6017" />
                    <RANKING order="6" place="-1" resultid="4797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7230" />
                    <RANKING order="2" place="2" resultid="7243" />
                    <RANKING order="3" place="3" resultid="5614" />
                    <RANKING order="4" place="4" resultid="5802" />
                    <RANKING order="5" place="5" resultid="2641" />
                    <RANKING order="6" place="6" resultid="2451" />
                    <RANKING order="7" place="7" resultid="5591" />
                    <RANKING order="8" place="8" resultid="5868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3521" />
                    <RANKING order="2" place="2" resultid="3526" />
                    <RANKING order="3" place="3" resultid="6867" />
                    <RANKING order="4" place="4" resultid="3333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7271" />
                    <RANKING order="2" place="2" resultid="6838" />
                    <RANKING order="3" place="3" resultid="3193" />
                    <RANKING order="4" place="4" resultid="5791" />
                    <RANKING order="5" place="5" resultid="3185" />
                    <RANKING order="6" place="6" resultid="4638" />
                    <RANKING order="7" place="7" resultid="2330" />
                    <RANKING order="8" place="8" resultid="5086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3616" />
                    <RANKING order="2" place="2" resultid="3028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5608" />
                    <RANKING order="2" place="2" resultid="4630" />
                    <RANKING order="3" place="3" resultid="6402" />
                    <RANKING order="4" place="4" resultid="3929" />
                    <RANKING order="5" place="5" resultid="5663" />
                    <RANKING order="6" place="6" resultid="4004" />
                    <RANKING order="7" place="7" resultid="7289" />
                    <RANKING order="8" place="8" resultid="1998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1077" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1078" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1063" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8885" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8886" daytime="16:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8887" daytime="16:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8888" daytime="16:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8889" daytime="16:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8890" daytime="16:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8891" daytime="16:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8892" daytime="16:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8893" daytime="16:15" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1147" daytime="18:15" gender="F" number="6" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3377" />
                    <RANKING order="2" place="2" resultid="2231" />
                    <RANKING order="3" place="3" resultid="4843" />
                    <RANKING order="4" place="4" resultid="2508" />
                    <RANKING order="5" place="5" resultid="5619" />
                    <RANKING order="6" place="6" resultid="5785" />
                    <RANKING order="7" place="-1" resultid="5655" />
                    <RANKING order="8" place="-1" resultid="6139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6187" />
                    <RANKING order="2" place="2" resultid="6216" />
                    <RANKING order="3" place="3" resultid="6202" />
                    <RANKING order="4" place="4" resultid="4813" />
                    <RANKING order="5" place="5" resultid="5554" />
                    <RANKING order="6" place="-1" resultid="3663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1950" />
                    <RANKING order="2" place="2" resultid="4245" />
                    <RANKING order="3" place="3" resultid="5561" />
                    <RANKING order="4" place="4" resultid="6195" />
                    <RANKING order="5" place="5" resultid="4851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6392" />
                    <RANKING order="2" place="2" resultid="1792" />
                    <RANKING order="3" place="3" resultid="2148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3137" />
                    <RANKING order="2" place="2" resultid="6282" />
                    <RANKING order="3" place="3" resultid="5573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6844" />
                    <RANKING order="2" place="2" resultid="6144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3466" />
                    <RANKING order="2" place="2" resultid="7272" />
                    <RANKING order="3" place="3" resultid="6022" />
                    <RANKING order="4" place="4" resultid="2241" />
                    <RANKING order="5" place="-1" resultid="2331" />
                    <RANKING order="6" place="-1" resultid="3194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4005" />
                    <RANKING order="2" place="-1" resultid="1999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1160" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1161" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1162" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1163" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1164" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8936" daytime="18:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8937" daytime="18:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8938" daytime="18:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8939" daytime="19:10" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2015-11-14" daytime="09:00" name="BLOK II" number="2" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1222" daytime="09:30" gender="F" number="10" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1223" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3603" />
                    <RANKING order="2" place="2" resultid="4176" />
                    <RANKING order="3" place="3" resultid="2837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2232" />
                    <RANKING order="2" place="2" resultid="6243" />
                    <RANKING order="3" place="3" resultid="7004" />
                    <RANKING order="4" place="4" resultid="2509" />
                    <RANKING order="5" place="5" resultid="5779" />
                    <RANKING order="6" place="-1" resultid="7159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2517" />
                    <RANKING order="2" place="2" resultid="4963" />
                    <RANKING order="3" place="3" resultid="3866" />
                    <RANKING order="4" place="4" resultid="5555" />
                    <RANKING order="5" place="5" resultid="3750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5562" />
                    <RANKING order="2" place="2" resultid="2769" />
                    <RANKING order="3" place="3" resultid="3203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6393" />
                    <RANKING order="2" place="2" resultid="3924" />
                    <RANKING order="3" place="3" resultid="2444" />
                    <RANKING order="4" place="4" resultid="2615" />
                    <RANKING order="5" place="5" resultid="3457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2643" />
                    <RANKING order="2" place="2" resultid="6283" />
                    <RANKING order="3" place="3" resultid="5574" />
                    <RANKING order="4" place="4" resultid="2862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3970" />
                    <RANKING order="2" place="2" resultid="3402" />
                    <RANKING order="3" place="3" resultid="2346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6839" />
                    <RANKING order="2" place="2" resultid="7361" />
                    <RANKING order="3" place="3" resultid="6023" />
                    <RANKING order="4" place="4" resultid="3186" />
                    <RANKING order="5" place="5" resultid="2339" />
                    <RANKING order="6" place="6" resultid="6875" />
                    <RANKING order="7" place="7" resultid="2242" />
                    <RANKING order="8" place="8" resultid="2332" />
                    <RANKING order="9" place="-1" resultid="5793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3002" />
                    <RANKING order="2" place="2" resultid="3162" />
                    <RANKING order="3" place="3" resultid="3336" />
                    <RANKING order="4" place="4" resultid="2351" />
                    <RANKING order="5" place="5" resultid="1819" />
                    <RANKING order="6" place="-1" resultid="6164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7291" />
                    <RANKING order="2" place="2" resultid="2001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1235" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1236" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1237" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1238" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8966" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8967" daytime="09:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8968" daytime="09:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8969" daytime="09:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8970" daytime="09:55" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="12:20" gender="F" number="16" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1325" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1326" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6244" />
                    <RANKING order="2" place="2" resultid="3379" />
                    <RANKING order="3" place="3" resultid="2233" />
                    <RANKING order="4" place="4" resultid="3960" />
                    <RANKING order="5" place="5" resultid="7012" />
                    <RANKING order="6" place="6" resultid="5786" />
                    <RANKING order="7" place="-1" resultid="2510" />
                    <RANKING order="8" place="-1" resultid="3346" />
                    <RANKING order="9" place="-1" resultid="7005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3985" />
                    <RANKING order="2" place="2" resultid="6189" />
                    <RANKING order="3" place="3" resultid="6204" />
                    <RANKING order="4" place="4" resultid="4971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1328" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1329" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1330" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="1331" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3403" />
                    <RANKING order="2" place="2" resultid="6145" />
                    <RANKING order="3" place="3" resultid="6869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1332" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7274" />
                    <RANKING order="2" place="2" resultid="3187" />
                    <RANKING order="3" place="3" resultid="2243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1333" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1334" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1335" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1336" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1337" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1338" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1339" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1340" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9022" daytime="12:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9023" daytime="12:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9024" daytime="12:30" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1239" daytime="10:00" gender="M" number="11" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1240" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5948" />
                    <RANKING order="2" place="2" resultid="6337" />
                    <RANKING order="3" place="3" resultid="4151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3169" />
                    <RANKING order="2" place="2" resultid="4165" />
                    <RANKING order="3" place="3" resultid="7365" />
                    <RANKING order="4" place="4" resultid="3850" />
                    <RANKING order="5" place="5" resultid="1778" />
                    <RANKING order="6" place="-1" resultid="4171" />
                    <RANKING order="7" place="-1" resultid="7025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3858" />
                    <RANKING order="2" place="2" resultid="4764" />
                    <RANKING order="3" place="3" resultid="6209" />
                    <RANKING order="4" place="-1" resultid="7060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6260" />
                    <RANKING order="2" place="2" resultid="3534" />
                    <RANKING order="3" place="3" resultid="3912" />
                    <RANKING order="4" place="4" resultid="2651" />
                    <RANKING order="5" place="5" resultid="7382" />
                    <RANKING order="6" place="6" resultid="2685" />
                    <RANKING order="7" place="7" resultid="2101" />
                    <RANKING order="8" place="8" resultid="4771" />
                    <RANKING order="9" place="9" resultid="5810" />
                    <RANKING order="10" place="-1" resultid="3731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4956" />
                    <RANKING order="2" place="2" resultid="4232" />
                    <RANKING order="3" place="3" resultid="2729" />
                    <RANKING order="4" place="4" resultid="1895" />
                    <RANKING order="5" place="5" resultid="5774" />
                    <RANKING order="6" place="6" resultid="3422" />
                    <RANKING order="7" place="7" resultid="5879" />
                    <RANKING order="8" place="8" resultid="2812" />
                    <RANKING order="9" place="-1" resultid="4947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2797" />
                    <RANKING order="2" place="2" resultid="4622" />
                    <RANKING order="3" place="3" resultid="2193" />
                    <RANKING order="4" place="4" resultid="2461" />
                    <RANKING order="5" place="5" resultid="7311" />
                    <RANKING order="6" place="6" resultid="3950" />
                    <RANKING order="7" place="7" resultid="5547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3392" />
                    <RANKING order="2" place="2" resultid="6862" />
                    <RANKING order="3" place="3" resultid="6237" />
                    <RANKING order="4" place="4" resultid="5094" />
                    <RANKING order="5" place="5" resultid="3384" />
                    <RANKING order="6" place="6" resultid="5679" />
                    <RANKING order="7" place="-1" resultid="3885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5863" />
                    <RANKING order="2" place="2" resultid="2981" />
                    <RANKING order="3" place="3" resultid="4667" />
                    <RANKING order="4" place="4" resultid="3567" />
                    <RANKING order="5" place="5" resultid="2323" />
                    <RANKING order="6" place="-1" resultid="3154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2184" />
                    <RANKING order="2" place="2" resultid="2938" />
                    <RANKING order="3" place="3" resultid="3561" />
                    <RANKING order="4" place="4" resultid="3016" />
                    <RANKING order="5" place="5" resultid="2577" />
                    <RANKING order="6" place="6" resultid="2591" />
                    <RANKING order="7" place="7" resultid="1976" />
                    <RANKING order="8" place="-1" resultid="5725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1249" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3488" />
                    <RANKING order="2" place="2" resultid="3021" />
                    <RANKING order="3" place="3" resultid="2480" />
                    <RANKING order="4" place="4" resultid="2274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1786" />
                    <RANKING order="2" place="2" resultid="2314" />
                    <RANKING order="3" place="3" resultid="1991" />
                    <RANKING order="4" place="4" resultid="3327" />
                    <RANKING order="5" place="-1" resultid="2954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6366" />
                    <RANKING order="2" place="2" resultid="3826" />
                    <RANKING order="3" place="3" resultid="5849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1254" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1255" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8971" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8972" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8973" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8974" daytime="10:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8975" daytime="10:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8976" daytime="10:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8977" daytime="10:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8978" daytime="10:35" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1256" daytime="10:35" gender="F" number="12" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1257" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2782" />
                    <RANKING order="2" place="2" resultid="5625" />
                    <RANKING order="3" place="3" resultid="7135" />
                    <RANKING order="4" place="4" resultid="6342" />
                    <RANKING order="5" place="5" resultid="4184" />
                    <RANKING order="6" place="6" resultid="4177" />
                    <RANKING order="7" place="7" resultid="1812" />
                    <RANKING order="8" place="8" resultid="6895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4872" />
                    <RANKING order="2" place="2" resultid="1939" />
                    <RANKING order="3" place="3" resultid="7128" />
                    <RANKING order="4" place="4" resultid="3416" />
                    <RANKING order="5" place="5" resultid="3378" />
                    <RANKING order="6" place="6" resultid="5969" />
                    <RANKING order="7" place="7" resultid="5910" />
                    <RANKING order="8" place="8" resultid="3947" />
                    <RANKING order="9" place="9" resultid="2080" />
                    <RANKING order="10" place="10" resultid="7167" />
                    <RANKING order="11" place="11" resultid="5109" />
                    <RANKING order="12" place="12" resultid="6140" />
                    <RANKING order="13" place="13" resultid="6030" />
                    <RANKING order="14" place="-1" resultid="5656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3441" />
                    <RANKING order="2" place="2" resultid="4964" />
                    <RANKING order="3" place="3" resultid="4814" />
                    <RANKING order="4" place="4" resultid="5905" />
                    <RANKING order="5" place="5" resultid="6203" />
                    <RANKING order="6" place="6" resultid="3682" />
                    <RANKING order="7" place="7" resultid="4791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1951" />
                    <RANKING order="2" place="2" resultid="4753" />
                    <RANKING order="3" place="3" resultid="6196" />
                    <RANKING order="4" place="4" resultid="4263" />
                    <RANKING order="5" place="5" resultid="4852" />
                    <RANKING order="6" place="6" resultid="3204" />
                    <RANKING order="7" place="-1" resultid="4255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2149" />
                    <RANKING order="2" place="2" resultid="7256" />
                    <RANKING order="3" place="3" resultid="2776" />
                    <RANKING order="4" place="4" resultid="6019" />
                    <RANKING order="5" place="5" resultid="7378" />
                    <RANKING order="6" place="6" resultid="4798" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7244" />
                    <RANKING order="2" place="2" resultid="5615" />
                    <RANKING order="3" place="3" resultid="6284" />
                    <RANKING order="4" place="4" resultid="5869" />
                    <RANKING order="5" place="-1" resultid="5669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3528" />
                    <RANKING order="2" place="2" resultid="6845" />
                    <RANKING order="3" place="3" resultid="3334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7273" />
                    <RANKING order="2" place="2" resultid="3195" />
                    <RANKING order="3" place="3" resultid="2340" />
                    <RANKING order="4" place="4" resultid="2333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6403" />
                    <RANKING order="2" place="2" resultid="3931" />
                    <RANKING order="3" place="3" resultid="5665" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1269" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1270" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1271" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1272" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8979" daytime="10:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8980" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8981" daytime="10:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8982" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8983" daytime="10:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8984" daytime="10:50" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1358" daytime="13:05" gender="F" number="18" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1375" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8604" />
                    <RANKING order="2" place="-1" resultid="7527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1376" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6300" />
                    <RANKING order="2" place="2" resultid="2871" />
                    <RANKING order="3" place="3" resultid="5826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1377" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3626" />
                    <RANKING order="2" place="2" resultid="5598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1378" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7400" />
                    <RANKING order="2" place="2" resultid="6913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1379" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1380" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9031" daytime="13:05" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1307" daytime="11:45" gender="M" number="15" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1308" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5949" />
                    <RANKING order="2" place="2" resultid="5634" />
                    <RANKING order="3" place="3" resultid="1803" />
                    <RANKING order="4" place="4" resultid="5533" />
                    <RANKING order="5" place="5" resultid="2120" />
                    <RANKING order="6" place="6" resultid="6346" />
                    <RANKING order="7" place="7" resultid="3357" />
                    <RANKING order="8" place="-1" resultid="5080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4720" />
                    <RANKING order="2" place="2" resultid="5769" />
                    <RANKING order="3" place="3" resultid="3594" />
                    <RANKING order="4" place="4" resultid="5105" />
                    <RANKING order="5" place="5" resultid="4837" />
                    <RANKING order="6" place="6" resultid="4879" />
                    <RANKING order="7" place="7" resultid="2852" />
                    <RANKING order="8" place="8" resultid="7366" />
                    <RANKING order="9" place="9" resultid="4914" />
                    <RANKING order="10" place="10" resultid="7144" />
                    <RANKING order="11" place="11" resultid="3495" />
                    <RANKING order="12" place="12" resultid="4217" />
                    <RANKING order="13" place="13" resultid="3851" />
                    <RANKING order="14" place="14" resultid="3170" />
                    <RANKING order="15" place="15" resultid="1779" />
                    <RANKING order="16" place="16" resultid="7026" />
                    <RANKING order="17" place="17" resultid="4918" />
                    <RANKING order="18" place="18" resultid="1934" />
                    <RANKING order="19" place="19" resultid="2131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7190" />
                    <RANKING order="2" place="2" resultid="2113" />
                    <RANKING order="3" place="3" resultid="2086" />
                    <RANKING order="4" place="4" resultid="3720" />
                    <RANKING order="5" place="5" resultid="7240" />
                    <RANKING order="6" place="6" resultid="4714" />
                    <RANKING order="7" place="7" resultid="4765" />
                    <RANKING order="8" place="8" resultid="5922" />
                    <RANKING order="9" place="9" resultid="2748" />
                    <RANKING order="10" place="10" resultid="6210" />
                    <RANKING order="11" place="11" resultid="4780" />
                    <RANKING order="12" place="12" resultid="4887" />
                    <RANKING order="13" place="-1" resultid="5980" />
                    <RANKING order="14" place="-1" resultid="7359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4010" />
                    <RANKING order="2" place="2" resultid="2806" />
                    <RANKING order="3" place="3" resultid="3690" />
                    <RANKING order="4" place="4" resultid="2599" />
                    <RANKING order="5" place="5" resultid="6261" />
                    <RANKING order="6" place="6" resultid="2154" />
                    <RANKING order="7" place="7" resultid="5944" />
                    <RANKING order="8" place="8" resultid="5719" />
                    <RANKING order="9" place="9" resultid="2661" />
                    <RANKING order="10" place="10" resultid="2017" />
                    <RANKING order="11" place="11" resultid="3796" />
                    <RANKING order="12" place="12" resultid="4865" />
                    <RANKING order="13" place="13" resultid="3942" />
                    <RANKING order="14" place="14" resultid="3701" />
                    <RANKING order="15" place="15" resultid="2102" />
                    <RANKING order="16" place="16" resultid="2398" />
                    <RANKING order="17" place="17" resultid="4772" />
                    <RANKING order="18" place="-1" resultid="2040" />
                    <RANKING order="19" place="-1" resultid="3706" />
                    <RANKING order="20" place="-1" resultid="3732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2703" />
                    <RANKING order="2" place="2" resultid="4283" />
                    <RANKING order="3" place="3" resultid="2266" />
                    <RANKING order="4" place="4" resultid="4233" />
                    <RANKING order="5" place="5" resultid="3557" />
                    <RANKING order="6" place="6" resultid="3784" />
                    <RANKING order="7" place="7" resultid="7374" />
                    <RANKING order="8" place="8" resultid="3423" />
                    <RANKING order="9" place="9" resultid="4271" />
                    <RANKING order="10" place="10" resultid="5965" />
                    <RANKING order="11" place="11" resultid="6177" />
                    <RANKING order="12" place="12" resultid="7048" />
                    <RANKING order="13" place="13" resultid="4786" />
                    <RANKING order="14" place="-1" resultid="4922" />
                    <RANKING order="15" place="-1" resultid="6352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4830" />
                    <RANKING order="2" place="2" resultid="3352" />
                    <RANKING order="3" place="3" resultid="3835" />
                    <RANKING order="4" place="4" resultid="4822" />
                    <RANKING order="5" place="5" resultid="4073" />
                    <RANKING order="6" place="6" resultid="2055" />
                    <RANKING order="7" place="7" resultid="4077" />
                    <RANKING order="8" place="8" resultid="6857" />
                    <RANKING order="9" place="9" resultid="5818" />
                    <RANKING order="10" place="10" resultid="2462" />
                    <RANKING order="11" place="11" resultid="4289" />
                    <RANKING order="12" place="12" resultid="4927" />
                    <RANKING order="13" place="13" resultid="6290" />
                    <RANKING order="14" place="14" resultid="2010" />
                    <RANKING order="15" place="15" resultid="1901" />
                    <RANKING order="16" place="-1" resultid="4623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4225" />
                    <RANKING order="2" place="2" resultid="2047" />
                    <RANKING order="3" place="3" resultid="6152" />
                    <RANKING order="4" place="4" resultid="7305" />
                    <RANKING order="5" place="5" resultid="3233" />
                    <RANKING order="6" place="6" resultid="6863" />
                    <RANKING order="7" place="-1" resultid="3586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5099" />
                    <RANKING order="2" place="2" resultid="3792" />
                    <RANKING order="3" place="3" resultid="7114" />
                    <RANKING order="4" place="4" resultid="2607" />
                    <RANKING order="5" place="5" resultid="3991" />
                    <RANKING order="6" place="6" resultid="2571" />
                    <RANKING order="7" place="7" resultid="2301" />
                    <RANKING order="8" place="-1" resultid="3479" />
                    <RANKING order="9" place="-1" resultid="3568" />
                    <RANKING order="10" place="-1" resultid="5864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1316" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2185" />
                    <RANKING order="2" place="2" resultid="3966" />
                    <RANKING order="3" place="3" resultid="2939" />
                    <RANKING order="4" place="4" resultid="4660" />
                    <RANKING order="5" place="5" resultid="3012" />
                    <RANKING order="6" place="6" resultid="1908" />
                    <RANKING order="7" place="7" resultid="5646" />
                    <RANKING order="8" place="8" resultid="2525" />
                    <RANKING order="9" place="9" resultid="2578" />
                    <RANKING order="10" place="10" resultid="3146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1317" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2678" />
                    <RANKING order="2" place="2" resultid="2035" />
                    <RANKING order="3" place="3" resultid="3512" />
                    <RANKING order="4" place="4" resultid="2308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1318" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1787" />
                    <RANKING order="2" place="2" resultid="4647" />
                    <RANKING order="3" place="3" resultid="3364" />
                    <RANKING order="4" place="4" resultid="1882" />
                    <RANKING order="5" place="5" resultid="7263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1319" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6382" />
                    <RANKING order="2" place="2" resultid="2995" />
                    <RANKING order="3" place="3" resultid="3827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1320" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1321" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1322" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1323" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9008" daytime="11:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9009" daytime="11:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9010" daytime="11:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9011" daytime="11:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9012" daytime="11:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9013" daytime="12:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9014" daytime="12:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9015" daytime="12:05" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9016" daytime="12:05" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9017" daytime="12:10" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9018" daytime="12:10" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="9019" daytime="12:10" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="9020" daytime="12:15" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="9021" daytime="12:15" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1341" daytime="12:35" gender="M" number="17" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1342" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6906" />
                    <RANKING order="2" place="2" resultid="1804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4683" />
                    <RANKING order="2" place="2" resultid="7041" />
                    <RANKING order="3" place="3" resultid="4909" />
                    <RANKING order="4" place="4" resultid="2202" />
                    <RANKING order="5" place="5" resultid="4159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7191" />
                    <RANKING order="2" place="2" resultid="2542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6882" />
                    <RANKING order="2" place="2" resultid="3913" />
                    <RANKING order="3" place="3" resultid="4895" />
                    <RANKING order="4" place="4" resultid="2652" />
                    <RANKING order="5" place="5" resultid="2686" />
                    <RANKING order="6" place="6" resultid="5811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7318" />
                    <RANKING order="2" place="2" resultid="6223" />
                    <RANKING order="3" place="3" resultid="2210" />
                    <RANKING order="4" place="4" resultid="1874" />
                    <RANKING order="5" place="5" resultid="6178" />
                    <RANKING order="6" place="-1" resultid="4978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3918" />
                    <RANKING order="2" place="2" resultid="6133" />
                    <RANKING order="3" place="3" resultid="3409" />
                    <RANKING order="4" place="4" resultid="3180" />
                    <RANKING order="5" place="5" resultid="3951" />
                    <RANKING order="6" place="-1" resultid="2866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4807" />
                    <RANKING order="2" place="2" resultid="6832" />
                    <RANKING order="3" place="3" resultid="5932" />
                    <RANKING order="4" place="4" resultid="3587" />
                    <RANKING order="5" place="5" resultid="6850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6268" />
                    <RANKING order="2" place="2" resultid="3503" />
                    <RANKING order="3" place="3" resultid="7328" />
                    <RANKING order="4" place="4" resultid="2585" />
                    <RANKING order="5" place="5" resultid="2324" />
                    <RANKING order="6" place="-1" resultid="2407" />
                    <RANKING order="7" place="-1" resultid="3155" />
                    <RANKING order="8" place="-1" resultid="3480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1350" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3562" />
                    <RANKING order="2" place="2" resultid="5856" />
                    <RANKING order="3" place="3" resultid="1968" />
                    <RANKING order="4" place="4" resultid="2063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1351" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1928" />
                    <RANKING order="2" place="2" resultid="1915" />
                    <RANKING order="3" place="3" resultid="3022" />
                    <RANKING order="4" place="4" resultid="2625" />
                    <RANKING order="5" place="-1" resultid="2488" />
                    <RANKING order="6" place="-1" resultid="5698" />
                    <RANKING order="7" place="-1" resultid="7283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1355" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1356" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1357" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9025" daytime="12:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9026" daytime="12:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9027" daytime="12:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9028" daytime="12:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9029" daytime="12:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9030" daytime="13:00" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1381" daytime="13:10" gender="M" number="19" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1382" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2163" />
                    <RANKING order="2" place="-1" resultid="5988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1383" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3628" />
                    <RANKING order="2" place="2" resultid="7900" />
                    <RANKING order="3" place="3" resultid="7529" />
                    <RANKING order="4" place="4" resultid="3760" />
                    <RANKING order="5" place="5" resultid="2873" />
                    <RANKING order="6" place="6" resultid="8606" />
                    <RANKING order="7" place="7" resultid="4932" />
                    <RANKING order="8" place="8" resultid="5954" />
                    <RANKING order="9" place="9" resultid="7404" />
                    <RANKING order="10" place="10" resultid="8607" />
                    <RANKING order="11" place="11" resultid="3761" />
                    <RANKING order="12" place="12" resultid="2165" />
                    <RANKING order="13" place="-1" resultid="7067" />
                    <RANKING order="14" place="-1" resultid="7902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1384" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6914" />
                    <RANKING order="2" place="2" resultid="6168" />
                    <RANKING order="3" place="3" resultid="6301" />
                    <RANKING order="4" place="4" resultid="7402" />
                    <RANKING order="5" place="5" resultid="4295" />
                    <RANKING order="6" place="6" resultid="5824" />
                    <RANKING order="7" place="7" resultid="3671" />
                    <RANKING order="8" place="8" resultid="3240" />
                    <RANKING order="9" place="9" resultid="6303" />
                    <RANKING order="10" place="-1" resultid="2433" />
                    <RANKING order="11" place="-1" resultid="5743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1385" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2709" />
                    <RANKING order="2" place="2" resultid="3630" />
                    <RANKING order="3" place="3" resultid="2967" />
                    <RANKING order="4" place="4" resultid="2358" />
                    <RANKING order="5" place="-1" resultid="2875" />
                    <RANKING order="6" place="-1" resultid="2023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1386" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4677" />
                    <RANKING order="2" place="2" resultid="7405" />
                    <RANKING order="3" place="3" resultid="3036" />
                    <RANKING order="4" place="-1" resultid="3632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1387" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6418" />
                    <RANKING order="2" place="2" resultid="2552" />
                    <RANKING order="3" place="3" resultid="2360" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9032" daytime="13:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9033" daytime="13:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9034" daytime="13:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9035" daytime="13:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1273" daytime="10:50" gender="M" number="13" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1274" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5875" />
                    <RANKING order="2" place="2" resultid="6905" />
                    <RANKING order="3" place="3" resultid="5542" />
                    <RANKING order="4" place="4" resultid="2858" />
                    <RANKING order="5" place="5" resultid="5079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2094" />
                    <RANKING order="2" place="2" resultid="5768" />
                    <RANKING order="3" place="3" resultid="2138" />
                    <RANKING order="4" place="4" resultid="6327" />
                    <RANKING order="5" place="5" resultid="4710" />
                    <RANKING order="6" place="6" resultid="2791" />
                    <RANKING order="7" place="7" resultid="7143" />
                    <RANKING order="8" place="8" resultid="7040" />
                    <RANKING order="9" place="9" resultid="2072" />
                    <RANKING order="10" place="10" resultid="4158" />
                    <RANKING order="11" place="11" resultid="3891" />
                    <RANKING order="12" place="12" resultid="4617" />
                    <RANKING order="13" place="13" resultid="1933" />
                    <RANKING order="14" place="14" resultid="2130" />
                    <RANKING order="15" place="-1" resultid="5072" />
                    <RANKING order="16" place="-1" resultid="5926" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3712" />
                    <RANKING order="2" place="2" resultid="2143" />
                    <RANKING order="3" place="3" resultid="5117" />
                    <RANKING order="4" place="4" resultid="7175" />
                    <RANKING order="5" place="5" resultid="2473" />
                    <RANKING order="6" place="6" resultid="5898" />
                    <RANKING order="7" place="7" resultid="7183" />
                    <RANKING order="8" place="8" resultid="2846" />
                    <RANKING order="9" place="9" resultid="5921" />
                    <RANKING order="10" place="10" resultid="5587" />
                    <RANKING order="11" place="11" resultid="2747" />
                    <RANKING order="12" place="12" resultid="4779" />
                    <RANKING order="13" place="13" resultid="2541" />
                    <RANKING order="14" place="14" resultid="4952" />
                    <RANKING order="15" place="15" resultid="4201" />
                    <RANKING order="16" place="16" resultid="4886" />
                    <RANKING order="17" place="17" resultid="2549" />
                    <RANKING order="18" place="-1" resultid="2726" />
                    <RANKING order="19" place="-1" resultid="3371" />
                    <RANKING order="20" place="-1" resultid="3859" />
                    <RANKING order="21" place="-1" resultid="5581" />
                    <RANKING order="22" place="-1" resultid="7239" />
                    <RANKING order="23" place="-1" resultid="7358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1773" />
                    <RANKING order="2" place="2" resultid="6881" />
                    <RANKING order="3" place="3" resultid="2805" />
                    <RANKING order="4" place="4" resultid="5915" />
                    <RANKING order="5" place="5" resultid="2502" />
                    <RANKING order="6" place="6" resultid="5943" />
                    <RANKING order="7" place="7" resultid="3689" />
                    <RANKING order="8" place="8" resultid="3700" />
                    <RANKING order="9" place="9" resultid="3757" />
                    <RANKING order="10" place="10" resultid="3978" />
                    <RANKING order="11" place="11" resultid="6276" />
                    <RANKING order="12" place="12" resultid="4864" />
                    <RANKING order="13" place="13" resultid="3879" />
                    <RANKING order="14" place="14" resultid="4941" />
                    <RANKING order="15" place="15" resultid="3696" />
                    <RANKING order="16" place="16" resultid="2107" />
                    <RANKING order="17" place="17" resultid="7299" />
                    <RANKING order="18" place="18" resultid="2397" />
                    <RANKING order="19" place="-1" resultid="3743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2702" />
                    <RANKING order="2" place="2" resultid="6222" />
                    <RANKING order="3" place="3" resultid="5730" />
                    <RANKING order="4" place="4" resultid="4688" />
                    <RANKING order="5" place="5" resultid="4282" />
                    <RANKING order="6" place="6" resultid="2670" />
                    <RANKING order="7" place="7" resultid="3783" />
                    <RANKING order="8" place="8" resultid="3905" />
                    <RANKING order="9" place="9" resultid="3216" />
                    <RANKING order="10" place="10" resultid="6006" />
                    <RANKING order="11" place="11" resultid="6000" />
                    <RANKING order="12" place="12" resultid="3936" />
                    <RANKING order="13" place="13" resultid="7250" />
                    <RANKING order="14" place="14" resultid="3956" />
                    <RANKING order="15" place="15" resultid="4240" />
                    <RANKING order="16" place="16" resultid="1896" />
                    <RANKING order="17" place="17" resultid="4760" />
                    <RANKING order="18" place="18" resultid="2423" />
                    <RANKING order="19" place="19" resultid="4785" />
                    <RANKING order="20" place="20" resultid="2160" />
                    <RANKING order="21" place="21" resultid="3226" />
                    <RANKING order="22" place="22" resultid="6230" />
                    <RANKING order="23" place="23" resultid="3238" />
                    <RANKING order="24" place="-1" resultid="2265" />
                    <RANKING order="25" place="-1" resultid="4921" />
                    <RANKING order="26" place="-1" resultid="5687" />
                    <RANKING order="27" place="-1" resultid="6351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4821" />
                    <RANKING order="2" place="2" resultid="4072" />
                    <RANKING order="3" place="3" resultid="3179" />
                    <RANKING order="4" place="4" resultid="3397" />
                    <RANKING order="5" place="5" resultid="2054" />
                    <RANKING order="6" place="6" resultid="2946" />
                    <RANKING order="7" place="7" resultid="7117" />
                    <RANKING order="8" place="8" resultid="2009" />
                    <RANKING order="9" place="9" resultid="7312" />
                    <RANKING order="10" place="10" resultid="2962" />
                    <RANKING order="11" place="11" resultid="3897" />
                    <RANKING order="12" place="12" resultid="2415" />
                    <RANKING order="13" place="13" resultid="5548" />
                    <RANKING order="14" place="14" resultid="1900" />
                    <RANKING order="15" place="15" resultid="7371" />
                    <RANKING order="16" place="-1" resultid="2798" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3886" />
                    <RANKING order="2" place="2" resultid="6899" />
                    <RANKING order="3" place="3" resultid="7107" />
                    <RANKING order="4" place="4" resultid="3455" />
                    <RANKING order="5" place="5" resultid="2046" />
                    <RANKING order="6" place="6" resultid="5091" />
                    <RANKING order="7" place="7" resultid="5931" />
                    <RANKING order="8" place="8" resultid="3580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3791" />
                    <RANKING order="2" place="2" resultid="2694" />
                    <RANKING order="3" place="3" resultid="5884" />
                    <RANKING order="4" place="4" resultid="7113" />
                    <RANKING order="5" place="5" resultid="2565" />
                    <RANKING order="6" place="6" resultid="7343" />
                    <RANKING order="7" place="7" resultid="3872" />
                    <RANKING order="8" place="8" resultid="3220" />
                    <RANKING order="9" place="9" resultid="7327" />
                    <RANKING order="10" place="10" resultid="7389" />
                    <RANKING order="11" place="-1" resultid="3132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3965" />
                    <RANKING order="2" place="2" resultid="1889" />
                    <RANKING order="3" place="3" resultid="2634" />
                    <RANKING order="4" place="4" resultid="3011" />
                    <RANKING order="5" place="5" resultid="5855" />
                    <RANKING order="6" place="6" resultid="2386" />
                    <RANKING order="7" place="7" resultid="3145" />
                    <RANKING order="8" place="8" resultid="2287" />
                    <RANKING order="9" place="9" resultid="1977" />
                    <RANKING order="10" place="10" resultid="2821" />
                    <RANKING order="11" place="11" resultid="3129" />
                    <RANKING order="12" place="-1" resultid="5707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3818" />
                    <RANKING order="2" place="2" resultid="7282" />
                    <RANKING order="3" place="3" resultid="3511" />
                    <RANKING order="4" place="4" resultid="6399" />
                    <RANKING order="5" place="5" resultid="1945" />
                    <RANKING order="6" place="6" resultid="2487" />
                    <RANKING order="7" place="7" resultid="2275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3843" />
                    <RANKING order="2" place="2" resultid="1881" />
                    <RANKING order="3" place="3" resultid="1992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7226" />
                    <RANKING order="2" place="2" resultid="7100" />
                    <RANKING order="3" place="3" resultid="7336" />
                    <RANKING order="4" place="4" resultid="2496" />
                    <RANKING order="5" place="5" resultid="1985" />
                    <RANKING order="6" place="6" resultid="2295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8985" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8986" daytime="10:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8987" daytime="10:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8988" daytime="11:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8989" daytime="11:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8990" daytime="11:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8991" daytime="11:05" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8992" daytime="11:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8993" daytime="11:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8994" daytime="11:15" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="8995" daytime="11:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="8996" daytime="11:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="8997" daytime="11:20" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="8998" daytime="11:20" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="8999" daytime="11:25" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="9000" daytime="11:25" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="09:10" gender="M" number="9" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1206" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5874" />
                    <RANKING order="2" place="2" resultid="5541" />
                    <RANKING order="3" place="3" resultid="5633" />
                    <RANKING order="4" place="4" resultid="6336" />
                    <RANKING order="5" place="5" resultid="5532" />
                    <RANKING order="6" place="6" resultid="2119" />
                    <RANKING order="7" place="7" resultid="6345" />
                    <RANKING order="8" place="8" resultid="3254" />
                    <RANKING order="9" place="-1" resultid="4150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2093" />
                    <RANKING order="2" place="2" resultid="4836" />
                    <RANKING order="3" place="3" resultid="2851" />
                    <RANKING order="4" place="4" resultid="4913" />
                    <RANKING order="5" place="5" resultid="4705" />
                    <RANKING order="6" place="6" resultid="4216" />
                    <RANKING order="7" place="7" resultid="4878" />
                    <RANKING order="8" place="8" resultid="3494" />
                    <RANKING order="9" place="-1" resultid="2201" />
                    <RANKING order="10" place="-1" resultid="4170" />
                    <RANKING order="11" place="-1" resultid="4717" />
                    <RANKING order="12" place="-1" resultid="5975" />
                    <RANKING order="13" place="-1" resultid="5984" />
                    <RANKING order="14" place="-1" resultid="5986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3473" />
                    <RANKING order="2" place="2" resultid="7174" />
                    <RANKING order="3" place="3" resultid="3719" />
                    <RANKING order="4" place="4" resultid="6889" />
                    <RANKING order="5" place="5" resultid="7238" />
                    <RANKING order="6" place="6" resultid="5586" />
                    <RANKING order="7" place="7" resultid="2845" />
                    <RANKING order="8" place="8" resultid="7182" />
                    <RANKING order="9" place="9" resultid="3210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4691" />
                    <RANKING order="2" place="2" resultid="6130" />
                    <RANKING order="3" place="3" resultid="3599" />
                    <RANKING order="4" place="4" resultid="2598" />
                    <RANKING order="5" place="5" resultid="1772" />
                    <RANKING order="6" place="6" resultid="2660" />
                    <RANKING order="7" place="7" resultid="6275" />
                    <RANKING order="8" place="8" resultid="2016" />
                    <RANKING order="9" place="9" resultid="3533" />
                    <RANKING order="10" place="10" resultid="5938" />
                    <RANKING order="11" place="11" resultid="3737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2669" />
                    <RANKING order="2" place="2" resultid="2426" />
                    <RANKING order="3" place="3" resultid="3556" />
                    <RANKING order="4" place="4" resultid="3904" />
                    <RANKING order="5" place="5" resultid="4276" />
                    <RANKING order="6" place="6" resultid="4270" />
                    <RANKING order="7" place="7" resultid="5964" />
                    <RANKING order="8" place="8" resultid="4759" />
                    <RANKING order="9" place="-1" resultid="2209" />
                    <RANKING order="10" place="-1" resultid="5686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3917" />
                    <RANKING order="2" place="2" resultid="4829" />
                    <RANKING order="3" place="3" resultid="3834" />
                    <RANKING order="4" place="4" resultid="3447" />
                    <RANKING order="5" place="5" resultid="6856" />
                    <RANKING order="6" place="6" resultid="5817" />
                    <RANKING order="7" place="7" resultid="2192" />
                    <RANKING order="8" place="8" resultid="4926" />
                    <RANKING order="9" place="9" resultid="3896" />
                    <RANKING order="10" place="10" resultid="2945" />
                    <RANKING order="11" place="11" resultid="2961" />
                    <RANKING order="12" place="-1" resultid="6334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7106" />
                    <RANKING order="2" place="2" resultid="4224" />
                    <RANKING order="3" place="3" resultid="5090" />
                    <RANKING order="4" place="4" resultid="6151" />
                    <RANKING order="5" place="5" resultid="7304" />
                    <RANKING order="6" place="6" resultid="8881" />
                    <RANKING order="7" place="7" resultid="3232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5098" />
                    <RANKING order="2" place="2" resultid="2693" />
                    <RANKING order="3" place="3" resultid="3502" />
                    <RANKING order="4" place="4" resultid="2980" />
                    <RANKING order="5" place="5" resultid="6376" />
                    <RANKING order="6" place="6" resultid="2564" />
                    <RANKING order="7" place="7" resultid="2606" />
                    <RANKING order="8" place="8" resultid="3990" />
                    <RANKING order="9" place="9" resultid="3219" />
                    <RANKING order="10" place="10" resultid="2300" />
                    <RANKING order="11" place="11" resultid="7388" />
                    <RANKING order="12" place="-1" resultid="3131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1907" />
                    <RANKING order="2" place="2" resultid="2062" />
                    <RANKING order="3" place="3" resultid="2633" />
                    <RANKING order="4" place="4" resultid="4659" />
                    <RANKING order="5" place="5" resultid="1967" />
                    <RANKING order="6" place="6" resultid="4653" />
                    <RANKING order="7" place="7" resultid="2590" />
                    <RANKING order="8" place="8" resultid="2820" />
                    <RANKING order="9" place="9" resultid="2286" />
                    <RANKING order="10" place="10" resultid="3128" />
                    <RANKING order="11" place="-1" resultid="5724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2034" />
                    <RANKING order="2" place="2" resultid="2677" />
                    <RANKING order="3" place="3" resultid="1914" />
                    <RANKING order="4" place="4" resultid="6355" />
                    <RANKING order="5" place="5" resultid="3817" />
                    <RANKING order="6" place="6" resultid="2624" />
                    <RANKING order="7" place="7" resultid="2307" />
                    <RANKING order="8" place="8" resultid="2479" />
                    <RANKING order="9" place="9" resultid="6360" />
                    <RANKING order="10" place="10" resultid="7321" />
                    <RANKING order="11" place="-1" resultid="5641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4646" />
                    <RANKING order="2" place="2" resultid="3363" />
                    <RANKING order="3" place="3" resultid="2953" />
                    <RANKING order="4" place="4" resultid="7262" />
                    <RANKING order="5" place="5" resultid="3326" />
                    <RANKING order="6" place="-1" resultid="3842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2994" />
                    <RANKING order="2" place="2" resultid="7099" />
                    <RANKING order="3" place="3" resultid="1958" />
                    <RANKING order="4" place="4" resultid="5848" />
                    <RANKING order="5" place="5" resultid="2495" />
                    <RANKING order="6" place="6" resultid="1984" />
                    <RANKING order="7" place="-1" resultid="2294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1219" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1221" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8954" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8955" daytime="09:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8956" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8957" daytime="09:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8958" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8959" daytime="09:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8960" daytime="09:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8961" daytime="09:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8962" daytime="09:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8963" daytime="09:25" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="8964" daytime="09:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="8965" daytime="09:30" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1187" daytime="09:00" gender="F" number="8" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7054" />
                    <RANKING order="2" place="2" resultid="6341" />
                    <RANKING order="3" place="3" resultid="7018" />
                    <RANKING order="4" place="4" resultid="5763" />
                    <RANKING order="5" place="5" resultid="7134" />
                    <RANKING order="6" place="6" resultid="2756" />
                    <RANKING order="7" place="7" resultid="2125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7218" />
                    <RANKING order="2" place="2" resultid="3573" />
                    <RANKING order="3" place="3" resultid="4871" />
                    <RANKING order="4" place="4" resultid="3430" />
                    <RANKING order="5" place="5" resultid="3415" />
                    <RANKING order="6" place="6" resultid="4844" />
                    <RANKING order="7" place="7" resultid="3959" />
                    <RANKING order="8" place="8" resultid="7166" />
                    <RANKING order="9" place="9" resultid="2079" />
                    <RANKING order="10" place="-1" resultid="4723" />
                    <RANKING order="11" place="-1" resultid="7158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2762" />
                    <RANKING order="2" place="2" resultid="4699" />
                    <RANKING order="3" place="3" resultid="2740" />
                    <RANKING order="4" place="4" resultid="3749" />
                    <RANKING order="5" place="-1" resultid="4016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2532" />
                    <RANKING order="2" place="2" resultid="2466" />
                    <RANKING order="3" place="3" resultid="6251" />
                    <RANKING order="4" place="4" resultid="4246" />
                    <RANKING order="5" place="5" resultid="5672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3548" />
                    <RANKING order="2" place="2" resultid="4210" />
                    <RANKING order="3" place="3" resultid="2775" />
                    <RANKING order="4" place="4" resultid="7255" />
                    <RANKING order="5" place="5" resultid="6018" />
                    <RANKING order="6" place="-1" resultid="6011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7231" />
                    <RANKING order="2" place="2" resultid="2453" />
                    <RANKING order="3" place="3" resultid="4204" />
                    <RANKING order="4" place="4" resultid="5593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3527" />
                    <RANKING order="2" place="2" resultid="6868" />
                    <RANKING order="3" place="3" resultid="2345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2987" />
                    <RANKING order="2" place="2" resultid="4639" />
                    <RANKING order="3" place="3" resultid="5087" />
                    <RANKING order="4" place="-1" resultid="5675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3030" />
                    <RANKING order="2" place="2" resultid="2350" />
                    <RANKING order="3" place="3" resultid="6163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5609" />
                    <RANKING order="2" place="2" resultid="3930" />
                    <RANKING order="3" place="3" resultid="4631" />
                    <RANKING order="4" place="4" resultid="2000" />
                    <RANKING order="5" place="-1" resultid="6363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5889" />
                    <RANKING order="2" place="2" resultid="1832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1202" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1203" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1204" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8948" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8949" daytime="09:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8950" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8951" daytime="09:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8952" daytime="09:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8953" daytime="09:10" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1290" daytime="11:25" gender="F" number="14" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1291" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2783" />
                    <RANKING order="2" place="2" resultid="7055" />
                    <RANKING order="3" place="3" resultid="5626" />
                    <RANKING order="4" place="4" resultid="7019" />
                    <RANKING order="5" place="5" resultid="4185" />
                    <RANKING order="6" place="6" resultid="3604" />
                    <RANKING order="7" place="7" resultid="1813" />
                    <RANKING order="8" place="8" resultid="7032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3574" />
                    <RANKING order="2" place="2" resultid="7219" />
                    <RANKING order="3" place="3" resultid="3810" />
                    <RANKING order="4" place="4" resultid="3431" />
                    <RANKING order="5" place="5" resultid="5970" />
                    <RANKING order="6" place="6" resultid="4845" />
                    <RANKING order="7" place="7" resultid="7011" />
                    <RANKING order="8" place="8" resultid="5780" />
                    <RANKING order="9" place="-1" resultid="7129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3436" />
                    <RANKING order="2" place="2" resultid="2763" />
                    <RANKING order="3" place="3" resultid="2518" />
                    <RANKING order="4" place="4" resultid="6188" />
                    <RANKING order="5" place="5" resultid="4021" />
                    <RANKING order="6" place="6" resultid="5556" />
                    <RANKING order="7" place="7" resultid="4017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2533" />
                    <RANKING order="2" place="2" resultid="6197" />
                    <RANKING order="3" place="3" resultid="6252" />
                    <RANKING order="4" place="4" resultid="2467" />
                    <RANKING order="5" place="5" resultid="4754" />
                    <RANKING order="6" place="6" resultid="4256" />
                    <RANKING order="7" place="7" resultid="4264" />
                    <RANKING order="8" place="8" resultid="6407" />
                    <RANKING order="9" place="9" resultid="4247" />
                    <RANKING order="10" place="10" resultid="2735" />
                    <RANKING order="11" place="11" resultid="4853" />
                    <RANKING order="12" place="12" resultid="2770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3549" />
                    <RANKING order="2" place="2" resultid="3925" />
                    <RANKING order="3" place="3" resultid="4904" />
                    <RANKING order="4" place="4" resultid="2445" />
                    <RANKING order="5" place="5" resultid="6012" />
                    <RANKING order="6" place="6" resultid="2616" />
                    <RANKING order="7" place="7" resultid="4799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7232" />
                    <RANKING order="2" place="2" resultid="7348" />
                    <RANKING order="3" place="3" resultid="2644" />
                    <RANKING order="4" place="4" resultid="5803" />
                    <RANKING order="5" place="5" resultid="4205" />
                    <RANKING order="6" place="6" resultid="2454" />
                    <RANKING order="7" place="7" resultid="5594" />
                    <RANKING order="8" place="8" resultid="5575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1298" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2391" />
                    <RANKING order="2" place="2" resultid="5794" />
                    <RANKING order="3" place="3" resultid="6024" />
                    <RANKING order="4" place="4" resultid="3196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1299" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3003" />
                    <RANKING order="2" place="2" resultid="3619" />
                    <RANKING order="3" place="3" resultid="1820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1300" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5610" />
                    <RANKING order="2" place="2" resultid="4632" />
                    <RANKING order="3" place="3" resultid="5569" />
                    <RANKING order="4" place="4" resultid="7292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1302" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1833" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1303" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1304" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1305" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1306" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9001" daytime="11:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9002" daytime="11:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9003" daytime="11:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9004" daytime="11:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9005" daytime="11:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9006" daytime="11:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9007" daytime="11:45" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2015-11-14" daytime="16:00" name="BLOK III" number="3" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="1440" daytime="17:00" gender="M" number="23" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1441" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5876" />
                    <RANKING order="2" place="2" resultid="5635" />
                    <RANKING order="3" place="3" resultid="5543" />
                    <RANKING order="4" place="4" resultid="6339" />
                    <RANKING order="5" place="5" resultid="5534" />
                    <RANKING order="6" place="6" resultid="3256" />
                    <RANKING order="7" place="-1" resultid="5081" />
                    <RANKING order="8" place="-1" resultid="6183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5770" />
                    <RANKING order="2" place="2" resultid="2095" />
                    <RANKING order="3" place="3" resultid="6328" />
                    <RANKING order="4" place="4" resultid="3614" />
                    <RANKING order="5" place="5" resultid="4706" />
                    <RANKING order="6" place="6" resultid="5107" />
                    <RANKING order="7" place="7" resultid="4711" />
                    <RANKING order="8" place="8" resultid="7145" />
                    <RANKING order="9" place="9" resultid="2139" />
                    <RANKING order="10" place="10" resultid="7368" />
                    <RANKING order="11" place="11" resultid="1922" />
                    <RANKING order="12" place="12" resultid="7042" />
                    <RANKING order="13" place="13" resultid="2792" />
                    <RANKING order="14" place="14" resultid="4919" />
                    <RANKING order="15" place="-1" resultid="1935" />
                    <RANKING order="16" place="-1" resultid="2203" />
                    <RANKING order="17" place="-1" resultid="4718" />
                    <RANKING order="18" place="-1" resultid="5073" />
                    <RANKING order="19" place="-1" resultid="5927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3713" />
                    <RANKING order="2" place="2" resultid="2114" />
                    <RANKING order="3" place="3" resultid="7192" />
                    <RANKING order="4" place="4" resultid="5981" />
                    <RANKING order="5" place="5" resultid="5118" />
                    <RANKING order="6" place="5" resultid="7176" />
                    <RANKING order="7" place="7" resultid="2144" />
                    <RANKING order="8" place="8" resultid="7184" />
                    <RANKING order="9" place="9" resultid="7241" />
                    <RANKING order="10" place="10" resultid="5899" />
                    <RANKING order="11" place="11" resultid="2847" />
                    <RANKING order="12" place="12" resultid="5923" />
                    <RANKING order="13" place="13" resultid="5582" />
                    <RANKING order="14" place="14" resultid="2750" />
                    <RANKING order="15" place="15" resultid="3211" />
                    <RANKING order="16" place="16" resultid="6212" />
                    <RANKING order="17" place="17" resultid="4781" />
                    <RANKING order="18" place="-1" resultid="4767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4692" />
                    <RANKING order="2" place="2" resultid="5916" />
                    <RANKING order="3" place="3" resultid="2807" />
                    <RANKING order="4" place="4" resultid="4011" />
                    <RANKING order="5" place="5" resultid="1774" />
                    <RANKING order="6" place="6" resultid="5945" />
                    <RANKING order="7" place="7" resultid="3702" />
                    <RANKING order="8" place="8" resultid="3691" />
                    <RANKING order="9" place="9" resultid="2155" />
                    <RANKING order="10" place="10" resultid="7383" />
                    <RANKING order="11" place="11" resultid="4896" />
                    <RANKING order="12" place="12" resultid="3979" />
                    <RANKING order="13" place="13" resultid="2018" />
                    <RANKING order="14" place="14" resultid="3880" />
                    <RANKING order="15" place="15" resultid="4866" />
                    <RANKING order="16" place="16" resultid="3744" />
                    <RANKING order="17" place="17" resultid="3943" />
                    <RANKING order="18" place="18" resultid="3798" />
                    <RANKING order="19" place="19" resultid="2108" />
                    <RANKING order="20" place="20" resultid="4774" />
                    <RANKING order="21" place="21" resultid="2399" />
                    <RANKING order="22" place="-1" resultid="3758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5731" />
                    <RANKING order="2" place="2" resultid="2704" />
                    <RANKING order="3" place="3" resultid="1875" />
                    <RANKING order="4" place="4" resultid="4284" />
                    <RANKING order="5" place="5" resultid="7268" />
                    <RANKING order="6" place="6" resultid="2267" />
                    <RANKING order="7" place="7" resultid="5713" />
                    <RANKING order="8" place="8" resultid="2671" />
                    <RANKING order="9" place="9" resultid="5800" />
                    <RANKING order="10" place="10" resultid="4277" />
                    <RANKING order="11" place="11" resultid="3906" />
                    <RANKING order="12" place="11" resultid="4235" />
                    <RANKING order="13" place="13" resultid="2211" />
                    <RANKING order="14" place="14" resultid="4272" />
                    <RANKING order="15" place="15" resultid="4761" />
                    <RANKING order="16" place="16" resultid="6179" />
                    <RANKING order="17" place="17" resultid="3425" />
                    <RANKING order="18" place="18" resultid="3227" />
                    <RANKING order="19" place="19" resultid="4787" />
                    <RANKING order="20" place="20" resultid="6231" />
                    <RANKING order="21" place="-1" resultid="2814" />
                    <RANKING order="22" place="-1" resultid="4923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3919" />
                    <RANKING order="2" place="2" resultid="4074" />
                    <RANKING order="3" place="3" resultid="5819" />
                    <RANKING order="4" place="4" resultid="2947" />
                    <RANKING order="5" place="5" resultid="4291" />
                    <RANKING order="6" place="6" resultid="2011" />
                    <RANKING order="7" place="7" resultid="6291" />
                    <RANKING order="8" place="8" resultid="2963" />
                    <RANKING order="9" place="9" resultid="2416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3888" />
                    <RANKING order="2" place="2" resultid="7108" />
                    <RANKING order="3" place="3" resultid="2048" />
                    <RANKING order="4" place="4" resultid="6153" />
                    <RANKING order="5" place="5" resultid="7306" />
                    <RANKING order="6" place="6" resultid="8882" />
                    <RANKING order="7" place="7" resultid="6833" />
                    <RANKING order="8" place="8" resultid="3581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6269" />
                    <RANKING order="2" place="2" resultid="5885" />
                    <RANKING order="3" place="3" resultid="7115" />
                    <RANKING order="4" place="4" resultid="6377" />
                    <RANKING order="5" place="5" resultid="4614" />
                    <RANKING order="6" place="6" resultid="7329" />
                    <RANKING order="7" place="7" resultid="2573" />
                    <RANKING order="8" place="8" resultid="3873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2187" />
                    <RANKING order="2" place="2" resultid="1890" />
                    <RANKING order="3" place="3" resultid="5857" />
                    <RANKING order="4" place="4" resultid="2526" />
                    <RANKING order="5" place="5" resultid="3147" />
                    <RANKING order="6" place="-1" resultid="2580" />
                    <RANKING order="7" place="-1" resultid="5708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6400" />
                    <RANKING order="2" place="2" resultid="1916" />
                    <RANKING order="3" place="3" resultid="3513" />
                    <RANKING order="4" place="4" resultid="1929" />
                    <RANKING order="5" place="5" resultid="7284" />
                    <RANKING order="6" place="6" resultid="6361" />
                    <RANKING order="7" place="-1" resultid="5699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1451" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1788" />
                    <RANKING order="2" place="2" resultid="3365" />
                    <RANKING order="3" place="3" resultid="2317" />
                    <RANKING order="4" place="4" resultid="1883" />
                    <RANKING order="5" place="5" resultid="7264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1452" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2997" />
                    <RANKING order="2" place="2" resultid="1960" />
                    <RANKING order="3" place="3" resultid="3829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1453" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1454" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1455" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1456" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9060" daytime="17:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9061" daytime="17:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9062" daytime="17:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9063" daytime="17:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9064" daytime="17:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9065" daytime="17:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9066" daytime="17:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9067" daytime="17:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9068" daytime="17:15" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9069" daytime="17:15" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9070" daytime="17:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="9071" daytime="17:20" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="9072" daytime="17:20" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="9073" daytime="17:20" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1457" daytime="17:25" gender="F" number="24" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1458" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5764" />
                    <RANKING order="2" place="2" resultid="2757" />
                    <RANKING order="3" place="3" resultid="6343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3576" />
                    <RANKING order="2" place="2" resultid="7221" />
                    <RANKING order="3" place="3" resultid="3433" />
                    <RANKING order="4" place="4" resultid="2234" />
                    <RANKING order="5" place="5" resultid="3417" />
                    <RANKING order="6" place="6" resultid="4846" />
                    <RANKING order="7" place="7" resultid="3961" />
                    <RANKING order="8" place="8" resultid="7169" />
                    <RANKING order="9" place="9" resultid="5110" />
                    <RANKING order="10" place="-1" resultid="2081" />
                    <RANKING order="11" place="-1" resultid="7161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1460" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2764" />
                    <RANKING order="2" place="2" resultid="4700" />
                    <RANKING order="3" place="3" resultid="2741" />
                    <RANKING order="4" place="-1" resultid="3752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1461" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2535" />
                    <RANKING order="2" place="2" resultid="2469" />
                    <RANKING order="3" place="3" resultid="4249" />
                    <RANKING order="4" place="4" resultid="6254" />
                    <RANKING order="5" place="-1" resultid="4266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1462" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3550" />
                    <RANKING order="2" place="2" resultid="4211" />
                    <RANKING order="3" place="3" resultid="4905" />
                    <RANKING order="4" place="4" resultid="7258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1463" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2455" />
                    <RANKING order="2" place="2" resultid="5596" />
                    <RANKING order="3" place="3" resultid="2863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1464" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3467" />
                    <RANKING order="2" place="2" resultid="2988" />
                    <RANKING order="3" place="3" resultid="3197" />
                    <RANKING order="4" place="4" resultid="4641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1466" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3033" />
                    <RANKING order="2" place="2" resultid="2353" />
                    <RANKING order="3" place="3" resultid="6166" />
                    <RANKING order="4" place="4" resultid="1822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5611" />
                    <RANKING order="2" place="2" resultid="3933" />
                    <RANKING order="3" place="3" resultid="4634" />
                    <RANKING order="4" place="4" resultid="5570" />
                    <RANKING order="5" place="5" resultid="2002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1468" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1469" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5891" />
                    <RANKING order="2" place="2" resultid="1835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1470" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1471" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1472" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1473" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9074" daytime="17:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9075" daytime="17:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9076" daytime="17:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9077" daytime="17:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9078" daytime="17:35" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1548" daytime="19:25" gender="M" number="29" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1549" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2164" />
                    <RANKING order="2" place="-1" resultid="7899" />
                    <RANKING order="3" place="-1" resultid="5987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1550" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3629" />
                    <RANKING order="2" place="2" resultid="7530" />
                    <RANKING order="3" place="3" resultid="2874" />
                    <RANKING order="4" place="4" resultid="3762" />
                    <RANKING order="5" place="5" resultid="5955" />
                    <RANKING order="6" place="6" resultid="4931" />
                    <RANKING order="7" place="7" resultid="8611" />
                    <RANKING order="8" place="8" resultid="7403" />
                    <RANKING order="9" place="9" resultid="2166" />
                    <RANKING order="10" place="10" resultid="3763" />
                    <RANKING order="11" place="-1" resultid="7068" />
                    <RANKING order="12" place="-1" resultid="7901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1551" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8610" />
                    <RANKING order="2" place="2" resultid="4857" />
                    <RANKING order="3" place="3" resultid="6918" />
                    <RANKING order="4" place="4" resultid="6302" />
                    <RANKING order="5" place="5" resultid="7401" />
                    <RANKING order="6" place="6" resultid="5744" />
                    <RANKING order="7" place="7" resultid="4296" />
                    <RANKING order="8" place="8" resultid="3239" />
                    <RANKING order="9" place="9" resultid="5823" />
                    <RANKING order="10" place="10" resultid="3670" />
                    <RANKING order="11" place="11" resultid="2432" />
                    <RANKING order="12" place="12" resultid="6304" />
                    <RANKING order="13" place="-1" resultid="8612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1552" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2708" />
                    <RANKING order="2" place="2" resultid="3631" />
                    <RANKING order="3" place="3" resultid="7120" />
                    <RANKING order="4" place="4" resultid="2968" />
                    <RANKING order="5" place="5" resultid="2876" />
                    <RANKING order="6" place="-1" resultid="2022" />
                    <RANKING order="7" place="-1" resultid="2359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1553" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1554" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6420" />
                    <RANKING order="2" place="2" resultid="7406" />
                    <RANKING order="3" place="3" resultid="2553" />
                    <RANKING order="4" place="4" resultid="2362" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9109" daytime="19:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9110" daytime="19:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9111" daytime="19:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9112" daytime="19:35" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1578" daytime="20:05" gender="M" number="31" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1579" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2260" />
                    <RANKING order="2" place="2" resultid="6908" />
                    <RANKING order="3" place="3" resultid="1806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1580" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4684" />
                    <RANKING order="2" place="2" resultid="4881" />
                    <RANKING order="3" place="3" resultid="4910" />
                    <RANKING order="4" place="4" resultid="2204" />
                    <RANKING order="5" place="5" resultid="3497" />
                    <RANKING order="6" place="6" resultid="1781" />
                    <RANKING order="7" place="-1" resultid="3172" />
                    <RANKING order="8" place="-1" resultid="4161" />
                    <RANKING order="9" place="-1" resultid="4173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1581" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7093" />
                    <RANKING order="2" place="2" resultid="3861" />
                    <RANKING order="3" place="3" resultid="2544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1582" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6884" />
                    <RANKING order="2" place="2" resultid="4012" />
                    <RANKING order="3" place="3" resultid="5720" />
                    <RANKING order="4" place="4" resultid="2663" />
                    <RANKING order="5" place="5" resultid="2654" />
                    <RANKING order="6" place="-1" resultid="3708" />
                    <RANKING order="7" place="-1" resultid="4897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6225" />
                    <RANKING order="2" place="2" resultid="2212" />
                    <RANKING order="3" place="3" resultid="7319" />
                    <RANKING order="4" place="4" resultid="4979" />
                    <RANKING order="5" place="-1" resultid="6002" />
                    <RANKING order="6" place="-1" resultid="4242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1584" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4824" />
                    <RANKING order="2" place="2" resultid="3411" />
                    <RANKING order="3" place="3" resultid="2800" />
                    <RANKING order="4" place="-1" resultid="2867" />
                    <RANKING order="5" place="-1" resultid="4625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6154" />
                    <RANKING order="2" place="2" resultid="4809" />
                    <RANKING order="3" place="3" resultid="8883" />
                    <RANKING order="4" place="4" resultid="6239" />
                    <RANKING order="5" place="5" resultid="5934" />
                    <RANKING order="6" place="6" resultid="6834" />
                    <RANKING order="7" place="7" resultid="3589" />
                    <RANKING order="8" place="-1" resultid="3386" />
                    <RANKING order="9" place="-1" resultid="6852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1586" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2696" />
                    <RANKING order="2" place="2" resultid="2409" />
                    <RANKING order="3" place="3" resultid="3482" />
                    <RANKING order="4" place="4" resultid="4669" />
                    <RANKING order="5" place="5" resultid="2612" />
                    <RANKING order="6" place="6" resultid="2586" />
                    <RANKING order="7" place="7" resultid="2326" />
                    <RANKING order="8" place="-1" resultid="3157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1587" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4662" />
                    <RANKING order="2" place="2" resultid="3564" />
                    <RANKING order="3" place="3" resultid="1970" />
                    <RANKING order="4" place="4" resultid="2941" />
                    <RANKING order="5" place="5" resultid="2527" />
                    <RANKING order="6" place="6" resultid="2593" />
                    <RANKING order="7" place="-1" resultid="1979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1588" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2680" />
                    <RANKING order="2" place="2" resultid="1917" />
                    <RANKING order="3" place="3" resultid="2627" />
                    <RANKING order="4" place="-1" resultid="2490" />
                    <RANKING order="5" place="-1" resultid="3024" />
                    <RANKING order="6" place="-1" resultid="5700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1589" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1590" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6383" />
                    <RANKING order="2" place="2" resultid="1961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1591" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1592" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1593" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1594" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9116" daytime="20:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9117" daytime="20:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9118" daytime="20:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9119" daytime="20:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9120" daytime="20:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9121" daytime="20:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9122" daytime="20:55" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1555" daytime="19:40" gender="F" number="30" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1562" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7056" />
                    <RANKING order="2" place="2" resultid="7021" />
                    <RANKING order="3" place="3" resultid="2758" />
                    <RANKING order="4" place="4" resultid="7034" />
                    <RANKING order="5" place="5" resultid="2840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1563" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6246" />
                    <RANKING order="2" place="2" resultid="7013" />
                    <RANKING order="3" place="3" resultid="2512" />
                    <RANKING order="4" place="4" resultid="5781" />
                    <RANKING order="5" place="-1" resultid="2235" />
                    <RANKING order="6" place="-1" resultid="3347" />
                    <RANKING order="7" place="-1" resultid="7007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1564" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2520" />
                    <RANKING order="2" place="2" resultid="6191" />
                    <RANKING order="3" place="3" resultid="4972" />
                    <RANKING order="4" place="-1" resultid="4794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1565" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1566" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3551" />
                    <RANKING order="2" place="2" resultid="6014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1567" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7350" />
                    <RANKING order="2" place="2" resultid="2646" />
                    <RANKING order="3" place="3" resultid="6286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1568" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6146" />
                    <RANKING order="2" place="2" resultid="6871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1569" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3468" />
                    <RANKING order="2" place="2" resultid="6026" />
                    <RANKING order="3" place="3" resultid="3189" />
                    <RANKING order="4" place="4" resultid="2245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1571" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1572" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1573" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1574" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1575" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1576" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1577" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9113" daytime="19:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9114" daytime="19:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9115" daytime="20:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1525" daytime="19:15" gender="F" number="28" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1542" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1543" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8608" />
                    <RANKING order="2" place="2" resultid="6299" />
                    <RANKING order="3" place="3" resultid="5825" />
                    <RANKING order="4" place="4" resultid="2872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1544" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3627" />
                    <RANKING order="2" place="-1" resultid="5597" />
                    <RANKING order="3" place="-1" resultid="6035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1545" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7399" />
                    <RANKING order="2" place="2" resultid="6917" />
                    <RANKING order="3" place="3" resultid="2356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1546" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1547" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9107" daytime="19:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9108" daytime="19:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1406" daytime="16:20" gender="M" number="21" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1407" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5950" />
                    <RANKING order="2" place="2" resultid="6338" />
                    <RANKING order="3" place="3" resultid="3255" />
                    <RANKING order="4" place="-1" resultid="4152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1408" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5106" />
                    <RANKING order="2" place="2" resultid="7367" />
                    <RANKING order="3" place="3" resultid="3171" />
                    <RANKING order="4" place="4" resultid="4166" />
                    <RANKING order="5" place="5" resultid="2073" />
                    <RANKING order="6" place="6" resultid="3496" />
                    <RANKING order="7" place="7" resultid="3852" />
                    <RANKING order="8" place="8" resultid="7027" />
                    <RANKING order="9" place="9" resultid="3892" />
                    <RANKING order="10" place="10" resultid="2132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1409" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2087" />
                    <RANKING order="2" place="2" resultid="3860" />
                    <RANKING order="3" place="3" resultid="3721" />
                    <RANKING order="4" place="4" resultid="6211" />
                    <RANKING order="5" place="5" resultid="6159" />
                    <RANKING order="6" place="6" resultid="2749" />
                    <RANKING order="7" place="-1" resultid="4766" />
                    <RANKING order="8" place="-1" resultid="4888" />
                    <RANKING order="9" place="-1" resultid="7061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6262" />
                    <RANKING order="2" place="2" resultid="3535" />
                    <RANKING order="3" place="3" resultid="2653" />
                    <RANKING order="4" place="4" resultid="3797" />
                    <RANKING order="5" place="5" resultid="2687" />
                    <RANKING order="6" place="6" resultid="4942" />
                    <RANKING order="7" place="7" resultid="3707" />
                    <RANKING order="8" place="8" resultid="3726" />
                    <RANKING order="9" place="9" resultid="7300" />
                    <RANKING order="10" place="10" resultid="2103" />
                    <RANKING order="11" place="11" resultid="3733" />
                    <RANKING order="12" place="12" resultid="4773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4957" />
                    <RANKING order="2" place="2" resultid="5712" />
                    <RANKING order="3" place="3" resultid="4234" />
                    <RANKING order="4" place="4" resultid="2730" />
                    <RANKING order="5" place="5" resultid="3937" />
                    <RANKING order="6" place="6" resultid="7375" />
                    <RANKING order="7" place="7" resultid="3424" />
                    <RANKING order="8" place="8" resultid="1897" />
                    <RANKING order="9" place="9" resultid="2430" />
                    <RANKING order="10" place="10" resultid="2419" />
                    <RANKING order="11" place="11" resultid="5775" />
                    <RANKING order="12" place="12" resultid="5880" />
                    <RANKING order="13" place="13" resultid="2813" />
                    <RANKING order="14" place="14" resultid="7049" />
                    <RANKING order="15" place="-1" resultid="3785" />
                    <RANKING order="16" place="-1" resultid="4948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1412" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2799" />
                    <RANKING order="2" place="2" resultid="4624" />
                    <RANKING order="3" place="3" resultid="3181" />
                    <RANKING order="4" place="4" resultid="2194" />
                    <RANKING order="5" place="5" resultid="4290" />
                    <RANKING order="6" place="6" resultid="3898" />
                    <RANKING order="7" place="7" resultid="3952" />
                    <RANKING order="8" place="8" resultid="5549" />
                    <RANKING order="9" place="9" resultid="1902" />
                    <RANKING order="10" place="-1" resultid="7313" />
                    <RANKING order="11" place="-1" resultid="7372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3887" />
                    <RANKING order="2" place="2" resultid="3393" />
                    <RANKING order="3" place="3" resultid="4808" />
                    <RANKING order="4" place="4" resultid="6864" />
                    <RANKING order="5" place="5" resultid="5095" />
                    <RANKING order="6" place="6" resultid="3385" />
                    <RANKING order="7" place="7" resultid="5680" />
                    <RANKING order="8" place="-1" resultid="3234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5100" />
                    <RANKING order="2" place="2" resultid="5865" />
                    <RANKING order="3" place="3" resultid="4668" />
                    <RANKING order="4" place="4" resultid="3569" />
                    <RANKING order="5" place="5" resultid="2325" />
                    <RANKING order="6" place="6" resultid="3992" />
                    <RANKING order="7" place="7" resultid="2302" />
                    <RANKING order="8" place="8" resultid="7390" />
                    <RANKING order="9" place="-1" resultid="2572" />
                    <RANKING order="10" place="-1" resultid="2982" />
                    <RANKING order="11" place="-1" resultid="3156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1415" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2186" />
                    <RANKING order="2" place="2" resultid="2940" />
                    <RANKING order="3" place="3" resultid="3017" />
                    <RANKING order="4" place="4" resultid="3563" />
                    <RANKING order="5" place="5" resultid="2635" />
                    <RANKING order="6" place="6" resultid="2579" />
                    <RANKING order="7" place="7" resultid="2592" />
                    <RANKING order="8" place="8" resultid="1978" />
                    <RANKING order="9" place="9" resultid="2387" />
                    <RANKING order="10" place="10" resultid="2288" />
                    <RANKING order="11" place="-1" resultid="5726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3489" />
                    <RANKING order="2" place="2" resultid="3023" />
                    <RANKING order="3" place="3" resultid="2481" />
                    <RANKING order="4" place="4" resultid="2276" />
                    <RANKING order="5" place="-1" resultid="5642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1417" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2316" />
                    <RANKING order="2" place="2" resultid="2955" />
                    <RANKING order="3" place="3" resultid="1993" />
                    <RANKING order="4" place="4" resultid="3328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1418" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6367" />
                    <RANKING order="2" place="2" resultid="2996" />
                    <RANKING order="3" place="3" resultid="3828" />
                    <RANKING order="4" place="4" resultid="5850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1420" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1421" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1422" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9043" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9044" daytime="16:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9045" daytime="16:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9046" daytime="16:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9047" daytime="16:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9048" daytime="16:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9049" daytime="16:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9050" daytime="16:40" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9051" daytime="16:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9052" daytime="16:45" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9053" daytime="16:50" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1388" daytime="16:00" gender="F" number="20" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1390" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2784" />
                    <RANKING order="2" place="2" resultid="7136" />
                    <RANKING order="3" place="3" resultid="1814" />
                    <RANKING order="4" place="4" resultid="3605" />
                    <RANKING order="5" place="5" resultid="4178" />
                    <RANKING order="6" place="6" resultid="2839" />
                    <RANKING order="7" place="7" resultid="4186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7130" />
                    <RANKING order="2" place="2" resultid="3811" />
                    <RANKING order="3" place="3" resultid="2511" />
                    <RANKING order="4" place="4" resultid="7006" />
                    <RANKING order="5" place="5" resultid="7168" />
                    <RANKING order="6" place="6" resultid="6031" />
                    <RANKING order="7" place="-1" resultid="7160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1392" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2519" />
                    <RANKING order="2" place="2" resultid="3867" />
                    <RANKING order="3" place="3" resultid="3683" />
                    <RANKING order="4" place="4" resultid="4965" />
                    <RANKING order="5" place="5" resultid="4815" />
                    <RANKING order="6" place="6" resultid="3751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1393" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2534" />
                    <RANKING order="2" place="2" resultid="4248" />
                    <RANKING order="3" place="3" resultid="4257" />
                    <RANKING order="4" place="4" resultid="6198" />
                    <RANKING order="5" place="5" resultid="5563" />
                    <RANKING order="6" place="6" resultid="2771" />
                    <RANKING order="7" place="7" resultid="3205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1394" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6394" />
                    <RANKING order="2" place="2" resultid="3542" />
                    <RANKING order="3" place="3" resultid="3926" />
                    <RANKING order="4" place="4" resultid="3458" />
                    <RANKING order="5" place="-1" resultid="2446" />
                    <RANKING order="6" place="-1" resultid="6013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1395" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7233" />
                    <RANKING order="2" place="2" resultid="5804" />
                    <RANKING order="3" place="3" resultid="4206" />
                    <RANKING order="4" place="4" resultid="2645" />
                    <RANKING order="5" place="5" resultid="5576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1396" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3971" />
                    <RANKING order="2" place="2" resultid="3523" />
                    <RANKING order="3" place="3" resultid="3404" />
                    <RANKING order="4" place="4" resultid="6870" />
                    <RANKING order="5" place="5" resultid="2347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6840" />
                    <RANKING order="2" place="2" resultid="7362" />
                    <RANKING order="3" place="3" resultid="5795" />
                    <RANKING order="4" place="4" resultid="3188" />
                    <RANKING order="5" place="5" resultid="2341" />
                    <RANKING order="6" place="6" resultid="6876" />
                    <RANKING order="7" place="7" resultid="2334" />
                    <RANKING order="8" place="-1" resultid="6025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3004" />
                    <RANKING order="2" place="2" resultid="3163" />
                    <RANKING order="3" place="3" resultid="6410" />
                    <RANKING order="4" place="4" resultid="2352" />
                    <RANKING order="5" place="5" resultid="3337" />
                    <RANKING order="6" place="6" resultid="6165" />
                    <RANKING order="7" place="7" resultid="1821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1399" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5664" />
                    <RANKING order="2" place="2" resultid="7293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1400" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1401" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1402" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1403" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1404" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1405" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9036" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9037" daytime="16:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9038" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9039" daytime="16:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9040" daytime="16:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9041" daytime="16:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9042" daytime="16:20" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1508" daytime="18:25" gender="M" number="27" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1509" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2259" />
                    <RANKING order="2" place="2" resultid="6907" />
                    <RANKING order="3" place="3" resultid="5636" />
                    <RANKING order="4" place="4" resultid="2859" />
                    <RANKING order="5" place="5" resultid="1805" />
                    <RANKING order="6" place="6" resultid="3358" />
                    <RANKING order="7" place="-1" resultid="6348" />
                    <RANKING order="8" place="-1" resultid="5082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2096" />
                    <RANKING order="2" place="2" resultid="3595" />
                    <RANKING order="3" place="3" resultid="5771" />
                    <RANKING order="4" place="4" resultid="6329" />
                    <RANKING order="5" place="5" resultid="2854" />
                    <RANKING order="6" place="6" resultid="2074" />
                    <RANKING order="7" place="7" resultid="4916" />
                    <RANKING order="8" place="8" resultid="4160" />
                    <RANKING order="9" place="9" resultid="2793" />
                    <RANKING order="10" place="10" resultid="7043" />
                    <RANKING order="11" place="11" resultid="2133" />
                    <RANKING order="12" place="-1" resultid="4167" />
                    <RANKING order="13" place="-1" resultid="4172" />
                    <RANKING order="14" place="-1" resultid="4219" />
                    <RANKING order="15" place="-1" resultid="5074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1511" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3714" />
                    <RANKING order="2" place="2" resultid="7092" />
                    <RANKING order="3" place="3" resultid="2145" />
                    <RANKING order="4" place="4" resultid="2475" />
                    <RANKING order="5" place="5" resultid="5900" />
                    <RANKING order="6" place="6" resultid="2848" />
                    <RANKING order="7" place="7" resultid="2543" />
                    <RANKING order="8" place="8" resultid="4202" />
                    <RANKING order="9" place="9" resultid="4889" />
                    <RANKING order="10" place="10" resultid="2550" />
                    <RANKING order="11" place="-1" resultid="5119" />
                    <RANKING order="12" place="-1" resultid="6891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1512" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6883" />
                    <RANKING order="2" place="2" resultid="5917" />
                    <RANKING order="3" place="3" resultid="3692" />
                    <RANKING order="4" place="4" resultid="2808" />
                    <RANKING order="5" place="5" resultid="3980" />
                    <RANKING order="6" place="6" resultid="2504" />
                    <RANKING order="7" place="7" resultid="3881" />
                    <RANKING order="8" place="8" resultid="6278" />
                    <RANKING order="9" place="9" resultid="4867" />
                    <RANKING order="10" place="10" resultid="6413" />
                    <RANKING order="11" place="11" resultid="3944" />
                    <RANKING order="12" place="12" resultid="4943" />
                    <RANKING order="13" place="13" resultid="2400" />
                    <RANKING order="14" place="-1" resultid="3745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1513" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2705" />
                    <RANKING order="2" place="2" resultid="4958" />
                    <RANKING order="3" place="3" resultid="6224" />
                    <RANKING order="4" place="4" resultid="3786" />
                    <RANKING order="5" place="5" resultid="4285" />
                    <RANKING order="6" place="6" resultid="4689" />
                    <RANKING order="7" place="7" resultid="1876" />
                    <RANKING order="8" place="8" resultid="7251" />
                    <RANKING order="9" place="9" resultid="6007" />
                    <RANKING order="10" place="10" resultid="3957" />
                    <RANKING order="11" place="11" resultid="1898" />
                    <RANKING order="12" place="12" resultid="4241" />
                    <RANKING order="13" place="13" resultid="6001" />
                    <RANKING order="14" place="14" resultid="5776" />
                    <RANKING order="15" place="15" resultid="6232" />
                    <RANKING order="16" place="16" resultid="3228" />
                    <RANKING order="17" place="-1" resultid="2268" />
                    <RANKING order="18" place="-1" resultid="3559" />
                    <RANKING order="19" place="-1" resultid="3907" />
                    <RANKING order="20" place="-1" resultid="5688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1514" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4823" />
                    <RANKING order="2" place="2" resultid="6134" />
                    <RANKING order="3" place="3" resultid="3837" />
                    <RANKING order="4" place="4" resultid="3398" />
                    <RANKING order="5" place="5" resultid="3449" />
                    <RANKING order="6" place="6" resultid="3182" />
                    <RANKING order="7" place="7" resultid="2057" />
                    <RANKING order="8" place="8" resultid="4078" />
                    <RANKING order="9" place="9" resultid="2948" />
                    <RANKING order="10" place="10" resultid="7314" />
                    <RANKING order="11" place="11" resultid="2012" />
                    <RANKING order="12" place="12" resultid="3899" />
                    <RANKING order="13" place="13" resultid="2417" />
                    <RANKING order="14" place="14" resultid="5550" />
                    <RANKING order="15" place="15" resultid="1903" />
                    <RANKING order="16" place="-1" resultid="2964" />
                    <RANKING order="17" place="-1" resultid="3353" />
                    <RANKING order="18" place="-1" resultid="9196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6900" />
                    <RANKING order="2" place="2" resultid="3453" />
                    <RANKING order="3" place="3" resultid="5933" />
                    <RANKING order="4" place="4" resultid="6238" />
                    <RANKING order="5" place="5" resultid="3342" />
                    <RANKING order="6" place="-1" resultid="6851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3793" />
                    <RANKING order="2" place="2" resultid="3505" />
                    <RANKING order="3" place="3" resultid="2408" />
                    <RANKING order="4" place="4" resultid="3373" />
                    <RANKING order="5" place="5" resultid="7344" />
                    <RANKING order="6" place="6" resultid="3874" />
                    <RANKING order="7" place="7" resultid="7330" />
                    <RANKING order="8" place="-1" resultid="3222" />
                    <RANKING order="9" place="-1" resultid="3481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3967" />
                    <RANKING order="2" place="2" resultid="1891" />
                    <RANKING order="3" place="3" resultid="5647" />
                    <RANKING order="4" place="4" resultid="3013" />
                    <RANKING order="5" place="5" resultid="2065" />
                    <RANKING order="6" place="6" resultid="2388" />
                    <RANKING order="7" place="7" resultid="3148" />
                    <RANKING order="8" place="8" resultid="2289" />
                    <RANKING order="9" place="-1" resultid="2636" />
                    <RANKING order="10" place="-1" resultid="2823" />
                    <RANKING order="11" place="-1" resultid="5858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1518" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3820" />
                    <RANKING order="2" place="2" resultid="7285" />
                    <RANKING order="3" place="3" resultid="1946" />
                    <RANKING order="4" place="4" resultid="2489" />
                    <RANKING order="5" place="5" resultid="2277" />
                    <RANKING order="6" place="-1" resultid="3610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1519" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1789" />
                    <RANKING order="2" place="2" resultid="3845" />
                    <RANKING order="3" place="3" resultid="3366" />
                    <RANKING order="4" place="4" resultid="1994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1520" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7227" />
                    <RANKING order="2" place="2" resultid="7337" />
                    <RANKING order="3" place="3" resultid="1987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1521" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1522" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1523" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1524" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9094" daytime="18:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9095" daytime="18:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9096" daytime="18:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9097" daytime="18:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9098" daytime="18:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9099" daytime="18:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9100" daytime="18:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9101" daytime="18:55" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9102" daytime="19:00" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9103" daytime="19:05" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9104" daytime="19:05" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="9105" daytime="19:10" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="9106" daytime="19:15" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1474" daytime="17:35" gender="M" number="25" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1475" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2382" />
                    <RANKING order="2" place="2" resultid="5544" />
                    <RANKING order="3" place="3" resultid="5535" />
                    <RANKING order="4" place="4" resultid="2121" />
                    <RANKING order="5" place="5" resultid="6347" />
                    <RANKING order="6" place="-1" resultid="4153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1476" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4838" />
                    <RANKING order="2" place="2" resultid="2853" />
                    <RANKING order="3" place="3" resultid="4915" />
                    <RANKING order="4" place="4" resultid="4218" />
                    <RANKING order="5" place="5" resultid="4880" />
                    <RANKING order="6" place="6" resultid="7146" />
                    <RANKING order="7" place="7" resultid="3853" />
                    <RANKING order="8" place="-1" resultid="1780" />
                    <RANKING order="9" place="-1" resultid="5976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1477" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7193" />
                    <RANKING order="2" place="2" resultid="3474" />
                    <RANKING order="3" place="3" resultid="6890" />
                    <RANKING order="4" place="4" resultid="7177" />
                    <RANKING order="5" place="5" resultid="3722" />
                    <RANKING order="6" place="6" resultid="5588" />
                    <RANKING order="7" place="7" resultid="3212" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1478" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4693" />
                    <RANKING order="2" place="2" resultid="2503" />
                    <RANKING order="3" place="3" resultid="2600" />
                    <RANKING order="4" place="4" resultid="3600" />
                    <RANKING order="5" place="5" resultid="6263" />
                    <RANKING order="6" place="6" resultid="5939" />
                    <RANKING order="7" place="7" resultid="2662" />
                    <RANKING order="8" place="8" resultid="2019" />
                    <RANKING order="9" place="9" resultid="6277" />
                    <RANKING order="10" place="-1" resultid="3536" />
                    <RANKING order="11" place="-1" resultid="3738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1479" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2672" />
                    <RANKING order="2" place="2" resultid="2427" />
                    <RANKING order="3" place="3" resultid="3558" />
                    <RANKING order="4" place="4" resultid="5966" />
                    <RANKING order="5" place="-1" resultid="4273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1480" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3920" />
                    <RANKING order="2" place="2" resultid="4831" />
                    <RANKING order="3" place="3" resultid="3836" />
                    <RANKING order="4" place="4" resultid="3448" />
                    <RANKING order="5" place="5" resultid="3410" />
                    <RANKING order="6" place="6" resultid="6858" />
                    <RANKING order="7" place="7" resultid="2056" />
                    <RANKING order="8" place="8" resultid="2195" />
                    <RANKING order="9" place="-1" resultid="4928" />
                    <RANKING order="10" place="-1" resultid="5820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7109" />
                    <RANKING order="2" place="2" resultid="4226" />
                    <RANKING order="3" place="3" resultid="5092" />
                    <RANKING order="4" place="4" resultid="7307" />
                    <RANKING order="5" place="5" resultid="3235" />
                    <RANKING order="6" place="-1" resultid="3588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5101" />
                    <RANKING order="2" place="2" resultid="2695" />
                    <RANKING order="3" place="3" resultid="6378" />
                    <RANKING order="4" place="4" resultid="2566" />
                    <RANKING order="5" place="5" resultid="2608" />
                    <RANKING order="6" place="6" resultid="3221" />
                    <RANKING order="7" place="7" resultid="3993" />
                    <RANKING order="8" place="8" resultid="7391" />
                    <RANKING order="9" place="-1" resultid="2303" />
                    <RANKING order="10" place="-1" resultid="2983" />
                    <RANKING order="11" place="-1" resultid="3504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4661" />
                    <RANKING order="2" place="2" resultid="2064" />
                    <RANKING order="3" place="3" resultid="1969" />
                    <RANKING order="4" place="4" resultid="4654" />
                    <RANKING order="5" place="5" resultid="2581" />
                    <RANKING order="6" place="6" resultid="2822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1484" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2679" />
                    <RANKING order="2" place="2" resultid="3819" />
                    <RANKING order="3" place="3" resultid="2036" />
                    <RANKING order="4" place="4" resultid="6356" />
                    <RANKING order="5" place="5" resultid="2626" />
                    <RANKING order="6" place="6" resultid="2309" />
                    <RANKING order="7" place="7" resultid="7322" />
                    <RANKING order="8" place="-1" resultid="2482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1485" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4648" />
                    <RANKING order="2" place="2" resultid="3844" />
                    <RANKING order="3" place="3" resultid="7265" />
                    <RANKING order="4" place="4" resultid="3329" />
                    <RANKING order="5" place="-1" resultid="2956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1486" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7101" />
                    <RANKING order="2" place="2" resultid="5851" />
                    <RANKING order="3" place="3" resultid="3041" />
                    <RANKING order="4" place="4" resultid="1986" />
                    <RANKING order="5" place="5" resultid="2296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1487" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1488" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1489" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1490" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9079" daytime="17:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9080" daytime="17:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9081" daytime="17:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9082" daytime="17:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9083" daytime="17:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9084" daytime="17:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9085" daytime="17:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9086" daytime="17:55" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9087" daytime="17:55" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1423" daytime="16:50" gender="F" number="22" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1424" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5627" />
                    <RANKING order="2" place="2" resultid="7137" />
                    <RANKING order="3" place="3" resultid="7020" />
                    <RANKING order="4" place="4" resultid="2126" />
                    <RANKING order="5" place="5" resultid="4187" />
                    <RANKING order="6" place="6" resultid="7033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7220" />
                    <RANKING order="2" place="2" resultid="4873" />
                    <RANKING order="3" place="3" resultid="3575" />
                    <RANKING order="4" place="4" resultid="4724" />
                    <RANKING order="5" place="5" resultid="1940" />
                    <RANKING order="6" place="6" resultid="3432" />
                    <RANKING order="7" place="7" resultid="6245" />
                    <RANKING order="8" place="8" resultid="5971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3986" />
                    <RANKING order="2" place="2" resultid="3442" />
                    <RANKING order="3" place="3" resultid="6190" />
                    <RANKING order="4" place="4" resultid="3437" />
                    <RANKING order="5" place="5" resultid="4966" />
                    <RANKING order="6" place="6" resultid="4022" />
                    <RANKING order="7" place="7" resultid="5906" />
                    <RANKING order="8" place="8" resultid="5557" />
                    <RANKING order="9" place="9" resultid="4792" />
                    <RANKING order="10" place="10" resultid="4018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6199" />
                    <RANKING order="2" place="2" resultid="6253" />
                    <RANKING order="3" place="3" resultid="2468" />
                    <RANKING order="4" place="4" resultid="4755" />
                    <RANKING order="5" place="5" resultid="4265" />
                    <RANKING order="6" place="6" resultid="5673" />
                    <RANKING order="7" place="7" resultid="2736" />
                    <RANKING order="8" place="8" resultid="4258" />
                    <RANKING order="9" place="9" resultid="4854" />
                    <RANKING order="10" place="-1" resultid="6408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3543" />
                    <RANKING order="2" place="2" resultid="7257" />
                    <RANKING order="3" place="3" resultid="2447" />
                    <RANKING order="4" place="4" resultid="7379" />
                    <RANKING order="5" place="5" resultid="4800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7234" />
                    <RANKING order="2" place="2" resultid="7245" />
                    <RANKING order="3" place="3" resultid="5595" />
                    <RANKING order="4" place="4" resultid="5870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3529" />
                    <RANKING order="2" place="2" resultid="3405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1431" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6841" />
                    <RANKING order="2" place="2" resultid="7275" />
                    <RANKING order="3" place="3" resultid="2392" />
                    <RANKING order="4" place="4" resultid="4640" />
                    <RANKING order="5" place="-1" resultid="5676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1432" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3005" />
                    <RANKING order="2" place="2" resultid="3620" />
                    <RANKING order="3" place="3" resultid="3032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4633" />
                    <RANKING order="2" place="2" resultid="3932" />
                    <RANKING order="3" place="3" resultid="7294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1435" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1436" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1437" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1438" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1439" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9054" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9055" daytime="16:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9056" daytime="16:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9057" daytime="16:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9058" daytime="17:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9059" daytime="17:00" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1491" daytime="18:00" gender="F" number="26" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1492" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2785" />
                    <RANKING order="2" place="2" resultid="5628" />
                    <RANKING order="3" place="3" resultid="4179" />
                    <RANKING order="4" place="4" resultid="3606" />
                    <RANKING order="5" place="5" resultid="1815" />
                    <RANKING order="6" place="6" resultid="6896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4874" />
                    <RANKING order="2" place="2" resultid="3418" />
                    <RANKING order="3" place="3" resultid="5911" />
                    <RANKING order="4" place="4" resultid="3948" />
                    <RANKING order="5" place="5" resultid="2082" />
                    <RANKING order="6" place="6" resultid="5787" />
                    <RANKING order="7" place="7" resultid="6141" />
                    <RANKING order="8" place="-1" resultid="5657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3443" />
                    <RANKING order="2" place="2" resultid="2765" />
                    <RANKING order="3" place="3" resultid="6217" />
                    <RANKING order="4" place="4" resultid="4816" />
                    <RANKING order="5" place="5" resultid="6205" />
                    <RANKING order="6" place="6" resultid="4023" />
                    <RANKING order="7" place="7" resultid="5907" />
                    <RANKING order="8" place="8" resultid="4793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1495" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1952" />
                    <RANKING order="2" place="2" resultid="4756" />
                    <RANKING order="3" place="3" resultid="5564" />
                    <RANKING order="4" place="4" resultid="2772" />
                    <RANKING order="5" place="5" resultid="3206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1496" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6395" />
                    <RANKING order="2" place="2" resultid="2150" />
                    <RANKING order="3" place="3" resultid="2777" />
                    <RANKING order="4" place="4" resultid="2617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1497" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7246" />
                    <RANKING order="2" place="2" resultid="3138" />
                    <RANKING order="3" place="3" resultid="6285" />
                    <RANKING order="4" place="4" resultid="7349" />
                    <RANKING order="5" place="5" resultid="4207" />
                    <RANKING order="6" place="6" resultid="2456" />
                    <RANKING order="7" place="7" resultid="5577" />
                    <RANKING order="8" place="-1" resultid="5670" />
                    <RANKING order="9" place="-1" resultid="5871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1498" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3972" />
                    <RANKING order="2" place="2" resultid="6846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1499" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7276" />
                    <RANKING order="2" place="2" resultid="3198" />
                    <RANKING order="3" place="3" resultid="5796" />
                    <RANKING order="4" place="4" resultid="2244" />
                    <RANKING order="5" place="5" resultid="2335" />
                    <RANKING order="6" place="-1" resultid="2342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1500" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6404" />
                    <RANKING order="2" place="2" resultid="4006" />
                    <RANKING order="3" place="3" resultid="2003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1502" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1503" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1504" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1505" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1506" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1507" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9088" daytime="18:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9089" daytime="18:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9090" daytime="18:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9091" daytime="18:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9092" daytime="18:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9093" daytime="18:25" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2015-11-15" daytime="09:00" name="BLOK IV" number="4" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1681" daytime="11:00" gender="M" number="37" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1682" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5951" />
                    <RANKING order="2" place="2" resultid="2123" />
                    <RANKING order="3" place="3" resultid="5537" />
                    <RANKING order="4" place="4" resultid="3257" />
                    <RANKING order="5" place="-1" resultid="4155" />
                    <RANKING order="6" place="-1" resultid="6184" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1683" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7369" />
                    <RANKING order="2" place="2" resultid="3173" />
                    <RANKING order="3" place="3" resultid="3498" />
                    <RANKING order="4" place="4" resultid="2075" />
                    <RANKING order="5" place="5" resultid="3854" />
                    <RANKING order="6" place="6" resultid="4840" />
                    <RANKING order="7" place="7" resultid="7028" />
                    <RANKING order="8" place="8" resultid="3893" />
                    <RANKING order="9" place="9" resultid="1936" />
                    <RANKING order="10" place="10" resultid="2134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1684" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2116" />
                    <RANKING order="2" place="2" resultid="2088" />
                    <RANKING order="3" place="3" resultid="5982" />
                    <RANKING order="4" place="4" resultid="3862" />
                    <RANKING order="5" place="5" resultid="7186" />
                    <RANKING order="6" place="6" resultid="6160" />
                    <RANKING order="7" place="7" resultid="4782" />
                    <RANKING order="8" place="8" resultid="6214" />
                    <RANKING order="9" place="9" resultid="2751" />
                    <RANKING order="10" place="10" resultid="4953" />
                    <RANKING order="11" place="-1" resultid="4768" />
                    <RANKING order="12" place="-1" resultid="4890" />
                    <RANKING order="13" place="-1" resultid="7062" />
                    <RANKING order="14" place="-1" resultid="7179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1685" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4013" />
                    <RANKING order="2" place="2" resultid="6885" />
                    <RANKING order="3" place="3" resultid="3709" />
                    <RANKING order="4" place="4" resultid="3601" />
                    <RANKING order="5" place="5" resultid="3538" />
                    <RANKING order="6" place="6" resultid="3799" />
                    <RANKING order="7" place="7" resultid="3759" />
                    <RANKING order="8" place="8" resultid="5946" />
                    <RANKING order="9" place="9" resultid="7384" />
                    <RANKING order="10" place="10" resultid="2689" />
                    <RANKING order="11" place="11" resultid="3697" />
                    <RANKING order="12" place="12" resultid="4868" />
                    <RANKING order="13" place="13" resultid="3727" />
                    <RANKING order="14" place="14" resultid="7301" />
                    <RANKING order="15" place="15" resultid="3739" />
                    <RANKING order="16" place="16" resultid="2104" />
                    <RANKING order="17" place="17" resultid="1925" />
                    <RANKING order="18" place="18" resultid="3734" />
                    <RANKING order="19" place="-1" resultid="6264" />
                    <RANKING order="20" place="-1" resultid="2021" />
                    <RANKING order="21" place="-1" resultid="4775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1686" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4959" />
                    <RANKING order="2" place="2" resultid="2707" />
                    <RANKING order="3" place="3" resultid="5714" />
                    <RANKING order="4" place="4" resultid="4287" />
                    <RANKING order="5" place="5" resultid="3938" />
                    <RANKING order="6" place="6" resultid="4236" />
                    <RANKING order="7" place="7" resultid="2731" />
                    <RANKING order="8" place="8" resultid="4278" />
                    <RANKING order="9" place="9" resultid="2674" />
                    <RANKING order="10" place="10" resultid="3426" />
                    <RANKING order="11" place="11" resultid="7376" />
                    <RANKING order="12" place="12" resultid="2431" />
                    <RANKING order="13" place="13" resultid="2816" />
                    <RANKING order="14" place="14" resultid="2420" />
                    <RANKING order="15" place="15" resultid="5881" />
                    <RANKING order="16" place="16" resultid="7050" />
                    <RANKING order="17" place="17" resultid="6233" />
                    <RANKING order="18" place="-1" resultid="4788" />
                    <RANKING order="19" place="-1" resultid="2270" />
                    <RANKING order="20" place="-1" resultid="4949" />
                    <RANKING order="21" place="-1" resultid="6003" />
                    <RANKING order="22" place="-1" resultid="6353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1687" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2801" />
                    <RANKING order="2" place="2" resultid="4626" />
                    <RANKING order="3" place="3" resultid="3900" />
                    <RANKING order="4" place="4" resultid="6292" />
                    <RANKING order="5" place="5" resultid="2197" />
                    <RANKING order="6" place="6" resultid="7315" />
                    <RANKING order="7" place="7" resultid="3954" />
                    <RANKING order="8" place="8" resultid="5551" />
                    <RANKING order="9" place="9" resultid="2014" />
                    <RANKING order="10" place="10" resultid="2966" />
                    <RANKING order="11" place="-1" resultid="4292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1688" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3889" />
                    <RANKING order="2" place="2" resultid="3394" />
                    <RANKING order="3" place="3" resultid="6155" />
                    <RANKING order="4" place="4" resultid="7309" />
                    <RANKING order="5" place="5" resultid="6865" />
                    <RANKING order="6" place="6" resultid="5681" />
                    <RANKING order="7" place="7" resultid="3582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1689" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3794" />
                    <RANKING order="2" place="2" resultid="5866" />
                    <RANKING order="3" place="3" resultid="3570" />
                    <RANKING order="4" place="4" resultid="7119" />
                    <RANKING order="5" place="5" resultid="2327" />
                    <RANKING order="6" place="6" resultid="2574" />
                    <RANKING order="7" place="7" resultid="2304" />
                    <RANKING order="8" place="-1" resultid="3159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1690" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2942" />
                    <RANKING order="2" place="2" resultid="2189" />
                    <RANKING order="3" place="3" resultid="3018" />
                    <RANKING order="4" place="4" resultid="3565" />
                    <RANKING order="5" place="5" resultid="4664" />
                    <RANKING order="6" place="6" resultid="2595" />
                    <RANKING order="7" place="7" resultid="2637" />
                    <RANKING order="8" place="8" resultid="2582" />
                    <RANKING order="9" place="9" resultid="2529" />
                    <RANKING order="10" place="10" resultid="1980" />
                    <RANKING order="11" place="11" resultid="2290" />
                    <RANKING order="12" place="-1" resultid="1909" />
                    <RANKING order="13" place="-1" resultid="5727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1691" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3490" />
                    <RANKING order="2" place="2" resultid="3026" />
                    <RANKING order="3" place="3" resultid="2483" />
                    <RANKING order="4" place="4" resultid="2311" />
                    <RANKING order="5" place="5" resultid="2279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1692" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1791" />
                    <RANKING order="2" place="2" resultid="2319" />
                    <RANKING order="3" place="3" resultid="4650" />
                    <RANKING order="4" place="4" resultid="2958" />
                    <RANKING order="5" place="5" resultid="3846" />
                    <RANKING order="6" place="6" resultid="1996" />
                    <RANKING order="7" place="7" resultid="3331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1693" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6368" />
                    <RANKING order="2" place="2" resultid="2999" />
                    <RANKING order="3" place="3" resultid="1963" />
                    <RANKING order="4" place="4" resultid="3831" />
                    <RANKING order="5" place="5" resultid="7338" />
                    <RANKING order="6" place="6" resultid="2500" />
                    <RANKING order="7" place="7" resultid="2297" />
                    <RANKING order="8" place="-1" resultid="5852" />
                    <RANKING order="9" place="-1" resultid="7103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1694" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5738" />
                    <RANKING order="2" place="2" resultid="5759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1695" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2833" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1696" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1697" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9159" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9160" daytime="11:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9161" daytime="11:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9162" daytime="11:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9163" daytime="11:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9164" daytime="11:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9165" daytime="11:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9166" daytime="11:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9167" daytime="11:15" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9168" daytime="11:15" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9169" daytime="11:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="9170" daytime="11:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="9171" daytime="11:20" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="9172" daytime="11:20" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1721" daytime="11:35" gender="F" number="39" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1728" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7057" />
                    <RANKING order="2" place="2" resultid="4181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1729" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3380" />
                    <RANKING order="2" place="2" resultid="2237" />
                    <RANKING order="3" place="3" resultid="3420" />
                    <RANKING order="4" place="4" resultid="4848" />
                    <RANKING order="5" place="5" resultid="2514" />
                    <RANKING order="6" place="6" resultid="5789" />
                    <RANKING order="7" place="7" resultid="6142" />
                    <RANKING order="8" place="8" resultid="5783" />
                    <RANKING order="9" place="-1" resultid="5620" />
                    <RANKING order="10" place="-1" resultid="5658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1730" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2767" />
                    <RANKING order="2" place="2" resultid="6218" />
                    <RANKING order="3" place="3" resultid="6207" />
                    <RANKING order="4" place="4" resultid="4817" />
                    <RANKING order="5" place="5" resultid="5558" />
                    <RANKING order="6" place="-1" resultid="4974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1731" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1953" />
                    <RANKING order="2" place="2" resultid="4251" />
                    <RANKING order="3" place="3" resultid="5566" />
                    <RANKING order="4" place="4" resultid="6295" />
                    <RANKING order="5" place="5" resultid="4856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1732" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6396" />
                    <RANKING order="2" place="2" resultid="4213" />
                    <RANKING order="3" place="3" resultid="2151" />
                    <RANKING order="4" place="4" resultid="2619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1733" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3139" />
                    <RANKING order="2" place="2" resultid="6287" />
                    <RANKING order="3" place="3" resultid="2458" />
                    <RANKING order="4" place="4" resultid="5579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1734" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3974" />
                    <RANKING order="2" place="2" resultid="6847" />
                    <RANKING order="3" place="3" resultid="6148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1735" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3470" />
                    <RANKING order="2" place="2" resultid="7278" />
                    <RANKING order="3" place="3" resultid="6027" />
                    <RANKING order="4" place="4" resultid="3200" />
                    <RANKING order="5" place="5" resultid="2247" />
                    <RANKING order="6" place="6" resultid="2337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1736" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6167" />
                    <RANKING order="2" place="2" resultid="1824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1737" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4636" />
                    <RANKING order="2" place="2" resultid="4007" />
                    <RANKING order="3" place="3" resultid="2005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1738" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1739" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1740" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1741" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1742" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1743" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9177" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9178" daytime="11:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9179" daytime="12:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9180" daytime="12:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9181" daytime="12:15" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1647" daytime="10:00" gender="M" number="35" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1648" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2383" />
                    <RANKING order="2" place="2" resultid="6349" />
                    <RANKING order="3" place="-1" resultid="4154" />
                    <RANKING order="4" place="-1" resultid="5638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1649" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4839" />
                    <RANKING order="2" place="2" resultid="2855" />
                    <RANKING order="3" place="3" resultid="4220" />
                    <RANKING order="4" place="4" resultid="4882" />
                    <RANKING order="5" place="5" resultid="7148" />
                    <RANKING order="6" place="-1" resultid="4174" />
                    <RANKING order="7" place="-1" resultid="5977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7094" />
                    <RANKING order="2" place="2" resultid="7195" />
                    <RANKING order="3" place="3" resultid="6892" />
                    <RANKING order="4" place="4" resultid="7178" />
                    <RANKING order="5" place="5" resultid="3723" />
                    <RANKING order="6" place="6" resultid="5589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4695" />
                    <RANKING order="2" place="2" resultid="2505" />
                    <RANKING order="3" place="3" resultid="5940" />
                    <RANKING order="4" place="4" resultid="6279" />
                    <RANKING order="5" place="5" resultid="2664" />
                    <RANKING order="6" place="-1" resultid="2020" />
                    <RANKING order="7" place="-1" resultid="2601" />
                    <RANKING order="8" place="-1" resultid="3537" />
                    <RANKING order="9" place="-1" resultid="2656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2673" />
                    <RANKING order="2" place="2" resultid="2428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1653" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4833" />
                    <RANKING order="2" place="2" resultid="3838" />
                    <RANKING order="3" place="3" resultid="3450" />
                    <RANKING order="4" place="4" resultid="3413" />
                    <RANKING order="5" place="5" resultid="6859" />
                    <RANKING order="6" place="6" resultid="2196" />
                    <RANKING order="7" place="7" resultid="5822" />
                    <RANKING order="8" place="8" resultid="2463" />
                    <RANKING order="9" place="9" resultid="2965" />
                    <RANKING order="10" place="10" resultid="2950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1654" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7110" />
                    <RANKING order="2" place="2" resultid="4227" />
                    <RANKING order="3" place="3" resultid="2050" />
                    <RANKING order="4" place="4" resultid="3591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1655" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2697" />
                    <RANKING order="2" place="2" resultid="2985" />
                    <RANKING order="3" place="3" resultid="6379" />
                    <RANKING order="4" place="4" resultid="2609" />
                    <RANKING order="5" place="5" resultid="2567" />
                    <RANKING order="6" place="6" resultid="4670" />
                    <RANKING order="7" place="7" resultid="2587" />
                    <RANKING order="8" place="8" resultid="3994" />
                    <RANKING order="9" place="9" resultid="7392" />
                    <RANKING order="10" place="-1" resultid="3158" />
                    <RANKING order="11" place="-1" resultid="3506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1656" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3968" />
                    <RANKING order="2" place="2" resultid="4663" />
                    <RANKING order="3" place="3" resultid="1972" />
                    <RANKING order="4" place="4" resultid="4655" />
                    <RANKING order="5" place="5" resultid="2824" />
                    <RANKING order="6" place="6" resultid="3149" />
                    <RANKING order="7" place="-1" resultid="5709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1657" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2681" />
                    <RANKING order="2" place="2" resultid="3821" />
                    <RANKING order="3" place="3" resultid="2037" />
                    <RANKING order="4" place="4" resultid="6357" />
                    <RANKING order="5" place="5" resultid="2629" />
                    <RANKING order="6" place="6" resultid="2310" />
                    <RANKING order="7" place="7" resultid="7323" />
                    <RANKING order="8" place="8" resultid="2278" />
                    <RANKING order="9" place="9" resultid="2492" />
                    <RANKING order="10" place="-1" resultid="5643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1658" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4649" />
                    <RANKING order="2" place="2" resultid="3367" />
                    <RANKING order="3" place="3" resultid="1995" />
                    <RANKING order="4" place="4" resultid="1886" />
                    <RANKING order="5" place="5" resultid="3330" />
                    <RANKING order="6" place="-1" resultid="2957" />
                    <RANKING order="7" place="-1" resultid="7266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1659" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3830" />
                    <RANKING order="2" place="2" resultid="2497" />
                    <RANKING order="3" place="3" resultid="1988" />
                    <RANKING order="4" place="-1" resultid="7102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1660" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1661" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1662" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1663" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9142" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9143" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9144" daytime="10:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9145" daytime="10:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9146" daytime="10:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9147" daytime="10:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9148" daytime="10:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9149" daytime="10:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9150" daytime="10:40" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1613" daytime="09:15" gender="M" number="33" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1614" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5877" />
                    <RANKING order="2" place="2" resultid="6909" />
                    <RANKING order="3" place="3" resultid="5637" />
                    <RANKING order="4" place="4" resultid="1807" />
                    <RANKING order="5" place="5" resultid="5536" />
                    <RANKING order="6" place="6" resultid="2122" />
                    <RANKING order="7" place="-1" resultid="5083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1615" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2097" />
                    <RANKING order="2" place="2" resultid="4685" />
                    <RANKING order="3" place="3" resultid="2140" />
                    <RANKING order="4" place="4" resultid="6330" />
                    <RANKING order="5" place="5" resultid="7044" />
                    <RANKING order="6" place="6" resultid="2205" />
                    <RANKING order="7" place="7" resultid="7147" />
                    <RANKING order="8" place="-1" resultid="3596" />
                    <RANKING order="9" place="-1" resultid="4707" />
                    <RANKING order="10" place="-1" resultid="5075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1616" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3715" />
                    <RANKING order="2" place="2" resultid="2115" />
                    <RANKING order="3" place="3" resultid="7194" />
                    <RANKING order="4" place="4" resultid="7185" />
                    <RANKING order="5" place="5" resultid="5120" />
                    <RANKING order="6" place="6" resultid="5901" />
                    <RANKING order="7" place="7" resultid="2545" />
                    <RANKING order="8" place="8" resultid="6213" />
                    <RANKING order="9" place="9" resultid="5583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1617" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4694" />
                    <RANKING order="2" place="2" resultid="5918" />
                    <RANKING order="3" place="3" resultid="2809" />
                    <RANKING order="4" place="4" resultid="3703" />
                    <RANKING order="5" place="5" resultid="4898" />
                    <RANKING order="6" place="6" resultid="5721" />
                    <RANKING order="7" place="7" resultid="2655" />
                    <RANKING order="8" place="8" resultid="2401" />
                    <RANKING order="9" place="9" resultid="5812" />
                    <RANKING order="10" place="-1" resultid="2109" />
                    <RANKING order="11" place="-1" resultid="2156" />
                    <RANKING order="12" place="-1" resultid="2688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2706" />
                    <RANKING order="2" place="2" resultid="6226" />
                    <RANKING order="3" place="3" resultid="5732" />
                    <RANKING order="4" place="4" resultid="1877" />
                    <RANKING order="5" place="5" resultid="4286" />
                    <RANKING order="6" place="6" resultid="7269" />
                    <RANKING order="7" place="7" resultid="2213" />
                    <RANKING order="8" place="8" resultid="2269" />
                    <RANKING order="9" place="9" resultid="4980" />
                    <RANKING order="10" place="10" resultid="6180" />
                    <RANKING order="11" place="-1" resultid="2815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3921" />
                    <RANKING order="2" place="2" resultid="6135" />
                    <RANKING order="3" place="3" resultid="3412" />
                    <RANKING order="4" place="4" resultid="5821" />
                    <RANKING order="5" place="5" resultid="2013" />
                    <RANKING order="6" place="6" resultid="2949" />
                    <RANKING order="7" place="7" resultid="3953" />
                    <RANKING order="8" place="-1" resultid="2868" />
                    <RANKING order="9" place="-1" resultid="4832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1620" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2049" />
                    <RANKING order="2" place="2" resultid="7308" />
                    <RANKING order="3" place="3" resultid="5935" />
                    <RANKING order="4" place="4" resultid="6835" />
                    <RANKING order="5" place="5" resultid="4810" />
                    <RANKING order="6" place="-1" resultid="3387" />
                    <RANKING order="7" place="-1" resultid="3590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1621" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6270" />
                    <RANKING order="2" place="2" resultid="5886" />
                    <RANKING order="3" place="3" resultid="3483" />
                    <RANKING order="4" place="4" resultid="7331" />
                    <RANKING order="5" place="-1" resultid="2410" />
                    <RANKING order="6" place="-1" resultid="2984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1622" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2188" />
                    <RANKING order="2" place="2" resultid="1971" />
                    <RANKING order="3" place="3" resultid="5859" />
                    <RANKING order="4" place="4" resultid="2066" />
                    <RANKING order="5" place="5" resultid="2594" />
                    <RANKING order="6" place="6" resultid="2528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1623" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1930" />
                    <RANKING order="2" place="2" resultid="1918" />
                    <RANKING order="3" place="3" resultid="3514" />
                    <RANKING order="4" place="4" resultid="7286" />
                    <RANKING order="5" place="5" resultid="2628" />
                    <RANKING order="6" place="6" resultid="2491" />
                    <RANKING order="7" place="-1" resultid="3025" />
                    <RANKING order="8" place="-1" resultid="5701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1624" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1790" />
                    <RANKING order="2" place="2" resultid="2318" />
                    <RANKING order="3" place="-1" resultid="1885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1625" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2998" />
                    <RANKING order="2" place="2" resultid="1962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1626" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1627" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1628" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1629" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9128" daytime="09:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9129" daytime="09:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9130" daytime="09:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9131" daytime="09:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9132" daytime="09:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9133" daytime="09:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9134" daytime="09:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9135" daytime="09:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9136" daytime="09:35" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9137" daytime="09:35" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1744" daytime="12:20" gender="M" number="40" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1745" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6910" />
                    <RANKING order="2" place="2" resultid="2860" />
                    <RANKING order="3" place="3" resultid="1808" />
                    <RANKING order="4" place="-1" resultid="3258" />
                    <RANKING order="5" place="-1" resultid="3359" />
                    <RANKING order="6" place="-1" resultid="5084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1746" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2098" />
                    <RANKING order="2" place="2" resultid="4221" />
                    <RANKING order="3" place="3" resultid="4911" />
                    <RANKING order="4" place="4" resultid="4162" />
                    <RANKING order="5" place="5" resultid="7045" />
                    <RANKING order="6" place="6" resultid="2135" />
                    <RANKING order="7" place="-1" resultid="2076" />
                    <RANKING order="8" place="-1" resultid="2206" />
                    <RANKING order="9" place="-1" resultid="3174" />
                    <RANKING order="10" place="-1" resultid="6331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1747" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7095" />
                    <RANKING order="2" place="2" resultid="3863" />
                    <RANKING order="3" place="3" resultid="5902" />
                    <RANKING order="4" place="4" resultid="4891" />
                    <RANKING order="5" place="5" resultid="3213" />
                    <RANKING order="6" place="6" resultid="2551" />
                    <RANKING order="7" place="-1" resultid="2146" />
                    <RANKING order="8" place="-1" resultid="2546" />
                    <RANKING order="9" place="-1" resultid="6893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1748" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6886" />
                    <RANKING order="2" place="2" resultid="3693" />
                    <RANKING order="3" place="3" resultid="5722" />
                    <RANKING order="4" place="4" resultid="3981" />
                    <RANKING order="5" place="5" resultid="3882" />
                    <RANKING order="6" place="6" resultid="2665" />
                    <RANKING order="7" place="7" resultid="3746" />
                    <RANKING order="8" place="8" resultid="3945" />
                    <RANKING order="9" place="9" resultid="2110" />
                    <RANKING order="10" place="10" resultid="6414" />
                    <RANKING order="11" place="11" resultid="7385" />
                    <RANKING order="12" place="12" resultid="5813" />
                    <RANKING order="13" place="13" resultid="2402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1749" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6227" />
                    <RANKING order="2" place="2" resultid="3787" />
                    <RANKING order="3" place="3" resultid="3908" />
                    <RANKING order="4" place="4" resultid="7252" />
                    <RANKING order="5" place="5" resultid="6008" />
                    <RANKING order="6" place="6" resultid="4243" />
                    <RANKING order="7" place="7" resultid="6234" />
                    <RANKING order="8" place="8" resultid="3229" />
                    <RANKING order="9" place="-1" resultid="2214" />
                    <RANKING order="10" place="-1" resultid="4960" />
                    <RANKING order="11" place="-1" resultid="4981" />
                    <RANKING order="12" place="-1" resultid="5689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1750" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6136" />
                    <RANKING order="2" place="2" resultid="3354" />
                    <RANKING order="3" place="3" resultid="4825" />
                    <RANKING order="4" place="4" resultid="3399" />
                    <RANKING order="5" place="5" resultid="2058" />
                    <RANKING order="6" place="6" resultid="3451" />
                    <RANKING order="7" place="7" resultid="9197" />
                    <RANKING order="8" place="-1" resultid="2464" />
                    <RANKING order="9" place="-1" resultid="4627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1751" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3454" />
                    <RANKING order="2" place="2" resultid="6901" />
                    <RANKING order="3" place="3" resultid="8884" />
                    <RANKING order="4" place="4" resultid="6156" />
                    <RANKING order="5" place="5" resultid="5936" />
                    <RANKING order="6" place="6" resultid="6240" />
                    <RANKING order="7" place="7" resultid="6836" />
                    <RANKING order="8" place="-1" resultid="3343" />
                    <RANKING order="9" place="-1" resultid="3388" />
                    <RANKING order="10" place="-1" resultid="3395" />
                    <RANKING order="11" place="-1" resultid="6853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1752" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6271" />
                    <RANKING order="2" place="2" resultid="3507" />
                    <RANKING order="3" place="3" resultid="2411" />
                    <RANKING order="4" place="4" resultid="3484" />
                    <RANKING order="5" place="5" resultid="7345" />
                    <RANKING order="6" place="6" resultid="3374" />
                    <RANKING order="7" place="7" resultid="3875" />
                    <RANKING order="8" place="8" resultid="2613" />
                    <RANKING order="9" place="9" resultid="3995" />
                    <RANKING order="10" place="10" resultid="3223" />
                    <RANKING order="11" place="11" resultid="7332" />
                    <RANKING order="12" place="12" resultid="2328" />
                    <RANKING order="13" place="-1" resultid="2568" />
                    <RANKING order="14" place="-1" resultid="2698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1753" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5648" />
                    <RANKING order="2" place="2" resultid="3014" />
                    <RANKING order="3" place="3" resultid="5860" />
                    <RANKING order="4" place="4" resultid="2067" />
                    <RANKING order="5" place="5" resultid="2389" />
                    <RANKING order="6" place="6" resultid="1981" />
                    <RANKING order="7" place="7" resultid="3150" />
                    <RANKING order="8" place="-1" resultid="1910" />
                    <RANKING order="9" place="-1" resultid="2291" />
                    <RANKING order="10" place="-1" resultid="2638" />
                    <RANKING order="11" place="-1" resultid="2825" />
                    <RANKING order="12" place="-1" resultid="4656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1754" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3822" />
                    <RANKING order="2" place="2" resultid="2682" />
                    <RANKING order="3" place="3" resultid="1919" />
                    <RANKING order="4" place="4" resultid="7287" />
                    <RANKING order="5" place="5" resultid="3611" />
                    <RANKING order="6" place="-1" resultid="1947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1755" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3368" />
                    <RANKING order="2" place="2" resultid="3847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1756" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6384" />
                    <RANKING order="2" place="2" resultid="7339" />
                    <RANKING order="3" place="-1" resultid="7228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1757" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1758" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1759" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1760" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9182" daytime="12:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9183" daytime="12:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9184" daytime="12:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9185" daytime="12:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9186" daytime="12:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9187" daytime="13:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9188" daytime="13:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9189" daytime="13:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9190" daytime="13:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9191" daytime="13:30" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9192" daytime="13:35" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1698" daytime="11:20" gender="X" number="38" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1715" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7524" />
                    <RANKING order="2" place="2" resultid="8601" />
                    <RANKING order="3" place="-1" resultid="7070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1716" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3624" />
                    <RANKING order="2" place="2" resultid="2555" />
                    <RANKING order="3" place="3" resultid="6298" />
                    <RANKING order="4" place="4" resultid="2870" />
                    <RANKING order="5" place="5" resultid="2753" />
                    <RANKING order="6" place="6" resultid="5953" />
                    <RANKING order="7" place="7" resultid="7066" />
                    <RANKING order="8" place="8" resultid="8603" />
                    <RANKING order="9" place="9" resultid="6307" />
                    <RANKING order="10" place="-1" resultid="5600" />
                    <RANKING order="11" place="-1" resultid="4802" />
                    <RANKING order="12" place="-1" resultid="5829" />
                    <RANKING order="13" place="-1" resultid="7526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1717" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8600" />
                    <RANKING order="2" place="2" resultid="7394" />
                    <RANKING order="3" place="3" resultid="4294" />
                    <RANKING order="4" place="4" resultid="6915" />
                    <RANKING order="5" place="5" resultid="3427" />
                    <RANKING order="6" place="6" resultid="6305" />
                    <RANKING order="7" place="7" resultid="4930" />
                    <RANKING order="8" place="8" resultid="6034" />
                    <RANKING order="9" place="9" resultid="5830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1718" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7396" />
                    <RANKING order="2" place="2" resultid="3242" />
                    <RANKING order="3" place="3" resultid="6916" />
                    <RANKING order="4" place="4" resultid="2877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1719" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3634" />
                    <RANKING order="2" place="2" resultid="7398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1720" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6421" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9173" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9174" daytime="11:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9175" daytime="11:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9176" daytime="11:35" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1595" daytime="09:00" gender="F" number="32" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1597" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5629" />
                    <RANKING order="2" place="2" resultid="2786" />
                    <RANKING order="3" place="3" resultid="7022" />
                    <RANKING order="4" place="4" resultid="7035" />
                    <RANKING order="5" place="5" resultid="2841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1941" />
                    <RANKING order="2" place="2" resultid="6247" />
                    <RANKING order="3" place="3" resultid="5912" />
                    <RANKING order="4" place="4" resultid="2513" />
                    <RANKING order="5" place="5" resultid="5782" />
                    <RANKING order="6" place="6" resultid="5788" />
                    <RANKING order="7" place="-1" resultid="3348" />
                    <RANKING order="8" place="-1" resultid="3812" />
                    <RANKING order="9" place="-1" resultid="7008" />
                    <RANKING order="10" place="-1" resultid="7014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3987" />
                    <RANKING order="2" place="2" resultid="6192" />
                    <RANKING order="3" place="3" resultid="3444" />
                    <RANKING order="4" place="4" resultid="2521" />
                    <RANKING order="5" place="5" resultid="6206" />
                    <RANKING order="6" place="6" resultid="4024" />
                    <RANKING order="7" place="-1" resultid="4973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6255" />
                    <RANKING order="2" place="2" resultid="4259" />
                    <RANKING order="3" place="3" resultid="4267" />
                    <RANKING order="4" place="4" resultid="2738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3544" />
                    <RANKING order="2" place="2" resultid="2448" />
                    <RANKING order="3" place="3" resultid="2618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7351" />
                    <RANKING order="2" place="2" resultid="2647" />
                    <RANKING order="3" place="-1" resultid="5805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3531" />
                    <RANKING order="2" place="2" resultid="3406" />
                    <RANKING order="3" place="3" resultid="6147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7277" />
                    <RANKING order="2" place="2" resultid="3190" />
                    <RANKING order="3" place="3" resultid="4642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3006" />
                    <RANKING order="2" place="2" resultid="3622" />
                    <RANKING order="3" place="3" resultid="3034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1606" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1607" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1608" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1609" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1610" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1611" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1612" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9123" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9124" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9125" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9126" daytime="09:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9127" daytime="09:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1630" daytime="09:40" gender="F" number="34" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1631" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5765" />
                    <RANKING order="2" place="2" resultid="2759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1632" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3577" />
                    <RANKING order="2" place="2" resultid="7222" />
                    <RANKING order="3" place="3" resultid="3419" />
                    <RANKING order="4" place="4" resultid="4847" />
                    <RANKING order="5" place="5" resultid="3962" />
                    <RANKING order="6" place="6" resultid="2083" />
                    <RANKING order="7" place="-1" resultid="2236" />
                    <RANKING order="8" place="-1" resultid="3349" />
                    <RANKING order="9" place="-1" resultid="7162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2766" />
                    <RANKING order="2" place="-1" resultid="2742" />
                    <RANKING order="3" place="-1" resultid="3753" />
                    <RANKING order="4" place="-1" resultid="4701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2536" />
                    <RANKING order="2" place="2" resultid="4250" />
                    <RANKING order="3" place="3" resultid="6256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3552" />
                    <RANKING order="2" place="2" resultid="4906" />
                    <RANKING order="3" place="3" resultid="4212" />
                    <RANKING order="4" place="4" resultid="7259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2457" />
                    <RANKING order="2" place="2" resultid="2864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1638" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3469" />
                    <RANKING order="2" place="2" resultid="2989" />
                    <RANKING order="3" place="3" resultid="2246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1639" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2354" />
                    <RANKING order="2" place="2" resultid="3035" />
                    <RANKING order="3" place="3" resultid="1823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1640" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5571" />
                    <RANKING order="2" place="2" resultid="6405" />
                    <RANKING order="3" place="3" resultid="2004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1641" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1642" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5893" />
                    <RANKING order="2" place="2" resultid="1836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1643" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1644" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1645" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1646" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9138" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9139" daytime="09:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9140" daytime="09:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9141" daytime="09:55" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1664" daytime="10:45" gender="F" number="36" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1665" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2787" />
                    <RANKING order="2" place="2" resultid="3607" />
                    <RANKING order="3" place="3" resultid="1816" />
                    <RANKING order="4" place="4" resultid="4180" />
                    <RANKING order="5" place="5" resultid="2842" />
                    <RANKING order="6" place="6" resultid="7036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1666" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4875" />
                    <RANKING order="2" place="2" resultid="7131" />
                    <RANKING order="3" place="3" resultid="3434" />
                    <RANKING order="4" place="4" resultid="7163" />
                    <RANKING order="5" place="5" resultid="7223" />
                    <RANKING order="6" place="6" resultid="3813" />
                    <RANKING order="7" place="7" resultid="6032" />
                    <RANKING order="8" place="-1" resultid="7170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1667" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3438" />
                    <RANKING order="2" place="2" resultid="2522" />
                    <RANKING order="3" place="3" resultid="3868" />
                    <RANKING order="4" place="4" resultid="3445" />
                    <RANKING order="5" place="5" resultid="3684" />
                    <RANKING order="6" place="6" resultid="3754" />
                    <RANKING order="7" place="7" resultid="4019" />
                    <RANKING order="8" place="8" resultid="4795" />
                    <RANKING order="9" place="-1" resultid="2743" />
                    <RANKING order="10" place="-1" resultid="4702" />
                    <RANKING order="11" place="-1" resultid="4967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1668" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2537" />
                    <RANKING order="2" place="2" resultid="6200" />
                    <RANKING order="3" place="3" resultid="4260" />
                    <RANKING order="4" place="4" resultid="5565" />
                    <RANKING order="5" place="5" resultid="4855" />
                    <RANKING order="6" place="6" resultid="2773" />
                    <RANKING order="7" place="7" resultid="3207" />
                    <RANKING order="8" place="8" resultid="4901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3927" />
                    <RANKING order="2" place="2" resultid="3545" />
                    <RANKING order="3" place="3" resultid="2778" />
                    <RANKING order="4" place="4" resultid="2449" />
                    <RANKING order="5" place="4" resultid="6015" />
                    <RANKING order="6" place="6" resultid="6020" />
                    <RANKING order="7" place="7" resultid="4801" />
                    <RANKING order="8" place="8" resultid="3459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1670" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7235" />
                    <RANKING order="2" place="2" resultid="5806" />
                    <RANKING order="3" place="3" resultid="2648" />
                    <RANKING order="4" place="4" resultid="5616" />
                    <RANKING order="5" place="5" resultid="4208" />
                    <RANKING order="6" place="6" resultid="5578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1671" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3524" />
                    <RANKING order="2" place="2" resultid="3973" />
                    <RANKING order="3" place="3" resultid="3407" />
                    <RANKING order="4" place="4" resultid="6873" />
                    <RANKING order="5" place="5" resultid="2348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1672" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7363" />
                    <RANKING order="2" place="2" resultid="6842" />
                    <RANKING order="3" place="3" resultid="5797" />
                    <RANKING order="4" place="4" resultid="2393" />
                    <RANKING order="5" place="5" resultid="3191" />
                    <RANKING order="6" place="6" resultid="3199" />
                    <RANKING order="7" place="7" resultid="6877" />
                    <RANKING order="8" place="8" resultid="2343" />
                    <RANKING order="9" place="9" resultid="2336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1673" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3164" />
                    <RANKING order="2" place="2" resultid="3007" />
                    <RANKING order="3" place="3" resultid="6411" />
                    <RANKING order="4" place="4" resultid="2355" />
                    <RANKING order="5" place="5" resultid="3338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1674" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6364" />
                    <RANKING order="2" place="2" resultid="5612" />
                    <RANKING order="3" place="3" resultid="4635" />
                    <RANKING order="4" place="4" resultid="5666" />
                    <RANKING order="5" place="5" resultid="7296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1675" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1676" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1677" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1678" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1679" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1680" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9151" daytime="10:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9152" daytime="10:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9153" daytime="10:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9154" daytime="10:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9155" daytime="10:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9156" daytime="10:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9157" daytime="10:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9158" daytime="10:55" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="DOL" nation="POL" region="DOL" clubid="4944" name="10 Brygada Kawalerii Pancernej Swietoszow" shortname="10 Brygada Kawalerii Pancernej">
          <CONTACT city="Świdnica" email="horbacz.marcin@wp.pl" name="Horbacz" phone="603672717" state="LUB" street="Buchałów 12c" zip="66-008" />
          <ATHLETES>
            <ATHLETE birthdate="1984-09-29" firstname="Radosław" gender="M" lastname="Stępień" nation="POL" athleteid="4950">
              <RESULTS>
                <RESULT eventid="1079" points="351" reactiontime="+90" swimtime="00:00:28.70" resultid="4951" heatid="8908" lane="1" entrytime="00:00:28.10" entrycourse="SCM" />
                <RESULT eventid="1273" points="302" reactiontime="+82" swimtime="00:01:06.92" resultid="4952" heatid="8992" lane="1" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="263" reactiontime="+77" swimtime="00:00:39.37" resultid="4953" heatid="9166" lane="3" entrytime="00:00:38.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-27" firstname="Natalia" gender="F" lastname="Szczęsnowicz" nation="POL" athleteid="4961">
              <RESULTS>
                <RESULT eventid="1062" points="433" reactiontime="+79" swimtime="00:00:30.71" resultid="4962" heatid="8892" lane="6" entrytime="00:00:29.65" entrycourse="SCM" />
                <RESULT eventid="1222" points="316" reactiontime="+87" swimtime="00:03:17.52" resultid="4963" heatid="8968" lane="6" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                    <SPLIT distance="100" swimtime="00:01:35.36" />
                    <SPLIT distance="150" swimtime="00:02:26.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="365" reactiontime="+89" swimtime="00:01:11.33" resultid="4964" heatid="8982" lane="7" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="319" reactiontime="+90" swimtime="00:01:31.25" resultid="4965" heatid="9037" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="322" reactiontime="+75" swimtime="00:00:35.55" resultid="4966" heatid="9058" lane="9" entrytime="00:00:34.30" entrycourse="SCM" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="4967" heatid="9157" lane="9" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-16" firstname="Marcin" gender="M" lastname="Horbacz" nation="POL" athleteid="4954">
              <RESULTS>
                <RESULT eventid="1113" points="492" reactiontime="+84" swimtime="00:02:18.84" resultid="4955" heatid="8930" lane="6" entrytime="00:02:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:06.70" />
                    <SPLIT distance="150" swimtime="00:01:45.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="446" reactiontime="+88" swimtime="00:02:37.62" resultid="4956" heatid="8978" lane="9" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                    <SPLIT distance="150" swimtime="00:01:55.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="472" reactiontime="+87" swimtime="00:01:11.38" resultid="4957" heatid="9044" lane="8" entrytime="00:02:30.00" entrycourse="SCM" />
                <RESULT eventid="1508" points="503" reactiontime="+87" swimtime="00:02:04.94" resultid="4958" heatid="9105" lane="2" entrytime="00:02:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="100" swimtime="00:01:01.53" />
                    <SPLIT distance="150" swimtime="00:01:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="487" reactiontime="+85" swimtime="00:00:32.08" resultid="4959" heatid="9159" lane="4" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="4960" heatid="9191" lane="3" entrytime="00:04:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-12-15" firstname="Oskar" gender="M" lastname="Bogucki" nation="POL" athleteid="4945">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="4946" heatid="8903" lane="0" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="4947" heatid="8975" lane="6" entrytime="00:03:10.00" entrycourse="SCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="4948" heatid="9049" lane="2" entrytime="00:01:25.00" entrycourse="SCM" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="4949" heatid="9168" lane="0" entrytime="00:00:37.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4776" name="Akademia Ruchu Andrzej Gadaś">
          <CONTACT name="Budek" phone="505831398" street="Sosnowskiego 6/24" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-12" firstname="Seweryna" gender="F" lastname="Afanasjew" nation="POL" athleteid="4796">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="4797" heatid="8886" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1256" points="124" reactiontime="+108" swimtime="00:01:42.08" resultid="4798" heatid="8979" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="93" reactiontime="+88" swimtime="00:02:05.13" resultid="4799" heatid="9001" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="68" reactiontime="+105" swimtime="00:00:59.63" resultid="4800" heatid="9054" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1664" points="125" reactiontime="+93" swimtime="00:00:57.45" resultid="4801" heatid="9152" lane="1" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-22" firstname="Andrzej" gender="M" lastname="Gadaś" nation="POL" athleteid="4777">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="4778" heatid="8908" lane="7" entrytime="00:00:28.06" />
                <RESULT eventid="1273" points="319" reactiontime="+81" swimtime="00:01:05.72" resultid="4779" heatid="8993" lane="8" entrytime="00:01:06.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="299" reactiontime="+80" swimtime="00:01:15.71" resultid="4780" heatid="9013" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="280" reactiontime="+89" swimtime="00:00:33.30" resultid="4781" heatid="9064" lane="0" entrytime="00:00:35.61" />
                <RESULT eventid="1681" points="337" reactiontime="+83" swimtime="00:00:36.27" resultid="4782" heatid="9168" lane="8" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-20" firstname="Robert" gender="M" lastname="Budek" nation="POL" athleteid="4783">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="4784" heatid="8904" lane="9" entrytime="00:00:30.50" />
                <RESULT eventid="1273" points="216" reactiontime="+107" swimtime="00:01:14.84" resultid="4785" heatid="8991" lane="8" entrytime="00:01:10.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="174" reactiontime="+104" swimtime="00:01:30.67" resultid="4786" heatid="9011" lane="4" entrytime="00:01:27.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="151" reactiontime="+107" swimtime="00:00:40.93" resultid="4787" heatid="9062" lane="4" entrytime="00:00:39.00" />
                <RESULT comment="K14 - Praca nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie) (Time: 11:11)" eventid="1681" reactiontime="+85" status="DSQ" swimtime="00:00:43.99" resultid="4788" heatid="9163" lane="0" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-13" firstname="Iza" gender="F" lastname="Chmielewska" nation="POL" athleteid="4789">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="4790" heatid="8888" lane="9" entrytime="00:00:39.80" />
                <RESULT eventid="1256" points="162" reactiontime="+90" swimtime="00:01:33.55" resultid="4791" heatid="8980" lane="8" entrytime="00:01:31.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="127" reactiontime="+108" swimtime="00:00:48.49" resultid="4792" heatid="9055" lane="2" entrytime="00:00:47.78" />
                <RESULT eventid="1491" points="138" reactiontime="+94" swimtime="00:03:34.04" resultid="4793" heatid="9090" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:40.71" />
                    <SPLIT distance="150" swimtime="00:02:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" status="DNS" swimtime="00:00:00.00" resultid="4794" heatid="9113" lane="4" entrytime="00:08:00.00" />
                <RESULT eventid="1664" points="83" reactiontime="+94" swimtime="00:01:05.83" resultid="4795" heatid="9152" lane="7" entrytime="00:01:08.16" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT comment="G4 - Wykonanie więcej niż jednego pociągnięcia ramioniem (lub obydwoma ramionami jednocześnie) (Time: 11:38)" eventid="1698" reactiontime="+74" status="DSQ" swimtime="00:02:51.37" resultid="4802" heatid="9174" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:01:39.10" />
                    <SPLIT distance="150" swimtime="00:02:10.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4783" number="1" reactiontime="+74" status="DSQ" />
                    <RELAYPOSITION athleteid="4796" number="2" reactiontime="+21" status="DSQ" />
                    <RELAYPOSITION athleteid="4777" number="3" reactiontime="+9" status="DSQ" />
                    <RELAYPOSITION athleteid="4789" number="4" reactiontime="+43" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="4803" heatid="8933" lane="9" entrytime="00:02:50.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4783" number="1" />
                    <RELAYPOSITION athleteid="4777" number="2" />
                    <RELAYPOSITION athleteid="4796" number="3" />
                    <RELAYPOSITION athleteid="4789" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5380" name="Aquasfera Masters Olsztyn">
          <CONTACT email="annamariaaneczka@gmail.com" name="Goździejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1984-06-13" firstname="Michał" gender="M" lastname="Kieres" nation="POL" athleteid="6208">
              <RESULTS>
                <RESULT eventid="1239" points="316" reactiontime="+81" swimtime="00:02:56.75" resultid="6209" heatid="8978" lane="7" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:08.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="316" reactiontime="+81" swimtime="00:01:14.32" resultid="6210" heatid="9017" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="342" reactiontime="+77" swimtime="00:01:19.45" resultid="6211" heatid="9053" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="292" reactiontime="+76" swimtime="00:00:32.85" resultid="6212" heatid="9069" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1613" points="272" reactiontime="+83" swimtime="00:01:14.70" resultid="6213" heatid="9135" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="323" reactiontime="+91" swimtime="00:00:36.78" resultid="6214" heatid="9170" lane="9" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="6265">
              <RESULTS>
                <RESULT eventid="1079" points="369" reactiontime="+82" swimtime="00:00:28.23" resultid="6266" heatid="8908" lane="8" entrytime="00:00:28.20" />
                <RESULT comment="Rekord Polski" eventid="1165" points="379" reactiontime="+85" swimtime="00:19:33.74" resultid="6267" heatid="8940" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                    <SPLIT distance="150" swimtime="00:01:51.45" />
                    <SPLIT distance="200" swimtime="00:02:29.68" />
                    <SPLIT distance="250" swimtime="00:03:08.00" />
                    <SPLIT distance="300" swimtime="00:03:46.84" />
                    <SPLIT distance="350" swimtime="00:04:25.53" />
                    <SPLIT distance="400" swimtime="00:05:04.64" />
                    <SPLIT distance="450" swimtime="00:05:43.69" />
                    <SPLIT distance="500" swimtime="00:06:22.84" />
                    <SPLIT distance="550" swimtime="00:07:02.23" />
                    <SPLIT distance="600" swimtime="00:07:41.34" />
                    <SPLIT distance="650" swimtime="00:08:20.61" />
                    <SPLIT distance="700" swimtime="00:08:59.83" />
                    <SPLIT distance="750" swimtime="00:09:38.78" />
                    <SPLIT distance="800" swimtime="00:10:18.11" />
                    <SPLIT distance="850" swimtime="00:10:57.62" />
                    <SPLIT distance="900" swimtime="00:11:37.39" />
                    <SPLIT distance="950" swimtime="00:12:17.03" />
                    <SPLIT distance="1000" swimtime="00:12:57.05" />
                    <SPLIT distance="1050" swimtime="00:13:36.99" />
                    <SPLIT distance="1100" swimtime="00:14:16.53" />
                    <SPLIT distance="1150" swimtime="00:14:56.17" />
                    <SPLIT distance="1200" swimtime="00:15:36.30" />
                    <SPLIT distance="1250" swimtime="00:16:16.14" />
                    <SPLIT distance="1300" swimtime="00:16:56.48" />
                    <SPLIT distance="1350" swimtime="00:17:36.64" />
                    <SPLIT distance="1400" swimtime="00:18:17.13" />
                    <SPLIT distance="1450" swimtime="00:18:56.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="299" reactiontime="+83" swimtime="00:02:42.28" resultid="6268" heatid="9030" lane="8" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:14.43" />
                    <SPLIT distance="150" swimtime="00:01:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="365" reactiontime="+83" swimtime="00:00:30.49" resultid="6269" heatid="9067" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1613" points="342" reactiontime="+81" swimtime="00:01:09.20" resultid="6270" heatid="9135" lane="9" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="357" reactiontime="+94" swimtime="00:04:59.07" resultid="6271" heatid="9190" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                    <SPLIT distance="150" swimtime="00:01:50.77" />
                    <SPLIT distance="200" swimtime="00:02:28.52" />
                    <SPLIT distance="250" swimtime="00:03:06.60" />
                    <SPLIT distance="300" swimtime="00:03:44.76" />
                    <SPLIT distance="350" swimtime="00:04:22.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-30" firstname="Karol" gender="M" lastname="Dziemian" nation="POL" athleteid="6228">
              <RESULTS>
                <RESULT eventid="1079" points="197" reactiontime="+97" swimtime="00:00:34.80" resultid="6229" heatid="8899" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1273" points="174" reactiontime="+97" swimtime="00:01:20.39" resultid="6230" heatid="8989" lane="9" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="141" reactiontime="+100" swimtime="00:00:41.79" resultid="6231" heatid="9061" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1508" points="169" reactiontime="+105" swimtime="00:02:59.66" resultid="6232" heatid="9097" lane="2" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                    <SPLIT distance="100" swimtime="00:01:25.17" />
                    <SPLIT distance="150" swimtime="00:02:12.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="185" reactiontime="+92" swimtime="00:00:44.25" resultid="6233" heatid="9162" lane="4" entrytime="00:00:44.00" />
                <RESULT eventid="1744" points="146" reactiontime="+117" swimtime="00:06:42.49" resultid="6234" heatid="9182" lane="5" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                    <SPLIT distance="100" swimtime="00:01:35.74" />
                    <SPLIT distance="150" swimtime="00:02:27.37" />
                    <SPLIT distance="200" swimtime="00:03:18.66" />
                    <SPLIT distance="250" swimtime="00:04:09.70" />
                    <SPLIT distance="300" swimtime="00:05:01.20" />
                    <SPLIT distance="350" swimtime="00:05:53.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="6280">
              <RESULTS>
                <RESULT eventid="1096" points="260" reactiontime="+88" swimtime="00:03:10.90" resultid="6281" heatid="8918" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:01:33.51" />
                    <SPLIT distance="150" swimtime="00:02:28.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="319" reactiontime="+92" swimtime="00:11:41.31" resultid="6282" heatid="8939" lane="0" entrytime="00:11:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:01:23.68" />
                    <SPLIT distance="150" swimtime="00:02:07.90" />
                    <SPLIT distance="200" swimtime="00:02:52.20" />
                    <SPLIT distance="250" swimtime="00:03:36.75" />
                    <SPLIT distance="300" swimtime="00:04:20.92" />
                    <SPLIT distance="350" swimtime="00:05:04.85" />
                    <SPLIT distance="400" swimtime="00:05:48.72" />
                    <SPLIT distance="450" swimtime="00:06:32.11" />
                    <SPLIT distance="500" swimtime="00:07:15.80" />
                    <SPLIT distance="550" swimtime="00:08:00.20" />
                    <SPLIT distance="600" swimtime="00:08:43.98" />
                    <SPLIT distance="650" swimtime="00:09:28.41" />
                    <SPLIT distance="700" swimtime="00:10:13.36" />
                    <SPLIT distance="750" swimtime="00:10:57.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="261" reactiontime="+98" swimtime="00:03:30.38" resultid="6283" heatid="8966" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                    <SPLIT distance="100" swimtime="00:01:42.24" />
                    <SPLIT distance="150" swimtime="00:02:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="335" reactiontime="+93" swimtime="00:01:13.41" resultid="6284" heatid="8982" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="322" reactiontime="+94" swimtime="00:02:41.54" resultid="6285" heatid="9089" lane="1" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:01:59.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="241" reactiontime="+96" swimtime="00:06:57.00" resultid="6286" heatid="9114" lane="7" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                    <SPLIT distance="100" swimtime="00:01:44.29" />
                    <SPLIT distance="150" swimtime="00:02:38.27" />
                    <SPLIT distance="200" swimtime="00:03:33.36" />
                    <SPLIT distance="250" swimtime="00:04:28.86" />
                    <SPLIT distance="300" swimtime="00:05:25.71" />
                    <SPLIT distance="350" swimtime="00:06:12.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="318" reactiontime="+83" swimtime="00:05:43.23" resultid="6287" heatid="9180" lane="4" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="100" swimtime="00:01:23.31" />
                    <SPLIT distance="150" swimtime="00:02:07.35" />
                    <SPLIT distance="200" swimtime="00:02:51.53" />
                    <SPLIT distance="250" swimtime="00:03:35.41" />
                    <SPLIT distance="300" swimtime="00:04:19.53" />
                    <SPLIT distance="350" swimtime="00:05:01.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="6248">
              <RESULTS>
                <RESULT eventid="1062" points="391" reactiontime="+88" swimtime="00:00:31.78" resultid="6249" heatid="8890" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1096" points="336" reactiontime="+87" swimtime="00:02:55.26" resultid="6250" heatid="8919" lane="3" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                    <SPLIT distance="100" swimtime="00:01:22.99" />
                    <SPLIT distance="150" swimtime="00:02:17.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="314" reactiontime="+76" swimtime="00:00:37.75" resultid="6251" heatid="8951" lane="5" entrytime="00:00:37.80" />
                <RESULT eventid="1290" points="359" reactiontime="+85" swimtime="00:01:19.71" resultid="6252" heatid="9005" lane="3" entrytime="00:01:21.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="356" reactiontime="+81" swimtime="00:00:34.37" resultid="6253" heatid="9057" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1457" points="293" reactiontime="+74" swimtime="00:01:22.81" resultid="6254" heatid="9076" lane="4" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="308" reactiontime="+86" swimtime="00:01:20.80" resultid="6255" heatid="9126" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="270" reactiontime="+78" swimtime="00:03:04.40" resultid="6256" heatid="9140" lane="6" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                    <SPLIT distance="100" swimtime="00:01:30.69" />
                    <SPLIT distance="150" swimtime="00:02:18.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-04-01" firstname="Piotr" gender="M" lastname="Konopacki" nation="POL" athleteid="6272">
              <RESULTS>
                <RESULT eventid="1079" points="394" reactiontime="+71" swimtime="00:00:27.62" resultid="6273" heatid="8910" lane="9" entrytime="00:00:27.66" />
                <RESULT eventid="1165" points="307" reactiontime="+86" swimtime="00:21:00.13" resultid="6274" heatid="8940" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:13.41" />
                    <SPLIT distance="150" swimtime="00:01:55.99" />
                    <SPLIT distance="200" swimtime="00:02:38.99" />
                    <SPLIT distance="250" swimtime="00:03:22.18" />
                    <SPLIT distance="300" swimtime="00:04:05.57" />
                    <SPLIT distance="350" swimtime="00:04:48.29" />
                    <SPLIT distance="400" swimtime="00:05:31.68" />
                    <SPLIT distance="450" swimtime="00:06:14.74" />
                    <SPLIT distance="500" swimtime="00:06:57.45" />
                    <SPLIT distance="550" swimtime="00:07:40.41" />
                    <SPLIT distance="600" swimtime="00:08:23.42" />
                    <SPLIT distance="650" swimtime="00:09:05.77" />
                    <SPLIT distance="700" swimtime="00:09:48.65" />
                    <SPLIT distance="750" swimtime="00:10:31.41" />
                    <SPLIT distance="800" swimtime="00:11:14.34" />
                    <SPLIT distance="850" swimtime="00:11:57.05" />
                    <SPLIT distance="900" swimtime="00:12:40.08" />
                    <SPLIT distance="950" swimtime="00:13:22.56" />
                    <SPLIT distance="1000" swimtime="00:14:05.34" />
                    <SPLIT distance="1050" swimtime="00:14:47.64" />
                    <SPLIT distance="1100" swimtime="00:15:29.85" />
                    <SPLIT distance="1150" swimtime="00:16:12.09" />
                    <SPLIT distance="1200" swimtime="00:16:53.81" />
                    <SPLIT distance="1250" swimtime="00:17:35.89" />
                    <SPLIT distance="1300" swimtime="00:18:18.03" />
                    <SPLIT distance="1350" swimtime="00:18:59.79" />
                    <SPLIT distance="1400" swimtime="00:19:42.04" />
                    <SPLIT distance="1450" swimtime="00:20:23.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="299" reactiontime="+77" swimtime="00:00:33.20" resultid="6275" heatid="8961" lane="6" entrytime="00:00:32.94" />
                <RESULT eventid="1273" points="347" reactiontime="+81" swimtime="00:01:03.93" resultid="6276" heatid="8995" lane="0" entrytime="00:01:02.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="279" swimtime="00:01:14.84" resultid="6277" heatid="9084" lane="9" entrytime="00:01:14.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="289" reactiontime="+81" swimtime="00:02:30.24" resultid="6278" heatid="9094" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:12.14" />
                    <SPLIT distance="150" swimtime="00:01:53.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="238" reactiontime="+77" swimtime="00:02:51.08" resultid="6279" heatid="9143" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="100" swimtime="00:01:23.22" />
                    <SPLIT distance="150" swimtime="00:02:08.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-13" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="6257">
              <RESULTS>
                <RESULT eventid="1079" points="444" reactiontime="+80" swimtime="00:00:26.54" resultid="6258" heatid="8905" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1113" points="378" reactiontime="+76" swimtime="00:02:31.59" resultid="6259" heatid="8929" lane="7" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="100" swimtime="00:01:12.35" />
                    <SPLIT distance="150" swimtime="00:01:54.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="450" reactiontime="+78" swimtime="00:02:37.16" resultid="6260" heatid="8978" lane="2" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:01:55.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="398" reactiontime="+79" swimtime="00:01:08.87" resultid="6261" heatid="9020" lane="9" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="469" reactiontime="+78" swimtime="00:01:11.57" resultid="6262" heatid="9052" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="302" reactiontime="+81" swimtime="00:01:12.94" resultid="6263" heatid="9084" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 11:18)" eventid="1681" reactiontime="+46" status="DSQ" swimtime="00:00:33.00" resultid="6264" heatid="9170" lane="2" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-01" firstname="Małgorzata" gender="F" lastname="Polito" nation="POL" athleteid="6215">
              <RESULTS>
                <RESULT eventid="1147" points="343" reactiontime="+87" swimtime="00:11:24.48" resultid="6216" heatid="8939" lane="8" entrytime="00:11:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:01:19.22" />
                    <SPLIT distance="150" swimtime="00:02:01.76" />
                    <SPLIT distance="200" swimtime="00:02:45.19" />
                    <SPLIT distance="250" swimtime="00:03:29.14" />
                    <SPLIT distance="300" swimtime="00:04:13.44" />
                    <SPLIT distance="350" swimtime="00:04:57.41" />
                    <SPLIT distance="400" swimtime="00:05:40.99" />
                    <SPLIT distance="450" swimtime="00:06:24.16" />
                    <SPLIT distance="500" swimtime="00:07:07.11" />
                    <SPLIT distance="550" swimtime="00:07:50.32" />
                    <SPLIT distance="600" swimtime="00:08:34.15" />
                    <SPLIT distance="650" swimtime="00:09:18.09" />
                    <SPLIT distance="700" swimtime="00:10:02.22" />
                    <SPLIT distance="750" swimtime="00:10:45.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="357" reactiontime="+84" swimtime="00:02:36.06" resultid="6217" heatid="9092" lane="6" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:01:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="344" reactiontime="+80" swimtime="00:05:34.50" resultid="6218" heatid="9181" lane="9" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                    <SPLIT distance="150" swimtime="00:02:02.01" />
                    <SPLIT distance="200" swimtime="00:02:45.27" />
                    <SPLIT distance="250" swimtime="00:03:27.13" />
                    <SPLIT distance="300" swimtime="00:04:10.15" />
                    <SPLIT distance="350" swimtime="00:04:53.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-12-05" firstname="Aleksandra" gender="F" lastname="Góralska" nation="POL" athleteid="6293">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="6294" heatid="8888" lane="3" entrytime="00:00:37.50" />
                <RESULT eventid="1721" points="219" reactiontime="+116" swimtime="00:06:28.78" resultid="6295" heatid="9179" lane="6" entrytime="00:06:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                    <SPLIT distance="100" swimtime="00:01:30.62" />
                    <SPLIT distance="150" swimtime="00:02:19.25" />
                    <SPLIT distance="200" swimtime="00:03:09.17" />
                    <SPLIT distance="250" swimtime="00:03:59.70" />
                    <SPLIT distance="300" swimtime="00:04:50.69" />
                    <SPLIT distance="350" swimtime="00:05:40.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-09" firstname="Marek" gender="M" lastname="Koźlikowski" nation="POL" athleteid="6235">
              <RESULTS>
                <RESULT eventid="1113" points="230" reactiontime="+95" swimtime="00:02:58.84" resultid="6236" heatid="8924" lane="4" entrytime="00:03:08.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:28.40" />
                    <SPLIT distance="150" swimtime="00:02:18.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="239" reactiontime="+107" swimtime="00:03:13.93" resultid="6237" heatid="8974" lane="8" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.52" />
                    <SPLIT distance="100" swimtime="00:01:35.18" />
                    <SPLIT distance="150" swimtime="00:02:25.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="265" reactiontime="+100" swimtime="00:02:34.55" resultid="6238" heatid="9097" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                    <SPLIT distance="150" swimtime="00:01:55.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="214" reactiontime="+101" swimtime="00:06:33.58" resultid="6239" heatid="9118" lane="5" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:39.70" />
                    <SPLIT distance="150" swimtime="00:02:34.19" />
                    <SPLIT distance="200" swimtime="00:03:27.16" />
                    <SPLIT distance="250" swimtime="00:04:19.17" />
                    <SPLIT distance="300" swimtime="00:05:11.23" />
                    <SPLIT distance="350" swimtime="00:05:53.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="240" reactiontime="+101" swimtime="00:05:41.54" resultid="6240" heatid="9186" lane="0" entrytime="00:06:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:18.70" />
                    <SPLIT distance="150" swimtime="00:02:02.22" />
                    <SPLIT distance="200" swimtime="00:02:46.94" />
                    <SPLIT distance="250" swimtime="00:03:31.97" />
                    <SPLIT distance="300" swimtime="00:04:16.67" />
                    <SPLIT distance="350" swimtime="00:05:00.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="6219">
              <RESULTS>
                <RESULT eventid="1079" points="467" reactiontime="+73" swimtime="00:00:26.11" resultid="6220" heatid="8911" lane="8" entrytime="00:00:26.80" />
                <RESULT eventid="1113" points="419" reactiontime="+82" swimtime="00:02:26.46" resultid="6221" heatid="8930" lane="7" entrytime="00:02:25.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="100" swimtime="00:01:11.19" />
                    <SPLIT distance="150" swimtime="00:01:53.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="504" reactiontime="+76" swimtime="00:00:56.45" resultid="6222" heatid="8998" lane="5" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="367" reactiontime="+88" swimtime="00:02:31.53" resultid="6223" heatid="9029" lane="7" entrytime="00:02:45.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:12.95" />
                    <SPLIT distance="150" swimtime="00:01:52.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="492" reactiontime="+82" swimtime="00:02:05.81" resultid="6224" heatid="9105" lane="6" entrytime="00:02:06.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="100" swimtime="00:01:01.32" />
                    <SPLIT distance="150" swimtime="00:01:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="384" reactiontime="+89" swimtime="00:05:23.81" resultid="6225" heatid="9122" lane="1" entrytime="00:05:17.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:10.57" />
                    <SPLIT distance="150" swimtime="00:01:56.29" />
                    <SPLIT distance="200" swimtime="00:02:39.94" />
                    <SPLIT distance="250" swimtime="00:03:26.01" />
                    <SPLIT distance="300" swimtime="00:04:12.55" />
                    <SPLIT distance="350" swimtime="00:04:49.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="461" reactiontime="+79" swimtime="00:01:02.70" resultid="6226" heatid="9136" lane="8" entrytime="00:01:03.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="486" reactiontime="+96" swimtime="00:04:29.80" resultid="6227" heatid="9192" lane="1" entrytime="00:04:31.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                    <SPLIT distance="150" swimtime="00:01:39.99" />
                    <SPLIT distance="200" swimtime="00:02:14.15" />
                    <SPLIT distance="250" swimtime="00:02:48.28" />
                    <SPLIT distance="300" swimtime="00:03:22.39" />
                    <SPLIT distance="350" swimtime="00:03:56.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="Piekut" nation="POL" athleteid="6241">
              <RESULTS>
                <RESULT eventid="1096" points="352" reactiontime="+85" swimtime="00:02:52.47" resultid="6242" heatid="8919" lane="0" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:19.85" />
                    <SPLIT distance="150" swimtime="00:02:10.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="331" reactiontime="+86" swimtime="00:03:14.37" resultid="6243" heatid="8966" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:34.89" />
                    <SPLIT distance="150" swimtime="00:02:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="393" reactiontime="+85" swimtime="00:02:43.28" resultid="6244" heatid="9024" lane="4" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="100" swimtime="00:01:18.73" />
                    <SPLIT distance="150" swimtime="00:02:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="378" reactiontime="+87" swimtime="00:00:33.71" resultid="6245" heatid="9058" lane="0" entrytime="00:00:34.20" />
                <RESULT eventid="1555" points="346" reactiontime="+94" swimtime="00:06:09.90" resultid="6246" heatid="9115" lane="7" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:22.99" />
                    <SPLIT distance="150" swimtime="00:02:12.17" />
                    <SPLIT distance="200" swimtime="00:03:00.40" />
                    <SPLIT distance="250" swimtime="00:03:52.03" />
                    <SPLIT distance="300" swimtime="00:04:43.89" />
                    <SPLIT distance="350" swimtime="00:05:27.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="375" reactiontime="+78" swimtime="00:01:15.67" resultid="6247" heatid="9127" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-18" firstname="Bogdan" gender="M" lastname="Milewski" nation="POL" athleteid="6288">
              <RESULTS>
                <RESULT eventid="1079" points="272" reactiontime="+94" swimtime="00:00:31.25" resultid="6289" heatid="8902" lane="0" entrytime="00:00:31.60" />
                <RESULT eventid="1307" points="246" reactiontime="+98" swimtime="00:01:20.78" resultid="6290" heatid="9012" lane="4" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="233" reactiontime="+89" swimtime="00:00:35.39" resultid="6291" heatid="9063" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1681" points="289" reactiontime="+101" swimtime="00:00:38.17" resultid="6292" heatid="9166" lane="0" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-26" firstname="Aleksandra" gender="F" lastname="Przybysz" nation="POL" athleteid="6201">
              <RESULTS>
                <RESULT eventid="1147" points="317" reactiontime="+75" swimtime="00:11:42.27" resultid="6202" heatid="8938" lane="3" entrytime="00:12:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                    <SPLIT distance="150" swimtime="00:02:06.63" />
                    <SPLIT distance="200" swimtime="00:02:50.84" />
                    <SPLIT distance="250" swimtime="00:03:34.85" />
                    <SPLIT distance="300" swimtime="00:04:19.48" />
                    <SPLIT distance="350" swimtime="00:05:03.72" />
                    <SPLIT distance="400" swimtime="00:05:48.16" />
                    <SPLIT distance="450" swimtime="00:06:31.86" />
                    <SPLIT distance="500" swimtime="00:07:16.00" />
                    <SPLIT distance="550" swimtime="00:08:00.66" />
                    <SPLIT distance="600" swimtime="00:08:45.71" />
                    <SPLIT distance="650" swimtime="00:09:30.39" />
                    <SPLIT distance="700" swimtime="00:10:15.06" />
                    <SPLIT distance="750" swimtime="00:10:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="322" reactiontime="+84" swimtime="00:01:14.38" resultid="6203" heatid="8981" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="240" reactiontime="+83" swimtime="00:03:12.41" resultid="6204" heatid="9024" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:33.36" />
                    <SPLIT distance="150" swimtime="00:02:22.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="323" reactiontime="+85" swimtime="00:02:41.43" resultid="6205" heatid="9091" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                    <SPLIT distance="150" swimtime="00:02:01.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="264" reactiontime="+89" swimtime="00:01:25.05" resultid="6206" heatid="9125" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="317" reactiontime="+90" swimtime="00:05:43.83" resultid="6207" heatid="9180" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:22.58" />
                    <SPLIT distance="150" swimtime="00:02:06.71" />
                    <SPLIT distance="200" swimtime="00:02:50.77" />
                    <SPLIT distance="250" swimtime="00:03:34.65" />
                    <SPLIT distance="300" swimtime="00:04:18.72" />
                    <SPLIT distance="350" swimtime="00:05:02.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="391" reactiontime="+82" swimtime="00:02:03.75" resultid="6301" heatid="9034" lane="4" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:07.86" />
                    <SPLIT distance="150" swimtime="00:01:36.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6265" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="6257" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="6219" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="6272" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="419" reactiontime="+73" swimtime="00:01:50.38" resultid="6302" heatid="9111" lane="5" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.89" />
                    <SPLIT distance="100" swimtime="00:00:56.36" />
                    <SPLIT distance="150" swimtime="00:01:23.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6257" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="6265" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="6272" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="6219" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="233" reactiontime="+75" swimtime="00:02:26.92" resultid="6303" heatid="9033" lane="2" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:21.57" />
                    <SPLIT distance="150" swimtime="00:01:54.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6288" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="6228" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="6208" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="6235" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="262" reactiontime="+80" swimtime="00:02:08.93" resultid="6304" heatid="9110" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:00:50.14" />
                    <SPLIT distance="150" swimtime="00:01:33.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6208" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="6235" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="6288" number="3" />
                    <RELAYPOSITION athleteid="6228" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1525" points="356" reactiontime="+84" swimtime="00:02:12.87" resultid="6299" heatid="9108" lane="6" entrytime="00:02:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:05.41" />
                    <SPLIT distance="150" swimtime="00:01:38.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6248" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="6241" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="6215" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="6201" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1358" points="350" reactiontime="+79" swimtime="00:02:27.56" resultid="6300" heatid="9031" lane="2" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="150" swimtime="00:01:53.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6248" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="6215" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="6241" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="6280" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="339" reactiontime="+80" swimtime="00:01:58.46" resultid="6297" heatid="8935" lane="7" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                    <SPLIT distance="100" swimtime="00:00:54.05" />
                    <SPLIT distance="150" swimtime="00:01:14.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6219" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="6257" number="2" reactiontime="+8" />
                    <RELAYPOSITION athleteid="6241" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="6248" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="330" reactiontime="+80" swimtime="00:02:10.91" resultid="6298" heatid="9176" lane="0" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                    <SPLIT distance="150" swimtime="00:01:44.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6248" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="6257" number="2" reactiontime="+13" />
                    <RELAYPOSITION athleteid="6241" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="6219" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1698" points="272" reactiontime="+67" swimtime="00:02:19.62" resultid="6305" heatid="9175" lane="3" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:15.01" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6272" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="6215" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="6265" number="3" reactiontime="+13" />
                    <RELAYPOSITION athleteid="6280" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1130" points="279" reactiontime="+76" swimtime="00:02:06.32" resultid="6306" heatid="8934" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="100" swimtime="00:00:57.88" />
                    <SPLIT distance="150" swimtime="00:01:32.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6272" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="6265" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="6280" number="3" reactiontime="+187" />
                    <RELAYPOSITION athleteid="6201" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1130" points="253" reactiontime="+96" swimtime="00:02:10.57" resultid="6296" heatid="8934" lane="9" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:05.48" />
                    <SPLIT distance="150" swimtime="00:01:39.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6235" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="6215" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="6228" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="6293" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1698" points="208" reactiontime="+70" swimtime="00:02:32.56" resultid="6307" heatid="9175" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:01:54.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6288" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="6208" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="6201" number="3" reactiontime="+5" />
                    <RELAYPOSITION athleteid="6293" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AQUNI" nation="SVK" region="ZSO" clubid="2215" name="AQUATICS Nitra">
          <ATHLETES>
            <ATHLETE birthdate="1970-02-03" firstname="Peter" gender="M" lastname="Čigáš" nation="SVK" license="SVK15844" athleteid="3446">
              <RESULTS>
                <RESULT eventid="1205" points="381" reactiontime="+174" swimtime="00:00:30.64" resultid="3447" heatid="8963" lane="1" entrytime="00:00:30.73" entrycourse="SCM" />
                <RESULT eventid="1474" points="397" reactiontime="+70" swimtime="00:01:06.57" resultid="3448" heatid="9086" lane="2" entrytime="00:01:05.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="411" reactiontime="+94" swimtime="00:02:13.63" resultid="3449" heatid="9103" lane="5" entrytime="00:02:12.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:06.24" />
                    <SPLIT distance="150" swimtime="00:01:39.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="389" reactiontime="+66" swimtime="00:02:25.35" resultid="3450" heatid="9149" lane="7" entrytime="00:02:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:11.22" />
                    <SPLIT distance="150" swimtime="00:01:48.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="376" reactiontime="+95" swimtime="00:04:53.98" resultid="3451" heatid="9191" lane="9" entrytime="00:04:48.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:09.38" />
                    <SPLIT distance="150" swimtime="00:01:46.13" />
                    <SPLIT distance="200" swimtime="00:02:23.32" />
                    <SPLIT distance="250" swimtime="00:03:00.20" />
                    <SPLIT distance="300" swimtime="00:04:16.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-05-08" firstname="Karol" gender="M" lastname="Lacko" nation="SVK" license="SVK16793" athleteid="3452">
              <RESULTS>
                <RESULT eventid="1508" points="399" reactiontime="+83" swimtime="00:02:14.97" resultid="3453" heatid="9103" lane="8" entrytime="00:02:16.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:05.89" />
                    <SPLIT distance="150" swimtime="00:01:40.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="408" reactiontime="+91" swimtime="00:04:45.99" resultid="3454" heatid="9190" lane="7" entrytime="00:04:55.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:08.77" />
                    <SPLIT distance="150" swimtime="00:01:44.88" />
                    <SPLIT distance="200" swimtime="00:02:20.62" />
                    <SPLIT distance="300" swimtime="00:03:32.95" />
                    <SPLIT distance="350" swimtime="00:04:09.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="388" reactiontime="+82" swimtime="00:01:01.60" resultid="3455" heatid="8994" lane="3" entrytime="00:01:03.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2032" name="Astoria Bydgoszcz">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-01" firstname="Wawrzyniec" gender="M" lastname="Mańczak" nation="POL" athleteid="2033">
              <RESULTS>
                <RESULT eventid="1205" points="166" reactiontime="+81" swimtime="00:00:40.43" resultid="2034" heatid="8958" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="1307" points="151" reactiontime="+115" swimtime="00:01:35.12" resultid="2035" heatid="9010" lane="6" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="145" reactiontime="+80" swimtime="00:01:33.11" resultid="2036" heatid="9081" lane="8" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="131" reactiontime="+80" swimtime="00:03:28.67" resultid="2037" heatid="9145" lane="5" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                    <SPLIT distance="100" swimtime="00:01:40.49" />
                    <SPLIT distance="150" swimtime="00:02:36.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="SLA" clubid="5746" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1990-10-09" firstname="Arkadiusz" gender="M" lastname="Kula" nation="POL" license="100611700280" athleteid="5766">
              <RESULTS>
                <RESULT eventid="1273" points="593" reactiontime="+70" swimtime="00:00:53.47" resultid="5768" heatid="9000" lane="7" entrytime="00:00:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="674" reactiontime="+67" swimtime="00:00:57.77" resultid="5769" heatid="9021" lane="3" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="592" reactiontime="+67" swimtime="00:00:25.96" resultid="5770" heatid="9073" lane="2" entrytime="00:00:25.80" />
                <RESULT eventid="1508" points="571" reactiontime="+78" swimtime="00:01:59.71" resultid="5771" heatid="9106" lane="0" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                    <SPLIT distance="100" swimtime="00:00:58.41" />
                    <SPLIT distance="150" swimtime="00:01:29.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1931-04-27" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" athleteid="5752">
              <RESULTS>
                <RESULT eventid="1079" points="36" reactiontime="+102" swimtime="00:01:01.22" resultid="5753" heatid="8895" lane="7" entrytime="00:01:00.21" />
                <RESULT eventid="1165" points="30" reactiontime="+97" swimtime="00:45:14.51" resultid="5754" heatid="8940" lane="5" entrytime="00:44:50.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.39" />
                    <SPLIT distance="100" swimtime="00:02:48.83" />
                    <SPLIT distance="150" swimtime="00:04:22.42" />
                    <SPLIT distance="200" swimtime="00:05:51.42" />
                    <SPLIT distance="250" swimtime="00:07:25.03" />
                    <SPLIT distance="300" swimtime="00:08:50.57" />
                    <SPLIT distance="350" swimtime="00:10:25.05" />
                    <SPLIT distance="400" swimtime="00:11:52.64" />
                    <SPLIT distance="450" swimtime="00:13:28.68" />
                    <SPLIT distance="500" swimtime="00:14:55.91" />
                    <SPLIT distance="550" swimtime="00:16:30.95" />
                    <SPLIT distance="600" swimtime="00:17:57.05" />
                    <SPLIT distance="650" swimtime="00:19:32.74" />
                    <SPLIT distance="700" swimtime="00:21:00.37" />
                    <SPLIT distance="750" swimtime="00:22:36.67" />
                    <SPLIT distance="800" swimtime="00:24:04.20" />
                    <SPLIT distance="850" swimtime="00:25:39.82" />
                    <SPLIT distance="900" swimtime="00:27:08.96" />
                    <SPLIT distance="950" swimtime="00:28:45.22" />
                    <SPLIT distance="1000" swimtime="00:30:12.59" />
                    <SPLIT distance="1050" swimtime="00:31:48.33" />
                    <SPLIT distance="1100" swimtime="00:33:14.50" />
                    <SPLIT distance="1150" swimtime="00:34:50.22" />
                    <SPLIT distance="1200" swimtime="00:36:16.94" />
                    <SPLIT distance="1250" swimtime="00:37:53.46" />
                    <SPLIT distance="1300" swimtime="00:39:20.54" />
                    <SPLIT distance="1350" swimtime="00:40:56.40" />
                    <SPLIT distance="1400" swimtime="00:42:22.73" />
                    <SPLIT distance="1450" swimtime="00:43:56.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="46" reactiontime="+104" swimtime="00:05:35.77" resultid="5755" heatid="8971" lane="4" entrytime="00:05:23.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.53" />
                    <SPLIT distance="100" swimtime="00:02:43.19" />
                    <SPLIT distance="150" swimtime="00:04:12.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="34" reactiontime="+100" swimtime="00:02:17.47" resultid="5756" heatid="8986" lane="7" entrytime="00:02:21.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="43" reactiontime="+90" swimtime="00:02:38.73" resultid="5757" heatid="9044" lane="9" entrytime="00:02:38.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="32" reactiontime="+96" swimtime="00:05:10.56" resultid="5758" heatid="9094" lane="4" entrytime="00:05:03.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.86" />
                    <SPLIT distance="100" swimtime="00:02:31.30" />
                    <SPLIT distance="150" swimtime="00:03:55.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="44" reactiontime="+109" swimtime="00:01:11.01" resultid="5759" heatid="9160" lane="1" entrytime="00:01:05.73" />
                <RESULT eventid="1744" points="33" reactiontime="+95" swimtime="00:10:56.63" resultid="5760" heatid="9182" lane="2" entrytime="00:10:46.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.70" />
                    <SPLIT distance="100" swimtime="00:02:46.21" />
                    <SPLIT distance="150" swimtime="00:04:13.08" />
                    <SPLIT distance="200" swimtime="00:05:35.44" />
                    <SPLIT distance="250" swimtime="00:06:58.17" />
                    <SPLIT distance="300" swimtime="00:08:20.76" />
                    <SPLIT distance="350" swimtime="00:09:42.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-06-20" firstname="Martyna" gender="F" lastname="Szkrobocz" nation="POL" license="100611600220" athleteid="5761">
              <RESULTS>
                <RESULT eventid="1062" points="483" reactiontime="+80" swimtime="00:00:29.62" resultid="5762" heatid="8892" lane="7" entrytime="00:00:29.70" />
                <RESULT eventid="1187" points="461" reactiontime="+73" swimtime="00:00:33.22" resultid="5763" heatid="8953" lane="6" entrytime="00:00:32.50" />
                <RESULT eventid="1457" points="486" reactiontime="+68" swimtime="00:01:09.98" resultid="5764" heatid="9078" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="519" reactiontime="+67" swimtime="00:02:28.36" resultid="5765" heatid="9141" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:51.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZS PWSZ R" nation="POL" region="SLA" clubid="3151" name="Azs Pwsz Raciborz">
          <CONTACT city="Racibórz" email="adip45@poczta.onet.pl" name="PIECHULA" state="ŚLĄSK" street="Słowackiego 55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-11-04" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="3152">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="3153" heatid="8925" lane="8" entrytime="00:03:04.70" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="3154" heatid="8974" lane="4" entrytime="00:03:19.80" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="3155" heatid="9028" lane="6" entrytime="00:03:07.50" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="3156" heatid="9048" lane="1" entrytime="00:01:29.80" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="3157" heatid="9119" lane="3" entrytime="00:06:29.60" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="3158" heatid="9146" lane="2" entrytime="00:03:11.60" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="3159" heatid="9165" lane="6" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LOD" nation="POL" region="LOD" clubid="5621" name="Azs Uł Pł">
          <CONTACT name="AZS UŁ PŁ" state="LOD" street="Styrska" />
          <ATHLETES>
            <ATHLETE birthdate="1994-04-30" firstname="Katarzyna" gender="F" lastname="Stasinowska" nation="POL" license="102305600024" athleteid="5622">
              <RESULTS>
                <RESULT eventid="1062" points="611" reactiontime="+69" swimtime="00:00:27.38" resultid="5623" heatid="8893" lane="5" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1096" points="501" reactiontime="+70" swimtime="00:02:33.37" resultid="5624" heatid="8920" lane="5" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="572" reactiontime="+72" swimtime="00:01:01.42" resultid="5625" heatid="8984" lane="3" entrytime="00:01:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="529" reactiontime="+72" swimtime="00:01:10.07" resultid="5626" heatid="9007" lane="6" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="587" reactiontime="+70" swimtime="00:00:29.11" resultid="5627" heatid="9059" lane="4" entrytime="00:00:28.80" entrycourse="SCM" />
                <RESULT eventid="1491" points="522" reactiontime="+72" swimtime="00:02:17.52" resultid="5628" heatid="9093" lane="5" entrytime="00:02:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:06.64" />
                    <SPLIT distance="150" swimtime="00:01:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="556" reactiontime="+73" swimtime="00:01:06.38" resultid="5629" heatid="9127" lane="4" entrytime="00:01:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4146" name="AZS WSB Dąbrowa Górnicza.">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="4147">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="4148" heatid="8913" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="4149" heatid="8945" lane="2" entrytime="00:21:20.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="4150" heatid="8962" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1239" points="278" reactiontime="+87" swimtime="00:03:04.40" resultid="4151" heatid="8977" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                    <SPLIT distance="100" swimtime="00:01:26.95" />
                    <SPLIT distance="150" swimtime="00:02:15.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="4152" heatid="9051" lane="2" entrytime="00:01:20.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="4153" heatid="9083" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="4154" heatid="9147" lane="6" entrytime="00:02:45.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="4155" heatid="9171" lane="5" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="HUN" clubid="2167" name="Budapesti Delfinek">
          <CONTACT city="Budapest" email="drpetergulyas@gmail.com" fax="+3612025040" name="dr. Gulyás Péter" phone="+36309492809" state="HUN" street="Alkotás u. 31. fszt. 4." zip="1123" />
          <ATHLETES>
            <ATHLETE birthdate="1951-10-09" firstname="Peter" gender="M" lastname="Gulyas" nation="HUN" athleteid="2181">
              <RESULTS>
                <RESULT eventid="1079" points="340" reactiontime="+74" swimtime="00:00:29.00" resultid="2182" heatid="8905" lane="4" entrytime="00:00:29.80" entrycourse="SCM" />
                <RESULT eventid="1113" points="255" reactiontime="+85" swimtime="00:02:52.78" resultid="2183" heatid="8925" lane="4" entrytime="00:02:55.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:23.72" />
                    <SPLIT distance="150" swimtime="00:02:13.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="255" reactiontime="+80" swimtime="00:03:09.90" resultid="2184" heatid="8975" lane="4" entrytime="00:03:06.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:01:29.25" />
                    <SPLIT distance="150" swimtime="00:02:18.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="319" reactiontime="+77" swimtime="00:01:14.14" resultid="2185" heatid="9015" lane="4" entrytime="00:01:14.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="288" reactiontime="+84" swimtime="00:01:24.14" resultid="2186" heatid="9050" lane="3" entrytime="00:01:22.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="272" reactiontime="+82" swimtime="00:00:33.61" resultid="2187" heatid="9066" lane="1" entrytime="00:00:32.74" entrycourse="SCM" />
                <RESULT eventid="1613" points="193" reactiontime="+84" swimtime="00:01:23.79" resultid="2188" heatid="9132" lane="1" entrytime="00:01:22.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="323" reactiontime="+75" swimtime="00:00:36.77" resultid="2189" heatid="9169" lane="3" entrytime="00:00:35.69" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CM UJ MAST" nation="POL" region="MAL" clubid="4040" name="Collegium Medicum UJ Masters Kraków" shortname="Collegium Medicum UJ Masters K">
          <CONTACT city="Kraków" email="jackwi@poczta.onet.pl" name="Kwiatkowski Jacek" phone="601648456" street="Łużycka 49" zip="30658" />
          <ATHLETES>
            <ATHLETE birthdate="1957-03-25" firstname="Jacek" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="4303">
              <RESULTS>
                <RESULT eventid="1079" points="218" reactiontime="+73" swimtime="00:00:33.62" resultid="4304" heatid="8902" lane="9" entrytime="00:00:31.68" entrycourse="SCM" />
                <RESULT eventid="1165" points="212" reactiontime="+115" swimtime="00:23:43.92" resultid="4305" heatid="8943" lane="0" entrytime="00:24:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.93" />
                    <SPLIT distance="150" swimtime="00:02:14.44" />
                    <SPLIT distance="200" swimtime="00:03:02.21" />
                    <SPLIT distance="250" swimtime="00:03:49.98" />
                    <SPLIT distance="300" swimtime="00:04:38.07" />
                    <SPLIT distance="350" swimtime="00:05:26.51" />
                    <SPLIT distance="400" swimtime="00:06:15.14" />
                    <SPLIT distance="450" swimtime="00:07:03.66" />
                    <SPLIT distance="500" swimtime="00:07:51.26" />
                    <SPLIT distance="550" swimtime="00:08:39.20" />
                    <SPLIT distance="600" swimtime="00:09:27.01" />
                    <SPLIT distance="650" swimtime="00:10:15.46" />
                    <SPLIT distance="700" swimtime="00:11:03.17" />
                    <SPLIT distance="750" swimtime="00:11:51.21" />
                    <SPLIT distance="800" swimtime="00:12:39.46" />
                    <SPLIT distance="850" swimtime="00:13:26.92" />
                    <SPLIT distance="900" swimtime="00:14:14.65" />
                    <SPLIT distance="950" swimtime="00:15:02.23" />
                    <SPLIT distance="1000" swimtime="00:15:50.31" />
                    <SPLIT distance="1050" swimtime="00:16:38.11" />
                    <SPLIT distance="1100" swimtime="00:17:26.03" />
                    <SPLIT distance="1150" swimtime="00:18:14.26" />
                    <SPLIT distance="1200" swimtime="00:19:01.72" />
                    <SPLIT distance="1250" swimtime="00:19:49.38" />
                    <SPLIT distance="1300" swimtime="00:20:37.18" />
                    <SPLIT distance="1350" swimtime="00:21:25.10" />
                    <SPLIT distance="1400" swimtime="00:22:13.22" />
                    <SPLIT distance="1450" swimtime="00:23:01.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-08-22" firstname="Mirosław" gender="M" lastname="Woźniak" nation="POL" athleteid="4075">
              <RESULTS>
                <RESULT eventid="1113" points="316" reactiontime="+93" swimtime="00:02:40.89" resultid="4076" heatid="8928" lane="4" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:15.40" />
                    <SPLIT distance="150" swimtime="00:02:02.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="339" reactiontime="+88" swimtime="00:01:12.65" resultid="4077" heatid="9017" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="295" reactiontime="+94" swimtime="00:02:29.13" resultid="4078" heatid="9101" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:09.52" />
                    <SPLIT distance="150" swimtime="00:01:49.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-29" firstname="Mariusz" gender="M" lastname="Baranik" nation="POL" athleteid="4070">
              <RESULTS>
                <RESULT eventid="1079" points="429" reactiontime="+81" swimtime="00:00:26.85" resultid="4071" heatid="8910" lane="8" entrytime="00:00:27.10" />
                <RESULT eventid="1273" points="431" reactiontime="+85" swimtime="00:00:59.47" resultid="4072" heatid="8996" lane="7" entrytime="00:01:01.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="390" reactiontime="+82" swimtime="00:01:09.28" resultid="4073" heatid="9017" lane="6" entrytime="00:01:10.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="423" reactiontime="+80" swimtime="00:00:29.04" resultid="4074" heatid="9070" lane="7" entrytime="00:00:29.10" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02711" nation="POL" region="SLA" clubid="2363" name="CSiR MOS Dąbrowa Górnicza">
          <CONTACT name="Waliczek Mariusz" phone="606448210" />
          <ATHLETES>
            <ATHLETE birthdate="1993-07-28" firstname="Łukasz" gender="M" lastname="Furman" nation="POL" license="102711700235" athleteid="2381">
              <RESULTS>
                <RESULT eventid="1474" points="611" reactiontime="+62" swimtime="00:00:57.66" resultid="2382" heatid="9087" lane="4" entrytime="00:00:56.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="578" reactiontime="+58" swimtime="00:02:07.32" resultid="2383" heatid="9150" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="100" swimtime="00:01:02.34" />
                    <SPLIT distance="150" swimtime="00:01:34.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DMLOD" nation="POL" region="LOD" clubid="2412" name="Delfin Masters Łódź">
          <CONTACT city="Łódź" email="cewa@poczta.fm" name="Cieplucha Ewa" phone="604627966" street="Retkińska 74 m 18" zip="94-004" />
          <ATHLETES>
            <ATHLETE birthdate="1974-04-11" firstname="Rafał" gender="M" lastname="Maciejewski" nation="POL" athleteid="2421">
              <RESULTS>
                <RESULT eventid="1079" points="249" reactiontime="+100" swimtime="00:00:32.19" resultid="2422" heatid="8901" lane="0" entrytime="00:00:32.01" />
                <RESULT eventid="1273" points="238" reactiontime="+92" swimtime="00:01:12.49" resultid="2423" heatid="8990" lane="0" entrytime="00:01:13.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-24" firstname="Piotr" gender="M" lastname="Gaede" nation="POL" athleteid="2418">
              <RESULTS>
                <RESULT eventid="1406" points="287" reactiontime="+86" swimtime="00:01:24.28" resultid="2419" heatid="9049" lane="4" entrytime="00:01:24.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="278" reactiontime="+89" swimtime="00:00:38.68" resultid="2420" heatid="9167" lane="0" entrytime="00:00:38.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-11" firstname="Arkadiusz" gender="M" lastname="Piecyk" nation="POL" athleteid="2424">
              <RESULTS>
                <RESULT eventid="1079" points="352" reactiontime="+94" swimtime="00:00:28.69" resultid="2425" heatid="8901" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1205" points="325" reactiontime="+73" swimtime="00:00:32.31" resultid="2426" heatid="8959" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1474" points="349" swimtime="00:01:09.48" resultid="2427" heatid="9083" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="315" reactiontime="+77" swimtime="00:02:35.84" resultid="2428" heatid="9147" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                    <SPLIT distance="150" swimtime="00:01:55.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-03-06" firstname="Tomasz" gender="M" lastname="Wiaderny" nation="POL" athleteid="2413">
              <RESULTS>
                <RESULT eventid="1079" points="218" reactiontime="+95" swimtime="00:00:33.65" resultid="2414" heatid="8902" lane="8" entrytime="00:00:31.50" />
                <RESULT eventid="1273" points="192" reactiontime="+93" swimtime="00:01:17.89" resultid="2415" heatid="8989" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="171" reactiontime="+104" swimtime="00:00:39.26" resultid="2416" heatid="9063" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1508" points="163" reactiontime="+96" swimtime="00:03:01.75" resultid="2417" heatid="9097" lane="3" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:11.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-02-25" firstname="Jacek" gender="M" lastname="Kadłubiec" nation="POL" athleteid="2429">
              <RESULTS>
                <RESULT eventid="1406" points="293" reactiontime="+112" swimtime="00:01:23.71" resultid="2430" heatid="9046" lane="1" entrytime="00:01:33.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="290" reactiontime="+100" swimtime="00:00:38.14" resultid="2431" heatid="9168" lane="7" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="267" reactiontime="+85" swimtime="00:02:08.14" resultid="2432" heatid="9109" lane="3" entrytime="00:02:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:05.57" />
                    <SPLIT distance="150" swimtime="00:01:36.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2413" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="2418" number="2" reactiontime="+8" />
                    <RELAYPOSITION athleteid="2429" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2421" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="2433" heatid="9032" lane="5" entrytime="00:02:36.99">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2424" number="1" />
                    <RELAYPOSITION athleteid="2429" number="2" />
                    <RELAYPOSITION athleteid="2413" number="3" />
                    <RELAYPOSITION athleteid="2421" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2990" name="Gdynia Masters">
          <CONTACT name="Mysiak" />
          <ATHLETES>
            <ATHLETE birthdate="1953-01-01" firstname="Leszek" gender="M" lastname="Kubicki" nation="POL" athleteid="3008">
              <RESULTS>
                <RESULT eventid="1079" points="250" reactiontime="+99" swimtime="00:00:32.16" resultid="3009" heatid="8899" lane="4" entrytime="00:00:34.15" />
                <RESULT eventid="1165" points="228" reactiontime="+100" swimtime="00:23:10.55" resultid="3010" heatid="8943" lane="8" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:20.24" />
                    <SPLIT distance="150" swimtime="00:02:05.20" />
                    <SPLIT distance="200" swimtime="00:02:51.23" />
                    <SPLIT distance="250" swimtime="00:03:37.26" />
                    <SPLIT distance="300" swimtime="00:04:23.62" />
                    <SPLIT distance="350" swimtime="00:05:09.75" />
                    <SPLIT distance="400" swimtime="00:05:55.68" />
                    <SPLIT distance="450" swimtime="00:06:42.00" />
                    <SPLIT distance="500" swimtime="00:07:28.63" />
                    <SPLIT distance="550" swimtime="00:08:14.81" />
                    <SPLIT distance="600" swimtime="00:09:01.62" />
                    <SPLIT distance="650" swimtime="00:09:48.53" />
                    <SPLIT distance="700" swimtime="00:10:34.97" />
                    <SPLIT distance="750" swimtime="00:11:22.13" />
                    <SPLIT distance="800" swimtime="00:12:09.05" />
                    <SPLIT distance="850" swimtime="00:12:56.23" />
                    <SPLIT distance="900" swimtime="00:13:43.06" />
                    <SPLIT distance="950" swimtime="00:14:29.87" />
                    <SPLIT distance="1000" swimtime="00:15:17.16" />
                    <SPLIT distance="1050" swimtime="00:16:03.90" />
                    <SPLIT distance="1100" swimtime="00:16:51.67" />
                    <SPLIT distance="1150" swimtime="00:17:39.44" />
                    <SPLIT distance="1200" swimtime="00:18:27.06" />
                    <SPLIT distance="1250" swimtime="00:19:14.64" />
                    <SPLIT distance="1300" swimtime="00:20:02.86" />
                    <SPLIT distance="1350" swimtime="00:20:50.17" />
                    <SPLIT distance="1400" swimtime="00:21:38.07" />
                    <SPLIT distance="1450" swimtime="00:22:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="220" reactiontime="+105" swimtime="00:01:14.44" resultid="3011" heatid="8990" lane="9" entrytime="00:01:14.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="194" reactiontime="+102" swimtime="00:01:27.41" resultid="3012" heatid="9011" lane="6" entrytime="00:01:28.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="214" reactiontime="+103" swimtime="00:02:45.91" resultid="3013" heatid="9098" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:17.75" />
                    <SPLIT distance="150" swimtime="00:02:01.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="208" reactiontime="+101" swimtime="00:05:58.22" resultid="3014" heatid="9186" lane="9" entrytime="00:06:02.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:21.23" />
                    <SPLIT distance="150" swimtime="00:02:06.49" />
                    <SPLIT distance="200" swimtime="00:02:52.43" />
                    <SPLIT distance="250" swimtime="00:03:39.43" />
                    <SPLIT distance="300" swimtime="00:04:26.18" />
                    <SPLIT distance="350" swimtime="00:05:13.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="3015">
              <RESULTS>
                <RESULT eventid="1239" points="202" reactiontime="+103" swimtime="00:03:25.33" resultid="3016" heatid="8974" lane="9" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                    <SPLIT distance="100" swimtime="00:01:37.19" />
                    <SPLIT distance="150" swimtime="00:02:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="234" reactiontime="+106" swimtime="00:01:30.15" resultid="3017" heatid="9047" lane="8" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="243" reactiontime="+98" swimtime="00:00:40.46" resultid="3018" heatid="9164" lane="7" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="2991">
              <RESULTS>
                <RESULT eventid="1079" points="111" reactiontime="+106" swimtime="00:00:42.05" resultid="2992" heatid="8898" lane="9" entrytime="00:00:38.50" />
                <RESULT eventid="1113" points="92" reactiontime="+121" swimtime="00:04:02.39" resultid="2993" heatid="8922" lane="7" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.59" />
                    <SPLIT distance="100" swimtime="00:02:01.30" />
                    <SPLIT distance="150" swimtime="00:03:07.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="83" reactiontime="+92" swimtime="00:00:50.86" resultid="2994" heatid="8956" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1307" points="114" reactiontime="+112" swimtime="00:01:44.22" resultid="2995" heatid="9009" lane="4" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="134" reactiontime="+114" swimtime="00:01:48.45" resultid="2996" heatid="9045" lane="2" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="96" reactiontime="+116" swimtime="00:00:47.55" resultid="2997" heatid="9061" lane="7" entrytime="00:00:46.50" />
                <RESULT eventid="1613" points="67" reactiontime="+111" swimtime="00:01:58.94" resultid="2998" heatid="9129" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="160" reactiontime="+106" swimtime="00:00:46.42" resultid="2999" heatid="9162" lane="5" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Hanka" gender="F" lastname="Kania" nation="POL" athleteid="3000">
              <RESULTS>
                <RESULT eventid="1096" points="154" reactiontime="+115" swimtime="00:03:47.16" resultid="3001" heatid="8917" lane="2" entrytime="00:03:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.73" />
                    <SPLIT distance="100" swimtime="00:01:49.37" />
                    <SPLIT distance="150" swimtime="00:02:52.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="193" reactiontime="+115" swimtime="00:03:52.77" resultid="3002" heatid="8968" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                    <SPLIT distance="100" swimtime="00:01:50.42" />
                    <SPLIT distance="150" swimtime="00:02:51.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="151" reactiontime="+112" swimtime="00:01:46.47" resultid="3003" heatid="9002" lane="3" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="187" reactiontime="+108" swimtime="00:01:48.92" resultid="3004" heatid="9038" lane="2" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="118" reactiontime="+114" swimtime="00:00:49.61" resultid="3005" heatid="9055" lane="8" entrytime="00:00:49.00" />
                <RESULT eventid="1595" points="109" reactiontime="+105" swimtime="00:01:53.99" resultid="3006" heatid="9124" lane="3" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="198" reactiontime="+112" swimtime="00:00:49.41" resultid="3007" heatid="9153" lane="3" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="Mikołajczyk" nation="POL" athleteid="3019">
              <RESULTS>
                <RESULT eventid="1113" points="115" reactiontime="+99" swimtime="00:03:45.13" resultid="3020" heatid="8923" lane="0" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.31" />
                    <SPLIT distance="100" swimtime="00:01:53.38" />
                    <SPLIT distance="150" swimtime="00:02:53.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="133" reactiontime="+104" swimtime="00:03:55.56" resultid="3021" heatid="8972" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.60" />
                    <SPLIT distance="100" swimtime="00:01:53.25" />
                    <SPLIT distance="150" swimtime="00:02:55.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="72" reactiontime="+103" swimtime="00:04:19.96" resultid="3022" heatid="9026" lane="2" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.52" />
                    <SPLIT distance="100" swimtime="00:02:03.90" />
                    <SPLIT distance="150" swimtime="00:03:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="132" reactiontime="+104" swimtime="00:01:49.08" resultid="3023" heatid="9045" lane="8" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="3024" heatid="9117" lane="6" entrytime="00:08:10.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="3025" heatid="9129" lane="7" entrytime="00:02:05.00" />
                <RESULT eventid="1681" points="144" reactiontime="+103" swimtime="00:00:48.11" resultid="3026" heatid="9162" lane="0" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Barbara" gender="F" lastname="Chomicka" nation="POL" athleteid="3027">
              <RESULTS>
                <RESULT eventid="1062" points="105" reactiontime="+105" swimtime="00:00:49.14" resultid="3028" heatid="8886" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1096" points="82" reactiontime="+107" swimtime="00:04:40.28" resultid="3029" heatid="8916" lane="4" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.73" />
                    <SPLIT distance="100" swimtime="00:02:19.85" />
                    <SPLIT distance="150" swimtime="00:03:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="115" reactiontime="+72" swimtime="00:00:52.65" resultid="3030" heatid="8949" lane="0" entrytime="00:00:57.00" />
                <RESULT eventid="1324" points="46" reactiontime="+108" swimtime="00:05:31.91" resultid="3031" heatid="9023" lane="8" entrytime="00:05:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.64" />
                    <SPLIT distance="100" swimtime="00:02:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="50" reactiontime="+109" swimtime="00:01:05.88" resultid="3032" heatid="9054" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1457" points="95" reactiontime="+70" swimtime="00:02:00.30" resultid="3033" heatid="9074" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="47" reactiontime="+107" swimtime="00:02:30.76" resultid="3034" heatid="9124" lane="9" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="87" reactiontime="+73" swimtime="00:04:28.23" resultid="3035" heatid="9138" lane="5" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.12" />
                    <SPLIT distance="100" swimtime="00:02:11.64" />
                    <SPLIT distance="150" swimtime="00:04:28.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="147" reactiontime="+98" swimtime="00:02:51.48" resultid="3036" heatid="9032" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.26" />
                    <SPLIT distance="100" swimtime="00:01:32.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2991" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="3015" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3019" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3008" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="5111" name="GKS Tychy">
          <CONTACT city="Tychy" email="guz166@wp.pl" internet="www.tyskifan.pl" name="Mróz Marek" phone="782-985-239" street="Gen. Ch. De Gaulle&apos;A 2" zip="43-100" />
          <ATHLETES>
            <ATHLETE birthdate="1983-05-05" firstname="Marek" gender="M" lastname="Mróz" nation="POL" athleteid="5115">
              <RESULTS>
                <RESULT eventid="1079" points="508" reactiontime="+71" swimtime="00:00:25.38" resultid="5116" heatid="8911" lane="5" entrytime="00:00:26.50" />
                <RESULT eventid="1273" points="508" reactiontime="+82" swimtime="00:00:56.29" resultid="5117" heatid="8999" lane="8" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="483" reactiontime="+75" swimtime="00:00:27.77" resultid="5118" heatid="9071" lane="5" entrytime="00:00:27.73" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="5119" heatid="9104" lane="7" entrytime="00:02:10.00" />
                <RESULT eventid="1613" points="422" reactiontime="+86" swimtime="00:01:04.56" resultid="5120" heatid="9135" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-16" firstname="Michał" gender="M" lastname="Spławiński" nation="POL" athleteid="5112" />
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1775" name="GVT">
          <ATHLETES>
            <ATHLETE birthdate="1979-09-26" firstname="Łukasz" gender="M" lastname="Malaczewski" nation="POL" athleteid="1770">
              <RESULTS>
                <RESULT eventid="1079" points="529" reactiontime="+75" swimtime="00:00:25.05" resultid="1771" heatid="8912" lane="5" entrytime="00:00:26.30" />
                <RESULT eventid="1205" points="365" reactiontime="+70" swimtime="00:00:31.07" resultid="1772" heatid="8963" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1273" points="512" reactiontime="+85" swimtime="00:00:56.17" resultid="1773" heatid="8998" lane="1" entrytime="00:00:59.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="422" reactiontime="+82" swimtime="00:00:29.05" resultid="1774" heatid="9070" lane="0" entrytime="00:00:29.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3175" name="IKS Konstancin">
          <CONTACT name="Juchno" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" athleteid="3176">
              <RESULTS>
                <RESULT eventid="1079" points="415" reactiontime="+73" swimtime="00:00:27.16" resultid="3177" heatid="8908" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1113" points="326" reactiontime="+82" swimtime="00:02:39.28" resultid="3178" heatid="8927" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:15.64" />
                    <SPLIT distance="150" swimtime="00:02:03.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="418" reactiontime="+79" swimtime="00:01:00.09" resultid="3179" heatid="8997" lane="0" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="212" reactiontime="+82" swimtime="00:03:01.92" resultid="3180" heatid="9029" lane="9" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:23.33" />
                    <SPLIT distance="150" swimtime="00:02:10.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="307" reactiontime="+87" swimtime="00:01:22.35" resultid="3181" heatid="9047" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="388" reactiontime="+83" swimtime="00:02:16.15" resultid="3182" heatid="9102" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:05.63" />
                    <SPLIT distance="150" swimtime="00:01:41.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-03" firstname="Rafal" gender="M" lastname="Juchno" nation="POL" license="103714700079" athleteid="4939">
              <RESULTS>
                <RESULT eventid="1079" points="364" reactiontime="+91" swimtime="00:00:28.37" resultid="4940" heatid="8907" lane="0" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="343" reactiontime="+95" swimtime="00:01:04.18" resultid="4941" heatid="8994" lane="2" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="274" reactiontime="+94" swimtime="00:01:25.56" resultid="4942" heatid="9049" lane="7" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="262" reactiontime="+101" swimtime="00:02:35.17" resultid="4943" heatid="9099" lane="3" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:14.59" />
                    <SPLIT distance="150" swimtime="00:01:57.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" region="WA" clubid="2602" name="K.S.niezrzeszeni.pl">
          <CONTACT name="K.S.niezrzeszeni.pl" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="2610">
              <RESULTS>
                <RESULT eventid="1165" points="155" reactiontime="+132" swimtime="00:26:22.47" resultid="2611" heatid="8942" lane="7" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="100" swimtime="00:01:33.99" />
                    <SPLIT distance="150" swimtime="00:02:25.07" />
                    <SPLIT distance="200" swimtime="00:03:16.55" />
                    <SPLIT distance="250" swimtime="00:04:08.45" />
                    <SPLIT distance="300" swimtime="00:05:00.96" />
                    <SPLIT distance="350" swimtime="00:05:53.30" />
                    <SPLIT distance="400" swimtime="00:06:46.59" />
                    <SPLIT distance="450" swimtime="00:07:39.60" />
                    <SPLIT distance="500" swimtime="00:08:32.71" />
                    <SPLIT distance="550" swimtime="00:09:25.22" />
                    <SPLIT distance="600" swimtime="00:10:18.19" />
                    <SPLIT distance="650" swimtime="00:11:10.94" />
                    <SPLIT distance="700" swimtime="00:12:02.86" />
                    <SPLIT distance="750" swimtime="00:12:54.77" />
                    <SPLIT distance="800" swimtime="00:13:47.36" />
                    <SPLIT distance="850" swimtime="00:14:40.62" />
                    <SPLIT distance="900" swimtime="00:15:34.47" />
                    <SPLIT distance="950" swimtime="00:16:28.26" />
                    <SPLIT distance="1000" swimtime="00:17:23.60" />
                    <SPLIT distance="1050" swimtime="00:18:17.72" />
                    <SPLIT distance="1100" swimtime="00:19:12.40" />
                    <SPLIT distance="1150" swimtime="00:20:06.43" />
                    <SPLIT distance="1200" swimtime="00:21:01.21" />
                    <SPLIT distance="1250" swimtime="00:21:55.54" />
                    <SPLIT distance="1300" swimtime="00:22:50.62" />
                    <SPLIT distance="1350" swimtime="00:23:44.21" />
                    <SPLIT distance="1400" swimtime="00:24:38.75" />
                    <SPLIT distance="1450" swimtime="00:25:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="116" reactiontime="+121" swimtime="00:08:02.87" resultid="2612" heatid="9117" lane="7" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.74" />
                    <SPLIT distance="100" swimtime="00:01:58.35" />
                    <SPLIT distance="150" swimtime="00:03:08.90" />
                    <SPLIT distance="200" swimtime="00:04:20.08" />
                    <SPLIT distance="250" swimtime="00:05:21.20" />
                    <SPLIT distance="300" swimtime="00:06:22.62" />
                    <SPLIT distance="350" swimtime="00:07:14.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="149" reactiontime="+125" swimtime="00:06:40.28" resultid="2613" heatid="9184" lane="3" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.68" />
                    <SPLIT distance="100" swimtime="00:01:35.33" />
                    <SPLIT distance="150" swimtime="00:02:27.02" />
                    <SPLIT distance="200" swimtime="00:03:18.94" />
                    <SPLIT distance="250" swimtime="00:04:11.23" />
                    <SPLIT distance="300" swimtime="00:05:02.59" />
                    <SPLIT distance="350" swimtime="00:05:54.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-08-26" firstname="Małgorzata" gender="F" lastname="Piechura" nation="POL" athleteid="2614">
              <RESULTS>
                <RESULT eventid="1222" points="184" reactiontime="+115" swimtime="00:03:56.55" resultid="2615" heatid="8968" lane="7" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.42" />
                    <SPLIT distance="100" swimtime="00:01:54.08" />
                    <SPLIT distance="150" swimtime="00:02:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="121" reactiontime="+122" swimtime="00:01:54.59" resultid="2616" heatid="9002" lane="0" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="129" reactiontime="+113" swimtime="00:03:38.71" resultid="2617" heatid="9089" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.01" />
                    <SPLIT distance="100" swimtime="00:01:47.27" />
                    <SPLIT distance="150" swimtime="00:02:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="76" reactiontime="+110" swimtime="00:02:08.85" resultid="2618" heatid="9124" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="123" reactiontime="+115" swimtime="00:07:50.72" resultid="2619" heatid="9178" lane="1" entrytime="00:07:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.74" />
                    <SPLIT distance="100" swimtime="00:01:47.04" />
                    <SPLIT distance="150" swimtime="00:02:46.92" />
                    <SPLIT distance="200" swimtime="00:03:49.86" />
                    <SPLIT distance="250" swimtime="00:04:50.70" />
                    <SPLIT distance="300" swimtime="00:05:53.62" />
                    <SPLIT distance="350" swimtime="00:06:54.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="2603">
              <RESULTS>
                <RESULT eventid="1079" points="180" reactiontime="+102" swimtime="00:00:35.82" resultid="2604" heatid="8894" lane="2" />
                <RESULT eventid="1165" points="190" reactiontime="+124" swimtime="00:24:36.59" resultid="2605" heatid="8942" lane="5" entrytime="00:25:21.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="100" swimtime="00:01:30.33" />
                    <SPLIT distance="150" swimtime="00:02:18.09" />
                    <SPLIT distance="200" swimtime="00:03:07.14" />
                    <SPLIT distance="250" swimtime="00:03:56.97" />
                    <SPLIT distance="300" swimtime="00:04:46.40" />
                    <SPLIT distance="350" swimtime="00:05:36.42" />
                    <SPLIT distance="400" swimtime="00:06:26.77" />
                    <SPLIT distance="450" swimtime="00:07:16.84" />
                    <SPLIT distance="500" swimtime="00:08:06.73" />
                    <SPLIT distance="550" swimtime="00:08:56.48" />
                    <SPLIT distance="600" swimtime="00:09:46.27" />
                    <SPLIT distance="650" swimtime="00:10:37.09" />
                    <SPLIT distance="700" swimtime="00:11:27.67" />
                    <SPLIT distance="750" swimtime="00:12:18.06" />
                    <SPLIT distance="800" swimtime="00:13:08.16" />
                    <SPLIT distance="850" swimtime="00:13:58.12" />
                    <SPLIT distance="900" swimtime="00:14:47.64" />
                    <SPLIT distance="950" swimtime="00:15:37.92" />
                    <SPLIT distance="1000" swimtime="00:16:27.35" />
                    <SPLIT distance="1050" swimtime="00:17:17.41" />
                    <SPLIT distance="1100" swimtime="00:18:07.23" />
                    <SPLIT distance="1150" swimtime="00:18:57.69" />
                    <SPLIT distance="1200" swimtime="00:19:47.41" />
                    <SPLIT distance="1250" swimtime="00:20:36.71" />
                    <SPLIT distance="1300" swimtime="00:21:25.53" />
                    <SPLIT distance="1350" swimtime="00:22:15.10" />
                    <SPLIT distance="1400" swimtime="00:23:04.06" />
                    <SPLIT distance="1450" swimtime="00:23:52.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="154" reactiontime="+66" swimtime="00:00:41.40" resultid="2606" heatid="8958" lane="1" entrytime="00:00:40.20" />
                <RESULT eventid="1307" points="154" reactiontime="+122" swimtime="00:01:34.40" resultid="2607" heatid="9011" lane="0" entrytime="00:01:30.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="165" reactiontime="+66" swimtime="00:01:29.07" resultid="2608" heatid="9081" lane="4" entrytime="00:01:28.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="174" reactiontime="+69" swimtime="00:03:09.87" resultid="2609" heatid="9146" lane="6" entrytime="00:03:10.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:21.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KS WAR" nation="POL" region="WIE" clubid="4520" name="Klub Sportowy Warta Poznań">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Thiem Jacek" state="WIE" street="Os. Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1957-10-01" firstname="Rusłana" gender="F" lastname="Dembecka" nation="POL" license="100115600353" athleteid="6874">
              <RESULTS>
                <RESULT eventid="1222" points="137" reactiontime="+120" swimtime="00:04:20.57" resultid="6875" heatid="8967" lane="3" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.23" />
                    <SPLIT distance="100" swimtime="00:02:08.08" />
                    <SPLIT distance="150" swimtime="00:03:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="143" reactiontime="+111" swimtime="00:01:59.18" resultid="6876" heatid="9038" lane="1" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="166" reactiontime="+104" swimtime="00:00:52.33" resultid="6877" heatid="9153" lane="6" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-23" firstname="Przemysław" gender="M" lastname="Kuca" nation="POL" license="S00115200198" athleteid="6902">
              <RESULTS>
                <RESULT eventid="1079" points="583" reactiontime="+69" swimtime="00:00:24.25" resultid="6903" heatid="8914" lane="3" entrytime="00:00:24.80" />
                <RESULT eventid="1113" points="587" reactiontime="+70" swimtime="00:02:10.89" resultid="6904" heatid="8931" lane="5" entrytime="00:02:11.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="150" swimtime="00:01:42.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="589" reactiontime="+69" swimtime="00:00:53.61" resultid="6905" heatid="9000" lane="3" entrytime="00:00:52.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="639" reactiontime="+70" swimtime="00:02:06.02" resultid="6906" heatid="9030" lane="4" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="150" swimtime="00:01:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="603" reactiontime="+73" swimtime="00:01:57.61" resultid="6907" heatid="9106" lane="6" entrytime="00:01:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                    <SPLIT distance="100" swimtime="00:00:57.91" />
                    <SPLIT distance="150" swimtime="00:01:28.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="592" reactiontime="+73" swimtime="00:04:40.34" resultid="6908" heatid="9122" lane="4" entrytime="00:04:38.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                    <SPLIT distance="100" swimtime="00:01:00.11" />
                    <SPLIT distance="150" swimtime="00:01:37.64" />
                    <SPLIT distance="200" swimtime="00:02:15.00" />
                    <SPLIT distance="250" swimtime="00:02:56.76" />
                    <SPLIT distance="300" swimtime="00:03:38.54" />
                    <SPLIT distance="350" swimtime="00:04:10.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="565" reactiontime="+69" swimtime="00:00:58.56" resultid="6909" heatid="9137" lane="8" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="594" reactiontime="+72" swimtime="00:04:12.49" resultid="6910" heatid="9192" lane="5" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                    <SPLIT distance="100" swimtime="00:01:00.38" />
                    <SPLIT distance="150" swimtime="00:01:32.79" />
                    <SPLIT distance="200" swimtime="00:02:05.44" />
                    <SPLIT distance="250" swimtime="00:02:37.77" />
                    <SPLIT distance="300" swimtime="00:03:10.04" />
                    <SPLIT distance="350" swimtime="00:03:41.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="Tomaszewski" nation="POL" athleteid="6887">
              <RESULTS>
                <RESULT eventid="1079" points="447" reactiontime="+80" swimtime="00:00:26.49" resultid="6888" heatid="8910" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="1205" points="375" reactiontime="+65" swimtime="00:00:30.80" resultid="6889" heatid="8963" lane="2" entrytime="00:00:30.60" />
                <RESULT eventid="1474" points="459" reactiontime="+73" swimtime="00:01:03.44" resultid="6890" heatid="9085" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="6891" heatid="9100" lane="2" entrytime="00:02:30.00" />
                <RESULT eventid="1647" points="415" reactiontime="+74" swimtime="00:02:22.25" resultid="6892" heatid="9148" lane="6" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:09.07" />
                    <SPLIT distance="150" swimtime="00:01:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="6893" heatid="9187" lane="2" entrytime="00:05:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" license="100115700346" athleteid="6854">
              <RESULTS>
                <RESULT eventid="1165" points="322" reactiontime="+93" swimtime="00:20:39.44" resultid="6855" heatid="8946" lane="2" entrytime="00:20:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:55.14" />
                    <SPLIT distance="200" swimtime="00:02:35.02" />
                    <SPLIT distance="250" swimtime="00:03:15.61" />
                    <SPLIT distance="350" swimtime="00:05:16.95" />
                    <SPLIT distance="400" swimtime="00:05:57.40" />
                    <SPLIT distance="450" swimtime="00:06:38.15" />
                    <SPLIT distance="500" swimtime="00:07:19.00" />
                    <SPLIT distance="550" swimtime="00:07:59.88" />
                    <SPLIT distance="650" swimtime="00:08:41.09" />
                    <SPLIT distance="700" swimtime="00:09:22.49" />
                    <SPLIT distance="750" swimtime="00:10:04.11" />
                    <SPLIT distance="800" swimtime="00:10:45.94" />
                    <SPLIT distance="850" swimtime="00:11:27.44" />
                    <SPLIT distance="900" swimtime="00:12:09.49" />
                    <SPLIT distance="950" swimtime="00:12:51.74" />
                    <SPLIT distance="1000" swimtime="00:13:34.39" />
                    <SPLIT distance="1050" swimtime="00:14:17.05" />
                    <SPLIT distance="1100" swimtime="00:14:59.75" />
                    <SPLIT distance="1150" swimtime="00:15:42.53" />
                    <SPLIT distance="1200" swimtime="00:16:25.35" />
                    <SPLIT distance="1250" swimtime="00:17:08.18" />
                    <SPLIT distance="1300" swimtime="00:17:51.43" />
                    <SPLIT distance="1350" swimtime="00:18:34.31" />
                    <SPLIT distance="1400" swimtime="00:19:17.56" />
                    <SPLIT distance="1450" swimtime="00:19:59.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="320" reactiontime="+76" swimtime="00:00:32.47" resultid="6856" heatid="8960" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1307" points="310" reactiontime="+82" swimtime="00:01:14.78" resultid="6857" heatid="9016" lane="9" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="306" reactiontime="+74" swimtime="00:01:12.57" resultid="6858" heatid="9084" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="298" reactiontime="+77" swimtime="00:02:38.81" resultid="6859" heatid="9148" lane="2" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.09" />
                    <SPLIT distance="150" swimtime="00:01:59.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" license="100115600357" athleteid="6843">
              <RESULTS>
                <RESULT eventid="1147" points="234" swimtime="00:12:57.72" resultid="6844" heatid="8938" lane="0" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                    <SPLIT distance="100" swimtime="00:01:26.43" />
                    <SPLIT distance="150" swimtime="00:02:13.74" />
                    <SPLIT distance="200" swimtime="00:03:01.29" />
                    <SPLIT distance="250" swimtime="00:03:49.78" />
                    <SPLIT distance="300" swimtime="00:04:39.42" />
                    <SPLIT distance="350" swimtime="00:05:29.16" />
                    <SPLIT distance="400" swimtime="00:06:19.84" />
                    <SPLIT distance="450" swimtime="00:07:10.16" />
                    <SPLIT distance="500" swimtime="00:08:00.28" />
                    <SPLIT distance="550" swimtime="00:08:50.47" />
                    <SPLIT distance="600" swimtime="00:09:40.54" />
                    <SPLIT distance="650" swimtime="00:10:30.42" />
                    <SPLIT distance="700" swimtime="00:11:20.71" />
                    <SPLIT distance="750" swimtime="00:12:10.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="232" swimtime="00:01:22.94" resultid="6845" heatid="8981" lane="0" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="244" swimtime="00:02:57.18" resultid="6846" heatid="9090" lane="3" entrytime="00:03:02.00" />
                <RESULT eventid="1721" points="233" swimtime="00:06:20.70" resultid="6847" heatid="9179" lane="2" entrytime="00:06:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:01:26.32" />
                    <SPLIT distance="150" swimtime="00:02:12.65" />
                    <SPLIT distance="200" swimtime="00:03:00.55" />
                    <SPLIT distance="250" swimtime="00:03:50.48" />
                    <SPLIT distance="300" swimtime="00:04:41.53" />
                    <SPLIT distance="350" swimtime="00:05:32.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" license="100115700354" athleteid="6878">
              <RESULTS>
                <RESULT eventid="1113" points="472" reactiontime="+72" swimtime="00:02:20.72" resultid="6879" heatid="8931" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                    <SPLIT distance="150" swimtime="00:01:47.74" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1165" points="538" reactiontime="+79" swimtime="00:17:25.16" resultid="6880" heatid="8947" lane="4" entrytime="00:17:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:01:06.96" />
                    <SPLIT distance="150" swimtime="00:01:41.98" />
                    <SPLIT distance="200" swimtime="00:02:17.04" />
                    <SPLIT distance="250" swimtime="00:02:52.32" />
                    <SPLIT distance="300" swimtime="00:03:27.74" />
                    <SPLIT distance="350" swimtime="00:04:02.90" />
                    <SPLIT distance="400" swimtime="00:04:38.51" />
                    <SPLIT distance="450" swimtime="00:05:13.63" />
                    <SPLIT distance="500" swimtime="00:05:49.21" />
                    <SPLIT distance="550" swimtime="00:06:24.88" />
                    <SPLIT distance="600" swimtime="00:07:00.57" />
                    <SPLIT distance="650" swimtime="00:07:35.73" />
                    <SPLIT distance="700" swimtime="00:08:10.86" />
                    <SPLIT distance="750" swimtime="00:08:46.27" />
                    <SPLIT distance="800" swimtime="00:09:21.47" />
                    <SPLIT distance="850" swimtime="00:09:56.71" />
                    <SPLIT distance="900" swimtime="00:10:31.59" />
                    <SPLIT distance="950" swimtime="00:11:06.52" />
                    <SPLIT distance="1000" swimtime="00:11:41.18" />
                    <SPLIT distance="1050" swimtime="00:12:16.11" />
                    <SPLIT distance="1100" swimtime="00:12:51.28" />
                    <SPLIT distance="1150" swimtime="00:13:26.12" />
                    <SPLIT distance="1200" swimtime="00:14:00.97" />
                    <SPLIT distance="1250" swimtime="00:14:35.78" />
                    <SPLIT distance="1300" swimtime="00:15:10.71" />
                    <SPLIT distance="1350" swimtime="00:15:45.30" />
                    <SPLIT distance="1400" swimtime="00:16:19.61" />
                    <SPLIT distance="1450" swimtime="00:16:53.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="493" reactiontime="+75" swimtime="00:00:56.87" resultid="6881" heatid="9000" lane="9" entrytime="00:00:56.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="490" reactiontime="+80" swimtime="00:02:17.67" resultid="6882" heatid="9030" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                    <SPLIT distance="150" swimtime="00:01:42.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="519" reactiontime="+83" swimtime="00:02:03.63" resultid="6883" heatid="9106" lane="1" entrytime="00:02:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:01.53" />
                    <SPLIT distance="150" swimtime="00:01:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="462" reactiontime="+85" swimtime="00:05:04.51" resultid="6884" heatid="9122" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:01:08.76" />
                    <SPLIT distance="150" swimtime="00:01:50.37" />
                    <SPLIT distance="200" swimtime="00:02:29.83" />
                    <SPLIT distance="250" swimtime="00:03:12.89" />
                    <SPLIT distance="300" swimtime="00:03:56.94" />
                    <SPLIT distance="350" swimtime="00:04:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="454" reactiontime="+78" swimtime="00:00:32.83" resultid="6885" heatid="9172" lane="8" entrytime="00:00:32.20" />
                <RESULT eventid="1744" points="541" reactiontime="+82" swimtime="00:04:20.35" resultid="6886" heatid="9192" lane="3" entrytime="00:04:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="100" swimtime="00:01:03.01" />
                    <SPLIT distance="150" swimtime="00:01:36.16" />
                    <SPLIT distance="200" swimtime="00:02:09.85" />
                    <SPLIT distance="250" swimtime="00:02:42.79" />
                    <SPLIT distance="300" swimtime="00:03:15.89" />
                    <SPLIT distance="350" swimtime="00:03:48.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Grażyna" gender="F" lastname="Cabaj-Drela" nation="POL" athleteid="6837">
              <RESULTS>
                <RESULT eventid="1062" points="306" reactiontime="+89" swimtime="00:00:34.46" resultid="6838" heatid="8889" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1222" points="325" reactiontime="+90" swimtime="00:03:15.53" resultid="6839" heatid="8969" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                    <SPLIT distance="100" swimtime="00:01:33.34" />
                    <SPLIT distance="150" swimtime="00:02:24.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="332" reactiontime="+87" swimtime="00:01:30.03" resultid="6840" heatid="9041" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1423" points="257" reactiontime="+90" swimtime="00:00:38.32" resultid="6841" heatid="9056" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1664" points="336" reactiontime="+87" swimtime="00:00:41.41" resultid="6842" heatid="9156" lane="6" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" license="100115700344" athleteid="6860">
              <RESULTS>
                <RESULT eventid="1113" points="255" reactiontime="+80" swimtime="00:02:52.82" resultid="6861" heatid="8926" lane="8" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:24.55" />
                    <SPLIT distance="150" swimtime="00:02:13.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="285" reactiontime="+85" swimtime="00:03:02.97" resultid="6862" heatid="8976" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:25.70" />
                    <SPLIT distance="150" swimtime="00:02:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="260" reactiontime="+84" swimtime="00:01:19.31" resultid="6863" heatid="9013" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="288" reactiontime="+79" swimtime="00:01:24.15" resultid="6864" heatid="9050" lane="9" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="281" reactiontime="+81" swimtime="00:00:38.52" resultid="6865" heatid="9166" lane="9" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="1001155700345" athleteid="6830">
              <RESULTS>
                <RESULT eventid="1113" points="187" reactiontime="+101" swimtime="00:03:11.47" resultid="6831" heatid="8924" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                    <SPLIT distance="100" swimtime="00:01:31.48" />
                    <SPLIT distance="150" swimtime="00:02:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="207" reactiontime="+108" swimtime="00:03:03.50" resultid="6832" heatid="9028" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                    <SPLIT distance="100" swimtime="00:01:28.49" />
                    <SPLIT distance="150" swimtime="00:02:15.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="182" reactiontime="+99" swimtime="00:00:38.43" resultid="6833" heatid="9063" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1578" points="179" reactiontime="+111" swimtime="00:06:57.26" resultid="6834" heatid="9118" lane="2" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                    <SPLIT distance="100" swimtime="00:01:36.10" />
                    <SPLIT distance="150" swimtime="00:02:35.18" />
                    <SPLIT distance="200" swimtime="00:03:31.86" />
                    <SPLIT distance="250" swimtime="00:04:32.48" />
                    <SPLIT distance="300" swimtime="00:05:30.38" />
                    <SPLIT distance="350" swimtime="00:06:15.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="217" reactiontime="+101" swimtime="00:01:20.53" resultid="6835" heatid="9131" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="203" reactiontime="+108" swimtime="00:06:00.75" resultid="6836" heatid="9186" lane="6" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:01:26.92" />
                    <SPLIT distance="150" swimtime="00:02:13.34" />
                    <SPLIT distance="200" swimtime="00:02:59.95" />
                    <SPLIT distance="250" swimtime="00:03:46.55" />
                    <SPLIT distance="300" swimtime="00:04:33.12" />
                    <SPLIT distance="350" swimtime="00:05:18.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-22" firstname="Małgorzata" gender="F" lastname="Putowska" nation="POL" athleteid="6866">
              <RESULTS>
                <RESULT eventid="1062" points="180" reactiontime="+125" swimtime="00:00:41.14" resultid="6867" heatid="8886" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="1187" points="123" reactiontime="+86" swimtime="00:00:51.51" resultid="6868" heatid="8949" lane="3" entrytime="00:00:49.00" />
                <RESULT eventid="1324" points="84" reactiontime="+124" swimtime="00:04:32.39" resultid="6869" heatid="9023" lane="7" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.65" />
                    <SPLIT distance="100" swimtime="00:02:04.65" />
                    <SPLIT distance="150" swimtime="00:03:18.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="166" reactiontime="+123" swimtime="00:01:53.31" resultid="6870" heatid="9038" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="122" reactiontime="+133" swimtime="00:08:42.66" resultid="6871" heatid="9113" lane="2" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.96" />
                    <SPLIT distance="150" swimtime="00:04:19.48" />
                    <SPLIT distance="200" swimtime="00:05:26.86" />
                    <SPLIT distance="250" swimtime="00:06:34.02" />
                    <SPLIT distance="300" swimtime="00:07:37.20" />
                    <SPLIT distance="350" swimtime="00:08:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="123" reactiontime="+83" swimtime="00:03:59.49" resultid="6872" heatid="9139" lane="8" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.15" />
                    <SPLIT distance="100" swimtime="00:01:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="216" reactiontime="+129" swimtime="00:00:47.99" resultid="6873" heatid="9154" lane="2" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-03-24" firstname="Paulina" gender="F" lastname="Danielska" nation="POL" athleteid="6894">
              <RESULTS>
                <RESULT eventid="1256" points="240" reactiontime="+94" swimtime="00:01:22.00" resultid="6895" heatid="8980" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="212" reactiontime="+95" swimtime="00:03:05.77" resultid="6896" heatid="9090" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                    <SPLIT distance="100" swimtime="00:01:27.22" />
                    <SPLIT distance="150" swimtime="00:02:16.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-22" firstname="Piotr" gender="M" lastname="Burzyński" nation="POL" athleteid="6848">
              <RESULTS>
                <RESULT eventid="1165" points="191" reactiontime="+127" swimtime="00:24:34.83" resultid="6849" heatid="8944" lane="8" entrytime="00:22:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:24.86" />
                    <SPLIT distance="150" swimtime="00:02:11.06" />
                    <SPLIT distance="200" swimtime="00:02:57.60" />
                    <SPLIT distance="250" swimtime="00:03:44.54" />
                    <SPLIT distance="300" swimtime="00:04:32.67" />
                    <SPLIT distance="350" swimtime="00:05:20.46" />
                    <SPLIT distance="400" swimtime="00:06:08.72" />
                    <SPLIT distance="450" swimtime="00:06:57.12" />
                    <SPLIT distance="500" swimtime="00:07:47.21" />
                    <SPLIT distance="550" swimtime="00:08:36.71" />
                    <SPLIT distance="600" swimtime="00:09:25.39" />
                    <SPLIT distance="650" swimtime="00:10:14.58" />
                    <SPLIT distance="700" swimtime="00:11:03.79" />
                    <SPLIT distance="750" swimtime="00:11:53.52" />
                    <SPLIT distance="800" swimtime="00:12:43.49" />
                    <SPLIT distance="850" swimtime="00:13:32.72" />
                    <SPLIT distance="900" swimtime="00:14:22.14" />
                    <SPLIT distance="950" swimtime="00:15:12.27" />
                    <SPLIT distance="1000" swimtime="00:16:02.68" />
                    <SPLIT distance="1050" swimtime="00:16:53.13" />
                    <SPLIT distance="1100" swimtime="00:17:43.00" />
                    <SPLIT distance="1150" swimtime="00:18:33.75" />
                    <SPLIT distance="1200" swimtime="00:19:25.27" />
                    <SPLIT distance="1250" swimtime="00:20:15.70" />
                    <SPLIT distance="1300" swimtime="00:21:06.94" />
                    <SPLIT distance="1350" swimtime="00:21:58.80" />
                    <SPLIT distance="1400" swimtime="00:22:50.72" />
                    <SPLIT distance="1450" swimtime="00:23:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="99" reactiontime="+119" swimtime="00:03:54.38" resultid="6850" heatid="9027" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.57" />
                    <SPLIT distance="100" swimtime="00:01:52.79" />
                    <SPLIT distance="150" swimtime="00:02:54.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="6851" heatid="9098" lane="7" entrytime="00:02:47.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="6852" heatid="9118" lane="6" entrytime="00:07:07.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="6853" heatid="9186" lane="7" entrytime="00:05:57.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-02" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" license="100115700350" athleteid="6897">
              <RESULTS>
                <RESULT eventid="1079" points="406" reactiontime="+77" swimtime="00:00:27.36" resultid="6898" heatid="8908" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="418" reactiontime="+76" swimtime="00:01:00.09" resultid="6899" heatid="8996" lane="6" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="414" reactiontime="+82" swimtime="00:02:13.32" resultid="6900" heatid="9103" lane="3" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:04.67" />
                    <SPLIT distance="150" swimtime="00:01:39.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="399" reactiontime="+83" swimtime="00:04:48.07" resultid="6901" heatid="9190" lane="2" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:47.14" />
                    <SPLIT distance="200" swimtime="00:02:24.12" />
                    <SPLIT distance="250" swimtime="00:03:00.81" />
                    <SPLIT distance="300" swimtime="00:03:37.11" />
                    <SPLIT distance="350" swimtime="00:04:13.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="417" reactiontime="+72" swimtime="00:02:01.14" resultid="6914" heatid="9034" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:01.53" />
                    <SPLIT distance="150" swimtime="00:01:32.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6887" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="6878" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="6897" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="6854" number="4" reactiontime="+80" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1548" points="443" reactiontime="+79" swimtime="00:01:48.31" resultid="6918" heatid="9111" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.59" />
                    <SPLIT distance="100" swimtime="00:00:52.69" />
                    <SPLIT distance="150" swimtime="00:01:21.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6887" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="6878" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="6854" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="6897" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1358" points="163" swimtime="00:03:10.38" resultid="6913" heatid="9031" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.57" />
                    <SPLIT distance="150" swimtime="00:02:30.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6874" number="1" />
                    <RELAYPOSITION athleteid="6837" number="2" />
                    <RELAYPOSITION athleteid="6866" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="6843" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="7">
              <RESULTS>
                <RESULT eventid="1525" points="191" reactiontime="+120" swimtime="00:02:43.54" resultid="6917" heatid="9108" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                    <SPLIT distance="150" swimtime="00:02:04.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6866" number="1" reactiontime="+120" />
                    <RELAYPOSITION athleteid="6837" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="6874" number="3" reactiontime="+92" />
                    <RELAYPOSITION athleteid="6843" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="134" reactiontime="+126" swimtime="00:02:41.40" resultid="6911" heatid="8933" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:32.25" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6866" number="1" reactiontime="+126" />
                    <RELAYPOSITION athleteid="6874" number="2" />
                    <RELAYPOSITION athleteid="6848" number="3" reactiontime="+84" />
                    <RELAYPOSITION athleteid="6860" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="278" swimtime="00:02:06.55" resultid="6912" heatid="8935" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="150" swimtime="00:01:39.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6843" number="1" />
                    <RELAYPOSITION athleteid="6837" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="6887" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="6878" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="1698" points="282" reactiontime="+65" swimtime="00:02:17.87" resultid="6915" heatid="9176" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="150" swimtime="00:01:39.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6887" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="6837" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="6878" number="3" reactiontime="+20" />
                    <RELAYPOSITION athleteid="6843" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="1698" points="136" reactiontime="+87" swimtime="00:02:55.88" resultid="6916" heatid="9174" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                    <SPLIT distance="100" swimtime="00:01:35.04" />
                    <SPLIT distance="150" swimtime="00:02:15.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6830" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="6874" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="6866" number="3" reactiontime="+85" />
                    <RELAYPOSITION athleteid="6860" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00304" nation="POL" region="LBS" clubid="5972" name="KORNER Zielona Góra">
          <CONTACT name="Rzeźniewski Marian" phone="508 223-896" />
          <ATHLETES>
            <ATHLETE birthdate="1987-01-01" firstname="Andrzej" gender="M" lastname="Dubiel" nation="POL" license="100304700306" athleteid="5985">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5986" heatid="8965" lane="5" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-09-03" firstname="Jakub" gender="M" lastname="Jasiński" nation="POL" license="100304700305" athleteid="5983">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5984" heatid="8965" lane="3" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-12-12" firstname="Adam" gender="M" lastname="Plutecki" nation="POL" license="100304700306" athleteid="5978">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="5979" heatid="8915" lane="2" entrytime="00:00:23.90" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="5980" heatid="9021" lane="4" entrytime="00:00:55.50" />
                <RESULT eventid="1440" points="496" reactiontime="+94" swimtime="00:00:27.53" resultid="5981" heatid="9073" lane="5" entrytime="00:00:24.50" />
                <RESULT eventid="1681" points="531" reactiontime="+72" swimtime="00:00:31.18" resultid="5982" heatid="9172" lane="4" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-21" firstname="Marcin" gender="M" lastname="Unold" nation="POL" license="100304700304" athleteid="5973">
              <RESULTS>
                <RESULT eventid="1079" points="624" reactiontime="+73" swimtime="00:00:23.70" resultid="5974" heatid="8915" lane="1" entrytime="00:00:24.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5975" heatid="8965" lane="4" entrytime="00:00:25.50" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="5976" heatid="9087" lane="5" entrytime="00:00:58.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="5977" heatid="9150" lane="5" entrytime="00:02:03.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="5987" heatid="9112" lane="3" entrytime="00:01:38.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5973" number="1" />
                    <RELAYPOSITION athleteid="5983" number="2" />
                    <RELAYPOSITION athleteid="5978" number="3" />
                    <RELAYPOSITION athleteid="5985" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="5988" heatid="9035" lane="4" entrytime="00:01:45.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5973" number="1" />
                    <RELAYPOSITION athleteid="5978" number="2" />
                    <RELAYPOSITION athleteid="5983" number="3" />
                    <RELAYPOSITION athleteid="5985" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AWBIA" nation="POL" region="LU" clubid="3165" name="KS AZS AWF Biała Podlaska">
          <CONTACT email="zielakko@gmail.com" name="Zieliński Kamil" phone="781529483" state="LUBEL" />
          <ATHLETES>
            <ATHLETE birthdate="1989-04-27" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="3166">
              <RESULTS>
                <RESULT eventid="1113" points="415" reactiontime="+70" swimtime="00:02:26.87" resultid="3167" heatid="8930" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:49.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="362" reactiontime="+78" swimtime="00:19:51.79" resultid="3168" heatid="8947" lane="8" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="150" swimtime="00:01:52.83" />
                    <SPLIT distance="200" swimtime="00:02:31.87" />
                    <SPLIT distance="250" swimtime="00:03:11.49" />
                    <SPLIT distance="300" swimtime="00:03:51.15" />
                    <SPLIT distance="350" swimtime="00:04:31.72" />
                    <SPLIT distance="400" swimtime="00:05:12.71" />
                    <SPLIT distance="450" swimtime="00:05:53.62" />
                    <SPLIT distance="500" swimtime="00:06:34.12" />
                    <SPLIT distance="550" swimtime="00:07:14.26" />
                    <SPLIT distance="600" swimtime="00:07:55.02" />
                    <SPLIT distance="650" swimtime="00:08:35.17" />
                    <SPLIT distance="700" swimtime="00:09:15.08" />
                    <SPLIT distance="750" swimtime="00:09:55.01" />
                    <SPLIT distance="800" swimtime="00:10:35.40" />
                    <SPLIT distance="850" swimtime="00:11:15.38" />
                    <SPLIT distance="900" swimtime="00:11:56.18" />
                    <SPLIT distance="950" swimtime="00:12:36.56" />
                    <SPLIT distance="1000" swimtime="00:13:16.37" />
                    <SPLIT distance="1050" swimtime="00:13:56.25" />
                    <SPLIT distance="1100" swimtime="00:14:36.09" />
                    <SPLIT distance="1150" swimtime="00:15:16.33" />
                    <SPLIT distance="1200" swimtime="00:15:55.97" />
                    <SPLIT distance="1250" swimtime="00:16:35.94" />
                    <SPLIT distance="1300" swimtime="00:17:15.76" />
                    <SPLIT distance="1350" swimtime="00:17:55.31" />
                    <SPLIT distance="1400" swimtime="00:18:34.92" />
                    <SPLIT distance="1450" swimtime="00:19:13.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="525" reactiontime="+72" swimtime="00:02:29.27" resultid="3169" heatid="8978" lane="5" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:50.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="434" reactiontime="+76" swimtime="00:01:06.87" resultid="3170" heatid="9021" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="526" reactiontime="+70" swimtime="00:01:08.86" resultid="3171" heatid="9053" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="3172" heatid="9121" lane="6" entrytime="00:05:30.00" />
                <RESULT eventid="1681" points="550" reactiontime="+72" swimtime="00:00:30.80" resultid="3173" heatid="9172" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="3174" heatid="9183" lane="9" entrytime="00:08:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WIE" clubid="3460" name="KS Czerwonak">
          <CONTACT city="Koziegłowy" email="ewaszala59@wp.pl" name="Ewa Szała" phone="509400316" street="Osiedle Leśne 13/21" zip="62-028" />
          <ATHLETES>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="3464">
              <RESULTS>
                <RESULT eventid="1096" points="290" reactiontime="+97" swimtime="00:03:03.94" resultid="3465" heatid="8919" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:26.06" />
                    <SPLIT distance="150" swimtime="00:02:19.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="294" reactiontime="+105" swimtime="00:12:00.81" resultid="3466" heatid="8937" lane="6" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:24.94" />
                    <SPLIT distance="150" swimtime="00:02:10.50" />
                    <SPLIT distance="200" swimtime="00:02:56.64" />
                    <SPLIT distance="250" swimtime="00:03:42.16" />
                    <SPLIT distance="300" swimtime="00:04:27.62" />
                    <SPLIT distance="350" swimtime="00:05:12.90" />
                    <SPLIT distance="400" swimtime="00:05:57.99" />
                    <SPLIT distance="450" swimtime="00:06:42.97" />
                    <SPLIT distance="500" swimtime="00:07:28.68" />
                    <SPLIT distance="550" swimtime="00:08:14.74" />
                    <SPLIT distance="600" swimtime="00:08:59.25" />
                    <SPLIT distance="650" swimtime="00:09:45.55" />
                    <SPLIT distance="700" swimtime="00:10:30.60" />
                    <SPLIT distance="750" swimtime="00:11:15.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="278" reactiontime="+93" swimtime="00:01:24.22" resultid="3467" heatid="9077" lane="0" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1555" points="313" reactiontime="+95" swimtime="00:06:22.45" resultid="3468" heatid="9114" lane="5" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:01:32.44" />
                    <SPLIT distance="150" swimtime="00:02:19.61" />
                    <SPLIT distance="200" swimtime="00:03:06.53" />
                    <SPLIT distance="250" swimtime="00:04:01.11" />
                    <SPLIT distance="300" swimtime="00:04:55.24" />
                    <SPLIT distance="350" swimtime="00:05:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="278" reactiontime="+89" swimtime="00:03:02.66" resultid="3469" heatid="9140" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:01:29.28" />
                    <SPLIT distance="150" swimtime="00:02:16.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="305" reactiontime="+74" swimtime="00:05:48.07" resultid="3470" heatid="9179" lane="3" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                    <SPLIT distance="100" swimtime="00:01:21.47" />
                    <SPLIT distance="150" swimtime="00:02:05.10" />
                    <SPLIT distance="200" swimtime="00:02:49.29" />
                    <SPLIT distance="250" swimtime="00:03:33.48" />
                    <SPLIT distance="300" swimtime="00:04:17.93" />
                    <SPLIT distance="350" swimtime="00:05:02.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01910" nation="POL" region="POM" clubid="1872" name="KS Delfin Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1971-11-04" firstname="Jakub" gender="M" lastname="Mańczak" nation="POL" license="101910200065" athleteid="1873">
              <RESULTS>
                <RESULT eventid="1341" points="283" reactiontime="+83" swimtime="00:02:45.28" resultid="1874" heatid="9030" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="150" swimtime="00:02:00.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="417" reactiontime="+69" swimtime="00:00:29.16" resultid="1875" heatid="9070" lane="9" entrytime="00:00:29.50" />
                <RESULT eventid="1508" points="384" reactiontime="+74" swimtime="00:02:16.67" resultid="1876" heatid="9102" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                    <SPLIT distance="100" swimtime="00:01:05.72" />
                    <SPLIT distance="150" swimtime="00:01:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="363" reactiontime="+65" swimtime="00:01:07.88" resultid="1877" heatid="9135" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04211" nation="POL" region="11" clubid="3263" name="KS Delfin Gliwice">
          <CONTACT email="ksdelfin@op,pl" name="Cupiał Jarosław" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Teodozja" gender="F" lastname="Gdula" nation="POL" athleteid="3335">
              <RESULTS>
                <RESULT eventid="1222" points="92" reactiontime="+91" swimtime="00:04:57.17" resultid="3336" heatid="8967" lane="1" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.05" />
                    <SPLIT distance="100" swimtime="00:02:24.63" />
                    <SPLIT distance="150" swimtime="00:03:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="87" reactiontime="+87" swimtime="00:02:20.25" resultid="3337" heatid="9037" lane="3" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="94" reactiontime="+95" swimtime="00:01:03.31" resultid="3338" heatid="9152" lane="2" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-10" firstname="Barbara" gender="F" lastname="Lipowska" nation="POL" athleteid="3332">
              <RESULTS>
                <RESULT eventid="1062" points="86" reactiontime="+95" swimtime="00:00:52.56" resultid="3333" heatid="8886" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1256" points="70" reactiontime="+96" swimtime="00:02:03.41" resultid="3334" heatid="8979" lane="7" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-11-23" firstname="Jerzy" gender="M" lastname="Marciniszko" nation="POL" athleteid="3324">
              <RESULTS>
                <RESULT eventid="1079" points="39" reactiontime="+97" swimtime="00:00:59.35" resultid="3325" heatid="8895" lane="1" entrytime="00:01:00.75" />
                <RESULT eventid="1205" points="36" reactiontime="+114" swimtime="00:01:06.90" resultid="3326" heatid="8955" lane="0" entrytime="00:01:09.21" />
                <RESULT eventid="1239" points="56" reactiontime="+99" swimtime="00:05:13.74" resultid="3327" heatid="8971" lane="5" entrytime="00:05:25.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.91" />
                    <SPLIT distance="100" swimtime="00:02:26.68" />
                    <SPLIT distance="150" swimtime="00:03:49.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="61" reactiontime="+100" swimtime="00:02:20.99" resultid="3328" heatid="9044" lane="1" entrytime="00:02:21.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="28" reactiontime="+105" swimtime="00:02:40.27" resultid="3329" heatid="9079" lane="2" entrytime="00:02:47.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="33" reactiontime="+107" swimtime="00:05:30.26" resultid="3330" heatid="9143" lane="6" entrytime="00:05:54.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.92" />
                    <SPLIT distance="100" swimtime="00:02:48.76" />
                    <SPLIT distance="150" swimtime="00:04:11.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="72" reactiontime="+96" swimtime="00:01:00.60" resultid="3331" heatid="9160" lane="2" entrytime="00:01:00.67" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" region="WIE" clubid="1942" name="KS Extreme Team Oborniki">
          <CONTACT city="Oborniki" email="janwol@poczta.onet.pl" name="Wolniewicz Janusz" phone="791064667" state="WIE" street="Czarnkowska 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="1943">
              <RESULTS>
                <RESULT eventid="1165" points="121" reactiontime="+99" swimtime="00:28:34.22" resultid="1944" heatid="8941" lane="5" entrytime="00:30:01.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                    <SPLIT distance="100" swimtime="00:01:42.97" />
                    <SPLIT distance="150" swimtime="00:02:40.44" />
                    <SPLIT distance="200" swimtime="00:03:37.63" />
                    <SPLIT distance="250" swimtime="00:04:34.69" />
                    <SPLIT distance="300" swimtime="00:05:31.38" />
                    <SPLIT distance="350" swimtime="00:06:26.71" />
                    <SPLIT distance="400" swimtime="00:07:22.57" />
                    <SPLIT distance="450" swimtime="00:08:18.33" />
                    <SPLIT distance="500" swimtime="00:09:14.90" />
                    <SPLIT distance="550" swimtime="00:10:12.05" />
                    <SPLIT distance="600" swimtime="00:11:09.20" />
                    <SPLIT distance="650" swimtime="00:12:05.95" />
                    <SPLIT distance="700" swimtime="00:13:02.73" />
                    <SPLIT distance="750" swimtime="00:13:59.76" />
                    <SPLIT distance="800" swimtime="00:14:57.48" />
                    <SPLIT distance="850" swimtime="00:15:54.50" />
                    <SPLIT distance="900" swimtime="00:16:51.23" />
                    <SPLIT distance="950" swimtime="00:17:49.80" />
                    <SPLIT distance="1000" swimtime="00:18:46.92" />
                    <SPLIT distance="1050" swimtime="00:19:45.98" />
                    <SPLIT distance="1100" swimtime="00:20:45.03" />
                    <SPLIT distance="1150" swimtime="00:21:42.79" />
                    <SPLIT distance="1200" swimtime="00:22:41.48" />
                    <SPLIT distance="1250" swimtime="00:23:40.36" />
                    <SPLIT distance="1300" swimtime="00:24:40.29" />
                    <SPLIT distance="1350" swimtime="00:25:38.85" />
                    <SPLIT distance="1400" swimtime="00:26:38.66" />
                    <SPLIT distance="1450" swimtime="00:27:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="153" reactiontime="+92" swimtime="00:01:23.87" resultid="1945" heatid="8988" lane="9" entrytime="00:01:25.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="121" reactiontime="+105" swimtime="00:03:20.85" resultid="1946" heatid="9096" lane="0" entrytime="00:03:24.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:35.37" />
                    <SPLIT distance="150" swimtime="00:02:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="1947" heatid="9183" lane="7" entrytime="00:07:34.47" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="JOKRA" nation="POL" region="MAL" clubid="2596" name="KS Masters Jordan Kraków">
          <CONTACT name="Chorążak" phone="504040816" />
          <ATHLETES>
            <ATHLETE birthdate="1978-06-10" firstname="Grzegorz" gender="M" lastname="Dadej" nation="POL" athleteid="2597">
              <RESULTS>
                <RESULT eventid="1205" points="372" reactiontime="+60" swimtime="00:00:30.88" resultid="2598" heatid="8963" lane="3" entrytime="00:00:30.50" />
                <RESULT eventid="1307" points="402" reactiontime="+81" swimtime="00:01:08.59" resultid="2599" heatid="9019" lane="9" entrytime="00:01:08.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="393" reactiontime="+70" swimtime="00:01:06.79" resultid="2600" heatid="9086" lane="1" entrytime="00:01:06.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="2601" heatid="9149" lane="6" entrytime="00:02:26.81" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" region="DOL" clubid="2190" name="KS Masters Polkowice">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="ul.Kolejowa 6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-02" firstname="Pavlo" gender="M" lastname="Vechirko" nation="POL" athleteid="2191">
              <RESULTS>
                <RESULT eventid="1205" points="243" reactiontime="+84" swimtime="00:00:35.58" resultid="2192" heatid="8960" lane="0" entrytime="00:00:34.70" entrycourse="SCM" />
                <RESULT eventid="1239" points="289" reactiontime="+108" swimtime="00:03:02.08" resultid="2193" heatid="8976" lane="7" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:28.73" />
                    <SPLIT distance="150" swimtime="00:02:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="293" reactiontime="+97" swimtime="00:01:23.69" resultid="2194" heatid="9050" lane="8" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="274" reactiontime="+96" swimtime="00:01:15.30" resultid="2195" heatid="9084" lane="0" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="260" reactiontime="+102" swimtime="00:02:46.05" resultid="2196" heatid="9148" lane="1" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:21.00" />
                    <SPLIT distance="150" swimtime="00:02:03.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="289" reactiontime="+81" swimtime="00:00:38.19" resultid="2197" heatid="9166" lane="2" entrytime="00:00:38.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" clubid="7125" name="KS REKIN Świebodzice">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztof" phone="606626274" state="DOL" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1995-07-17" firstname="Agnieszka" gender="F" lastname="Gajdowska" nation="POL" license="S02001100002" athleteid="7132">
              <RESULTS>
                <RESULT eventid="1062" points="598" reactiontime="+75" swimtime="00:00:27.57" resultid="7133" heatid="8893" lane="6" entrytime="00:00:27.50" entrycourse="SCM" />
                <RESULT eventid="1187" points="438" reactiontime="+89" swimtime="00:00:33.79" resultid="7134" heatid="8952" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1256" points="569" reactiontime="+73" swimtime="00:01:01.55" resultid="7135" heatid="8984" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="449" reactiontime="+69" swimtime="00:01:21.42" resultid="7136" heatid="9041" lane="4" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="476" reactiontime="+104" swimtime="00:00:31.21" resultid="7137" heatid="9058" lane="7" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-12-22" firstname="Jacek" gender="M" lastname="Hankus" nation="POL" athleteid="7140">
              <RESULTS>
                <RESULT eventid="1079" points="448" reactiontime="+84" swimtime="00:00:26.47" resultid="7141" heatid="8906" lane="5" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1113" points="367" reactiontime="+82" swimtime="00:02:33.03" resultid="7142" heatid="8926" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                    <SPLIT distance="100" swimtime="00:01:10.17" />
                    <SPLIT distance="150" swimtime="00:01:55.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="465" reactiontime="+78" swimtime="00:00:57.99" resultid="7143" heatid="8995" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="466" reactiontime="+77" swimtime="00:01:05.34" resultid="7144" heatid="9020" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="482" reactiontime="+80" swimtime="00:00:27.80" resultid="7145" heatid="9067" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1474" points="408" reactiontime="+63" swimtime="00:01:05.96" resultid="7146" heatid="9086" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="402" reactiontime="+79" swimtime="00:01:05.60" resultid="7147" heatid="9134" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="371" reactiontime="+60" swimtime="00:02:27.61" resultid="7148" heatid="9150" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:11.02" />
                    <SPLIT distance="150" swimtime="00:01:50.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-19" firstname="Paulina" gender="F" lastname="Madeja" nation="POL" athleteid="7164">
              <RESULTS>
                <RESULT eventid="1062" points="330" reactiontime="+97" swimtime="00:00:33.60" resultid="7165" heatid="8890" lane="3" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1187" points="285" reactiontime="+87" swimtime="00:00:38.97" resultid="7166" heatid="8951" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1256" points="294" reactiontime="+96" swimtime="00:01:16.68" resultid="7167" heatid="8982" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="252" reactiontime="+96" swimtime="00:01:38.64" resultid="7168" heatid="9042" lane="9" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="234" reactiontime="+86" swimtime="00:01:29.26" resultid="7169" heatid="9077" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="7170" heatid="9156" lane="0" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-12-12" firstname="Karolina" gender="F" lastname="Jahnz" nation="POL" athleteid="7149" />
            <ATHLETE birthdate="1982-11-09" firstname="Karol" gender="M" lastname="Żemier" nation="POL" athleteid="7187">
              <RESULTS>
                <RESULT eventid="1079" points="539" reactiontime="+74" swimtime="00:00:24.89" resultid="7188" heatid="8906" lane="6" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1113" points="482" reactiontime="+75" swimtime="00:02:19.76" resultid="7189" heatid="8926" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:01:04.12" />
                    <SPLIT distance="150" swimtime="00:01:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="561" reactiontime="+77" swimtime="00:01:01.41" resultid="7190" heatid="9016" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="462" reactiontime="+77" swimtime="00:02:20.34" resultid="7191" heatid="9028" lane="5" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                    <SPLIT distance="100" swimtime="00:01:05.74" />
                    <SPLIT distance="150" swimtime="00:01:43.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="536" reactiontime="+74" swimtime="00:00:26.83" resultid="7192" heatid="9067" lane="9" entrytime="00:00:32.20" />
                <RESULT eventid="1474" points="509" reactiontime="+67" swimtime="00:01:01.26" resultid="7193" heatid="9087" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="529" reactiontime="+78" swimtime="00:00:59.86" resultid="7194" heatid="9134" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="479" reactiontime="+63" swimtime="00:02:15.55" resultid="7195" heatid="9150" lane="0" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="150" swimtime="00:01:40.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-21" firstname="Alfred" gender="M" lastname="Żemier" nation="POL" athleteid="7171">
              <RESULTS>
                <RESULT eventid="1079" points="509" reactiontime="+82" swimtime="00:00:25.36" resultid="7172" heatid="8906" lane="3" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1113" points="407" reactiontime="+81" swimtime="00:02:27.87" resultid="7173" heatid="8926" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="100" swimtime="00:01:08.10" />
                    <SPLIT distance="150" swimtime="00:01:53.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="390" reactiontime="+70" swimtime="00:00:30.40" resultid="7174" heatid="8964" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1273" points="504" reactiontime="+76" swimtime="00:00:56.45" resultid="7175" heatid="8995" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="483" reactiontime="+78" swimtime="00:00:27.77" resultid="7176" heatid="9067" lane="0" entrytime="00:00:32.20" />
                <RESULT eventid="1474" points="395" reactiontime="+64" swimtime="00:01:06.70" resultid="7177" heatid="9087" lane="8" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="361" reactiontime="+65" swimtime="00:02:28.95" resultid="7178" heatid="9149" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:50.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="7179" heatid="9165" lane="4" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-16" firstname="Filip" gender="M" lastname="Żemier" nation="POL" athleteid="7180">
              <RESULTS>
                <RESULT eventid="1079" points="461" reactiontime="+66" swimtime="00:00:26.21" resultid="7181" heatid="8907" lane="9" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1205" points="280" reactiontime="+80" swimtime="00:00:33.95" resultid="7182" heatid="8961" lane="4" entrytime="00:00:32.50" />
                <RESULT eventid="1273" points="446" reactiontime="+72" swimtime="00:00:58.78" resultid="7183" heatid="8995" lane="3" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="418" reactiontime="+69" swimtime="00:00:29.15" resultid="7184" heatid="9066" lane="4" entrytime="00:00:32.20" />
                <RESULT eventid="1613" points="456" reactiontime="+80" swimtime="00:01:02.91" resultid="7185" heatid="9134" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="351" reactiontime="+71" swimtime="00:00:35.78" resultid="7186" heatid="9166" lane="8" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-07" firstname="Ewelina" gender="F" lastname="karska" nation="POL" athleteid="7156">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="7157" heatid="8891" lane="0" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="7158" heatid="8951" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="7159" heatid="8970" lane="9" entrytime="00:03:24.00" />
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="7160" heatid="9041" lane="3" entrytime="00:01:29.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="7161" heatid="9077" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="7162" heatid="9139" lane="4" entrytime="00:03:10.00" />
                <RESULT eventid="1664" points="425" reactiontime="+67" swimtime="00:00:38.29" resultid="7163" heatid="9156" lane="9" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-20" firstname="Veronica" gender="F" lastname="Campbell-Żemier" nation="POL" athleteid="7126">
              <RESULTS>
                <RESULT eventid="1062" points="543" reactiontime="+75" swimtime="00:00:28.48" resultid="7127" heatid="8891" lane="8" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1256" points="517" reactiontime="+79" swimtime="00:01:03.54" resultid="7128" heatid="8982" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z2 - Ukończenie poszczególnych odcinków niezgodnie z przepisami o dany stylu (Time: 11:44), G-8" eventid="1290" reactiontime="+77" status="DSQ" swimtime="00:01:14.30" resultid="7129" heatid="9005" lane="9" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="451" reactiontime="+78" swimtime="00:01:21.28" resultid="7130" heatid="9041" lane="5" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="464" reactiontime="+82" swimtime="00:00:37.20" resultid="7131" heatid="9156" lane="1" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Rekin Świebodzice B" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="496" reactiontime="+68" swimtime="00:01:54.31" resultid="7529" heatid="9035" lane="2" entrytime="00:01:50.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:01.84" />
                    <SPLIT distance="150" swimtime="00:01:29.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7171" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="7187" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="7140" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="7180" number="4" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="550" reactiontime="+74" swimtime="00:01:40.77" resultid="7530" heatid="9112" lane="7" entrytime="00:01:41.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.95" />
                    <SPLIT distance="100" swimtime="00:00:50.81" />
                    <SPLIT distance="150" swimtime="00:01:15.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7187" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="7140" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="7171" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="7180" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" name="Rekin Świebodzice A" number="1">
              <RESULTS>
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="7527" heatid="9031" lane="3" entrytime="00:02:16.58">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7156" number="1" />
                    <RELAYPOSITION athleteid="7126" number="2" />
                    <RELAYPOSITION athleteid="7149" number="3" />
                    <RELAYPOSITION athleteid="7164" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="7528" heatid="9108" lane="5" entrytime="00:02:03.08">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7126" number="1" />
                    <RELAYPOSITION athleteid="7164" number="2" />
                    <RELAYPOSITION athleteid="7149" number="3" />
                    <RELAYPOSITION athleteid="7156" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="Rekin Świebodzice A" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1130" points="480" reactiontime="+77" swimtime="00:01:45.47" resultid="7523" heatid="8935" lane="4" entrytime="00:01:47.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.23" />
                    <SPLIT distance="100" swimtime="00:00:53.48" />
                    <SPLIT distance="150" swimtime="00:01:18.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7140" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="7164" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="7149" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="7180" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="368" reactiontime="+88" swimtime="00:02:06.23" resultid="7524" heatid="9176" lane="3" entrytime="00:02:01.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                    <SPLIT distance="100" swimtime="00:01:14.93" />
                    <SPLIT distance="150" swimtime="00:01:41.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7164" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="7149" number="2" reactiontime="+17" />
                    <RELAYPOSITION athleteid="7180" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="7140" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Rekin Świebodzice B" number="1">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="7525" heatid="8935" lane="5" entrytime="00:01:49.68">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7171" number="1" />
                    <RELAYPOSITION athleteid="7126" number="2" />
                    <RELAYPOSITION athleteid="7187" number="3" />
                    <RELAYPOSITION athleteid="7156" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="7526" heatid="9176" lane="5" entrytime="00:02:00.54">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7171" number="1" />
                    <RELAYPOSITION athleteid="7156" number="2" />
                    <RELAYPOSITION athleteid="7187" number="3" />
                    <RELAYPOSITION athleteid="7126" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="ZAC" clubid="3672" name="KS Triathlon Szczecin">
          <CONTACT city="Szczecin" email="martahanczewska@yahoo.pl" name="Hanczewska" phone="664935249" street="Starego Wiarusa 6" zip="71-206" />
          <ATHLETES>
            <ATHLETE birthdate="1984-10-05" firstname="Marta" gender="F" lastname="Hanczewska" nation="POL" athleteid="3680">
              <RESULTS>
                <RESULT eventid="1062" points="325" reactiontime="+89" swimtime="00:00:33.80" resultid="3681" heatid="8890" lane="9" entrytime="00:00:33.09" />
                <RESULT eventid="1256" points="307" reactiontime="+95" swimtime="00:01:15.60" resultid="3682" heatid="8982" lane="8" entrytime="00:01:14.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="327" reactiontime="+92" swimtime="00:01:30.50" resultid="3683" heatid="9040" lane="4" entrytime="00:01:32.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="345" reactiontime="+88" swimtime="00:00:41.03" resultid="3684" heatid="9157" lane="8" entrytime="00:00:40.58" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="PO" clubid="4858" name="KU AZS UAM Poznań">
          <CONTACT city="Poznań" email="kukowalazs@gmail.com" name="Kowalik" phone="603965223" state="WLKP" street="Zagajnikowa 9" zip="61-602" />
          <ATHLETES>
            <ATHLETE birthdate="1977-03-14" firstname="Jarek" gender="M" lastname="Bystry" nation="POL" athleteid="4862">
              <RESULTS>
                <RESULT eventid="1079" points="345" reactiontime="+83" swimtime="00:00:28.86" resultid="4863" heatid="8905" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1273" points="346" reactiontime="+83" swimtime="00:01:04.00" resultid="4864" heatid="8993" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="290" reactiontime="+90" swimtime="00:01:16.45" resultid="4865" heatid="9013" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="303" reactiontime="+82" swimtime="00:00:32.43" resultid="4866" heatid="9064" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1508" points="285" reactiontime="+79" swimtime="00:02:30.95" resultid="4867" heatid="9100" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:11.55" />
                    <SPLIT distance="150" swimtime="00:01:51.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="293" reactiontime="+87" swimtime="00:00:37.99" resultid="4868" heatid="9162" lane="6" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-12-27" firstname="Bartosz" gender="M" lastname="Jankowiak" nation="POL" athleteid="4883">
              <RESULTS>
                <RESULT eventid="1079" points="295" reactiontime="+77" swimtime="00:00:30.41" resultid="4884" heatid="8903" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1113" points="214" reactiontime="+82" swimtime="00:03:03.27" resultid="4885" heatid="8926" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                    <SPLIT distance="100" swimtime="00:01:24.65" />
                    <SPLIT distance="150" swimtime="00:02:19.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="257" reactiontime="+84" swimtime="00:01:10.61" resultid="4886" heatid="8991" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="235" reactiontime="+83" swimtime="00:01:22.02" resultid="4887" heatid="9013" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="4888" heatid="9047" lane="3" entrytime="00:01:30.00" />
                <RESULT eventid="1508" points="229" reactiontime="+77" swimtime="00:02:42.32" resultid="4889" heatid="9099" lane="9" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:18.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="4890" heatid="9163" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1744" points="240" reactiontime="+89" swimtime="00:05:41.20" resultid="4891" heatid="9187" lane="3" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                    <SPLIT distance="100" swimtime="00:01:19.14" />
                    <SPLIT distance="150" swimtime="00:02:02.91" />
                    <SPLIT distance="200" swimtime="00:02:47.59" />
                    <SPLIT distance="300" swimtime="00:04:15.38" />
                    <SPLIT distance="350" swimtime="00:05:00.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="Sterczyński" nation="POL" license="103315200002" athleteid="4876">
              <RESULTS>
                <RESULT eventid="1113" points="477" reactiontime="+70" swimtime="00:02:20.25" resultid="4877" heatid="8930" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                    <SPLIT distance="100" swimtime="00:01:04.84" />
                    <SPLIT distance="150" swimtime="00:01:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="388" reactiontime="+69" swimtime="00:00:30.44" resultid="4878" heatid="8964" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1307" points="515" reactiontime="+72" swimtime="00:01:03.17" resultid="4879" heatid="9020" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="416" reactiontime="+65" swimtime="00:01:05.54" resultid="4880" heatid="9087" lane="9" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="431" reactiontime="+74" swimtime="00:05:11.54" resultid="4881" heatid="9122" lane="7" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:08.44" />
                    <SPLIT distance="150" swimtime="00:01:48.85" />
                    <SPLIT distance="200" swimtime="00:02:28.19" />
                    <SPLIT distance="250" swimtime="00:03:11.48" />
                    <SPLIT distance="300" swimtime="00:03:55.48" />
                    <SPLIT distance="350" swimtime="00:04:33.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="425" reactiontime="+68" swimtime="00:02:21.11" resultid="4882" heatid="9150" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:01:06.60" />
                    <SPLIT distance="150" swimtime="00:01:43.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="Stadnik" nation="POL" license="103315100003" athleteid="4869">
              <RESULTS>
                <RESULT eventid="1062" points="624" reactiontime="+75" swimtime="00:00:27.19" resultid="4870" heatid="8893" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1187" points="502" reactiontime="+71" swimtime="00:00:32.28" resultid="4871" heatid="8953" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="1256" points="637" reactiontime="+77" swimtime="00:00:59.27" resultid="4872" heatid="8984" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="547" reactiontime="+77" swimtime="00:00:29.80" resultid="4873" heatid="9059" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1491" points="526" reactiontime="+79" swimtime="00:02:17.18" resultid="4874" heatid="9093" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                    <SPLIT distance="150" swimtime="00:01:41.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="577" reactiontime="+77" swimtime="00:00:34.58" resultid="4875" heatid="9158" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06614" nation="POL" region="MAZ" clubid="4678" name="Legia Warszawa">
          <CONTACT email="janek@plywanielegia.pl" name="Peńsko" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1990-03-22" firstname="Mariusz" gender="M" lastname="Mikołajewski" nation="POL" athleteid="4719">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1307" points="675" reactiontime="+73" swimtime="00:00:57.75" resultid="4720" heatid="9021" lane="5" entrytime="00:00:58.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-21" firstname="Krzysztof" gender="M" lastname="Spyra" nation="POL" athleteid="4686">
              <RESULTS>
                <RESULT eventid="1079" points="442" reactiontime="+74" swimtime="00:00:26.58" resultid="4687" heatid="8912" lane="1" entrytime="00:00:26.41" />
                <RESULT eventid="1273" points="458" reactiontime="+86" swimtime="00:00:58.29" resultid="4688" heatid="8998" lane="0" entrytime="00:00:59.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="429" reactiontime="+85" swimtime="00:02:11.75" resultid="4689" heatid="9101" lane="3" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="100" swimtime="00:01:03.08" />
                    <SPLIT distance="150" swimtime="00:01:37.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-11" firstname="Katarzyna" gender="F" lastname="Ptaśińska" nation="POL" athleteid="7083" />
            <ATHLETE birthdate="1987-01-01" firstname="Patryk" gender="M" lastname="Wakuła" nation="POL" athleteid="4715">
              <RESULTS>
                <RESULT eventid="1079" points="525" reactiontime="+77" swimtime="00:00:25.11" resultid="4716" heatid="8913" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="4717" heatid="8965" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="4718" heatid="9072" lane="3" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-24" firstname="Michał" gender="M" lastname="Choiński" nation="POL" athleteid="4703">
              <RESULTS>
                <RESULT eventid="1079" points="468" reactiontime="+65" swimtime="00:00:26.08" resultid="4704" heatid="8915" lane="9" entrytime="00:00:24.30" />
                <RESULT eventid="1205" points="412" reactiontime="+70" swimtime="00:00:29.85" resultid="4705" heatid="8965" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1440" points="535" reactiontime="+72" swimtime="00:00:26.84" resultid="4706" heatid="9073" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="4707" heatid="9137" lane="6" entrytime="00:00:57.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-26" firstname="Tomasz" gender="M" lastname="Wilczęga" nation="POL" athleteid="4708">
              <RESULTS>
                <RESULT eventid="1079" points="505" reactiontime="+62" swimtime="00:00:25.43" resultid="4709" heatid="8913" lane="9" entrytime="00:00:26.10" />
                <RESULT eventid="1273" points="492" reactiontime="+66" swimtime="00:00:56.89" resultid="4710" heatid="8998" lane="4" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="496" reactiontime="+65" swimtime="00:00:27.53" resultid="4711" heatid="9071" lane="9" entrytime="00:00:28.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-07" firstname="Agnieszka" gender="F" lastname="Kaczmarek" nation="POL" athleteid="4696">
              <RESULTS>
                <RESULT eventid="1062" points="437" reactiontime="+91" swimtime="00:00:30.62" resultid="4697" heatid="8892" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1096" points="417" reactiontime="+93" swimtime="00:02:43.08" resultid="4698" heatid="8920" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:02:02.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="405" reactiontime="+124" swimtime="00:00:34.68" resultid="4699" heatid="8952" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1457" points="395" reactiontime="+74" swimtime="00:01:14.97" resultid="4700" heatid="9077" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="4701" heatid="9140" lane="8" entrytime="00:03:00.00" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="4702" heatid="9157" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-03-27" firstname="Agata" gender="F" lastname="Korc" nation="POL" athleteid="4721">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1062" points="709" reactiontime="+73" swimtime="00:00:26.06" resultid="4722" heatid="8893" lane="2" entrytime="00:00:27.80" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="4723" heatid="8952" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1423" points="476" reactiontime="+71" swimtime="00:00:31.21" resultid="4724" heatid="9059" lane="7" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" athleteid="4712">
              <RESULTS>
                <RESULT eventid="1079" points="444" reactiontime="+74" swimtime="00:00:26.55" resultid="4713" heatid="8912" lane="4" entrytime="00:00:26.25" />
                <RESULT eventid="1307" points="404" reactiontime="+72" swimtime="00:01:08.50" resultid="4714" heatid="9018" lane="5" entrytime="00:01:08.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-27" firstname="Jan" gender="M" lastname="Peńsko" nation="POL" athleteid="4682">
              <RESULTS>
                <RESULT eventid="1341" points="559" reactiontime="+81" swimtime="00:02:11.74" resultid="4683" heatid="9030" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="150" swimtime="00:01:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1578" points="590" reactiontime="+81" swimtime="00:04:40.65" resultid="4684" heatid="9122" lane="3" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:01:04.63" />
                    <SPLIT distance="150" swimtime="00:01:41.89" />
                    <SPLIT distance="200" swimtime="00:02:18.30" />
                    <SPLIT distance="250" swimtime="00:02:57.46" />
                    <SPLIT distance="300" swimtime="00:03:37.23" />
                    <SPLIT distance="350" swimtime="00:04:10.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="584" reactiontime="+82" swimtime="00:00:57.95" resultid="4685" heatid="9137" lane="1" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="4690">
              <RESULTS>
                <RESULT eventid="1205" points="571" reactiontime="+63" swimtime="00:00:26.77" resultid="4691" heatid="8965" lane="7" entrytime="00:00:27.27" />
                <RESULT comment="Rekord Polski" eventid="1440" points="595" reactiontime="+77" swimtime="00:00:25.91" resultid="4692" heatid="9062" lane="3" entrytime="00:00:39.39" />
                <RESULT comment="Rekord Polski" eventid="1474" points="584" reactiontime="+63" swimtime="00:00:58.53" resultid="4693" heatid="9087" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="553" reactiontime="+90" swimtime="00:00:58.99" resultid="4694" heatid="9133" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1647" points="540" reactiontime="+66" swimtime="00:02:10.23" resultid="4695" heatid="9150" lane="3" entrytime="00:02:13.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:37.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Nie regulaminowy skład sztafety" eventid="1548" reactiontime="+67" status="DSQ" swimtime="00:01:37.94" resultid="7899" heatid="9112" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                    <SPLIT distance="100" swimtime="00:00:49.31" />
                    <SPLIT distance="150" swimtime="00:01:13.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4690" number="1" reactiontime="+67" status="DSQ" />
                    <RELAYPOSITION athleteid="4682" number="2" reactiontime="+13" status="DSQ" />
                    <RELAYPOSITION athleteid="4712" number="3" reactiontime="+29" status="DSQ" />
                    <RELAYPOSITION athleteid="4719" number="4" reactiontime="+23" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="497" reactiontime="+74" swimtime="00:01:54.24" resultid="7900" heatid="9035" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:01:01.04" />
                    <SPLIT distance="150" swimtime="00:01:28.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4719" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4712" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="4708" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="4686" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="7901" heatid="9112" lane="2" entrytime="00:01:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4719" number="1" />
                    <RELAYPOSITION athleteid="4686" number="2" />
                    <RELAYPOSITION athleteid="4712" number="3" />
                    <RELAYPOSITION athleteid="4708" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="7902" heatid="9035" lane="6" entrytime="00:01:50.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4682" number="1" />
                    <RELAYPOSITION athleteid="4703" number="2" />
                    <RELAYPOSITION athleteid="4686" number="3" />
                    <RELAYPOSITION athleteid="4719" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1130" points="460" reactiontime="+76" swimtime="00:01:46.98" resultid="7903" heatid="8932" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                    <SPLIT distance="100" swimtime="00:00:57.53" />
                    <SPLIT distance="150" swimtime="00:01:22.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4721" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4696" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4708" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4690" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="LICHE" nation="POL" region="LBL" clubid="7216" name="Lider Chełm">
          <ATHLETES>
            <ATHLETE birthdate="1989-08-19" firstname="Agnieszka" gender="F" lastname="Kargol" nation="POL" license="100403100009" athleteid="7217">
              <RESULTS>
                <RESULT eventid="1187" points="558" reactiontime="+67" swimtime="00:00:31.18" resultid="7218" heatid="8953" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1290" points="506" reactiontime="+80" swimtime="00:01:11.12" resultid="7219" heatid="9007" lane="7" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="600" reactiontime="+80" swimtime="00:00:28.90" resultid="7220" heatid="9059" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1457" points="505" reactiontime="+70" swimtime="00:01:09.07" resultid="7221" heatid="9078" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="498" reactiontime="+72" swimtime="00:02:30.34" resultid="7222" heatid="9141" lane="3" entrytime="00:02:35.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:13.52" />
                    <SPLIT distance="150" swimtime="00:01:52.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="423" reactiontime="+79" swimtime="00:00:38.34" resultid="7223" heatid="9156" lane="7" entrytime="00:00:42.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1948" name="Masters Białystok">
          <CONTACT email="mbzgloszenia@gmail.pl" name="DOMINIKA MICHALIK" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="1949">
              <RESULTS>
                <RESULT eventid="1147" points="440" reactiontime="+86" swimtime="00:10:30.09" resultid="1950" heatid="8939" lane="5" entrytime="00:10:17.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                    <SPLIT distance="150" swimtime="00:01:50.06" />
                    <SPLIT distance="200" swimtime="00:02:28.65" />
                    <SPLIT distance="250" swimtime="00:03:07.88" />
                    <SPLIT distance="300" swimtime="00:03:46.89" />
                    <SPLIT distance="350" swimtime="00:04:25.90" />
                    <SPLIT distance="400" swimtime="00:05:04.98" />
                    <SPLIT distance="450" swimtime="00:05:44.52" />
                    <SPLIT distance="500" swimtime="00:06:24.15" />
                    <SPLIT distance="550" swimtime="00:07:03.99" />
                    <SPLIT distance="600" swimtime="00:07:44.58" />
                    <SPLIT distance="650" swimtime="00:08:25.19" />
                    <SPLIT distance="700" swimtime="00:09:06.27" />
                    <SPLIT distance="750" swimtime="00:09:49.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="451" reactiontime="+85" swimtime="00:01:06.47" resultid="1951" heatid="8984" lane="8" entrytime="00:01:05.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="468" reactiontime="+90" swimtime="00:02:22.61" resultid="1952" heatid="9093" lane="6" entrytime="00:02:19.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:09.43" />
                    <SPLIT distance="150" swimtime="00:01:46.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="469" reactiontime="+87" swimtime="00:05:01.66" resultid="1953" heatid="9181" lane="4" entrytime="00:04:57.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:01:50.23" />
                    <SPLIT distance="200" swimtime="00:02:28.54" />
                    <SPLIT distance="250" swimtime="00:03:07.49" />
                    <SPLIT distance="300" swimtime="00:03:46.55" />
                    <SPLIT distance="350" swimtime="00:04:24.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LBL" clubid="2261" name="Masters Chełm">
          <CONTACT city="Chełm" email="wepa56@interia.pl" name="Wepa Wieslaw" phone="663903089" state="LUBEL" street="Grunwaldzka 36" zip="22-100" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-01" firstname="Dariusz" gender="M" lastname="Rodewald" nation="POL" athleteid="2305">
              <RESULTS>
                <RESULT eventid="1079" points="94" reactiontime="+110" swimtime="00:00:44.55" resultid="2306" heatid="8894" lane="4" />
                <RESULT eventid="1205" points="72" reactiontime="+80" swimtime="00:00:53.32" resultid="2307" heatid="8954" lane="1" />
                <RESULT eventid="1307" points="74" reactiontime="+113" swimtime="00:02:00.55" resultid="2308" heatid="9008" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="68" swimtime="00:01:59.33" resultid="2309" heatid="9079" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="64" swimtime="00:04:24.58" resultid="2310" heatid="9143" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.20" />
                    <SPLIT distance="100" swimtime="00:02:09.66" />
                    <SPLIT distance="150" swimtime="00:03:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="75" reactiontime="+114" swimtime="00:00:59.62" resultid="2311" heatid="9159" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Elżbieta" gender="F" lastname="Dziwisz" nation="POL" athleteid="2349">
              <RESULTS>
                <RESULT eventid="1187" points="84" reactiontime="+96" swimtime="00:00:58.41" resultid="2350" heatid="8948" lane="6" />
                <RESULT eventid="1222" points="83" reactiontime="+115" swimtime="00:05:08.04" resultid="2351" heatid="8966" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.24" />
                    <SPLIT distance="100" swimtime="00:02:24.43" />
                    <SPLIT distance="150" swimtime="00:03:46.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="89" reactiontime="+116" swimtime="00:02:19.34" resultid="2352" heatid="9037" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="77" reactiontime="+92" swimtime="00:02:09.27" resultid="2353" heatid="9074" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="89" reactiontime="+98" swimtime="00:04:26.57" resultid="2354" heatid="9138" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.67" />
                    <SPLIT distance="100" swimtime="00:02:08.79" />
                    <SPLIT distance="150" swimtime="00:03:17.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="101" reactiontime="+106" swimtime="00:01:01.74" resultid="2355" heatid="9152" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Janusz" gender="M" lastname="Golik" nation="POL" athleteid="2312">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="2313" heatid="8921" lane="5" entrytime="00:04:30.00" />
                <RESULT eventid="1239" points="125" reactiontime="+117" swimtime="00:04:00.72" resultid="2314" heatid="8972" lane="2" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.59" />
                    <SPLIT distance="100" swimtime="00:01:57.02" />
                    <SPLIT distance="150" swimtime="00:03:00.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="60" reactiontime="+119" swimtime="00:04:36.38" resultid="2315" heatid="9026" lane="8" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.37" />
                    <SPLIT distance="100" swimtime="00:02:15.37" />
                    <SPLIT distance="150" swimtime="00:03:26.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="149" reactiontime="+112" swimtime="00:01:44.89" resultid="2316" heatid="9045" lane="6" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="94" reactiontime="+115" swimtime="00:00:47.84" resultid="2317" heatid="9061" lane="2" entrytime="00:00:46.00" />
                <RESULT eventid="1613" points="81" reactiontime="+116" swimtime="00:01:51.94" resultid="2318" heatid="9130" lane="0" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="172" reactiontime="+99" swimtime="00:00:45.33" resultid="2319" heatid="9163" lane="8" entrytime="00:00:43.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Ireneusz" gender="M" lastname="Sokołowski" nation="POL" athleteid="2298">
              <RESULTS>
                <RESULT eventid="1079" points="47" reactiontime="+142" swimtime="00:00:56.11" resultid="2299" heatid="8894" lane="3" />
                <RESULT eventid="1205" points="54" reactiontime="+133" swimtime="00:00:58.56" resultid="2300" heatid="8954" lane="6" />
                <RESULT eventid="1307" points="54" reactiontime="+130" swimtime="00:02:13.54" resultid="2301" heatid="9008" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="90" reactiontime="+143" swimtime="00:02:04.07" resultid="2302" heatid="9043" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="2303" heatid="9079" lane="1" />
                <RESULT eventid="1681" points="114" reactiontime="+124" swimtime="00:00:52.02" resultid="2304" heatid="9159" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Wieslaw" gender="M" lastname="Wepa" nation="POL" athleteid="2320">
              <RESULTS>
                <RESULT eventid="1079" points="133" reactiontime="+93" swimtime="00:00:39.66" resultid="2321" heatid="8897" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1165" points="99" reactiontime="+132" swimtime="00:30:31.92" resultid="2322" heatid="8941" lane="8" entrytime="00:34:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.65" />
                    <SPLIT distance="100" swimtime="00:01:46.46" />
                    <SPLIT distance="150" swimtime="00:03:48.62" />
                    <SPLIT distance="200" swimtime="00:04:48.25" />
                    <SPLIT distance="250" swimtime="00:06:49.46" />
                    <SPLIT distance="300" swimtime="00:07:50.98" />
                    <SPLIT distance="350" swimtime="00:08:50.43" />
                    <SPLIT distance="400" swimtime="00:09:52.07" />
                    <SPLIT distance="450" swimtime="00:10:53.90" />
                    <SPLIT distance="500" swimtime="00:11:53.16" />
                    <SPLIT distance="550" swimtime="00:12:53.81" />
                    <SPLIT distance="600" swimtime="00:13:53.72" />
                    <SPLIT distance="650" swimtime="00:14:55.58" />
                    <SPLIT distance="700" swimtime="00:15:57.36" />
                    <SPLIT distance="750" swimtime="00:16:58.56" />
                    <SPLIT distance="800" swimtime="00:17:58.89" />
                    <SPLIT distance="850" swimtime="00:18:59.68" />
                    <SPLIT distance="900" swimtime="00:20:01.07" />
                    <SPLIT distance="950" swimtime="00:21:03.20" />
                    <SPLIT distance="1000" swimtime="00:22:04.18" />
                    <SPLIT distance="1050" swimtime="00:23:06.42" />
                    <SPLIT distance="1100" swimtime="00:24:09.96" />
                    <SPLIT distance="1150" swimtime="00:25:12.90" />
                    <SPLIT distance="1200" swimtime="00:26:18.14" />
                    <SPLIT distance="1250" swimtime="00:27:22.19" />
                    <SPLIT distance="1300" swimtime="00:28:26.58" />
                    <SPLIT distance="1450" swimtime="00:29:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="141" reactiontime="+101" swimtime="00:03:51.11" resultid="2323" heatid="8972" lane="6" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.10" />
                    <SPLIT distance="100" swimtime="00:01:49.11" />
                    <SPLIT distance="150" swimtime="00:02:50.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="71" reactiontime="+99" swimtime="00:04:21.69" resultid="2324" heatid="9026" lane="0" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.12" />
                    <SPLIT distance="100" swimtime="00:01:57.70" />
                    <SPLIT distance="150" swimtime="00:03:09.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="138" reactiontime="+95" swimtime="00:01:47.43" resultid="2325" heatid="9044" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="100" reactiontime="+129" swimtime="00:08:26.48" resultid="2326" heatid="9116" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.82" />
                    <SPLIT distance="100" swimtime="00:02:02.59" />
                    <SPLIT distance="150" swimtime="00:03:15.53" />
                    <SPLIT distance="200" swimtime="00:04:29.56" />
                    <SPLIT distance="250" swimtime="00:05:29.63" />
                    <SPLIT distance="300" swimtime="00:06:34.69" />
                    <SPLIT distance="350" swimtime="00:07:31.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="160" reactiontime="+97" swimtime="00:00:46.42" resultid="2327" heatid="9161" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1744" points="90" reactiontime="+112" swimtime="00:07:52.69" resultid="2328" heatid="9182" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.22" />
                    <SPLIT distance="100" swimtime="00:01:41.29" />
                    <SPLIT distance="150" swimtime="00:02:38.66" />
                    <SPLIT distance="200" swimtime="00:03:42.25" />
                    <SPLIT distance="250" swimtime="00:04:44.78" />
                    <SPLIT distance="300" swimtime="00:05:48.11" />
                    <SPLIT distance="350" swimtime="00:06:50.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Iwona" gender="F" lastname="Chrzan" nation="POL" athleteid="2338">
              <RESULTS>
                <RESULT eventid="1222" points="146" reactiontime="+102" swimtime="00:04:15.38" resultid="2339" heatid="8966" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.93" />
                    <SPLIT distance="100" swimtime="00:02:02.29" />
                    <SPLIT distance="150" swimtime="00:03:08.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="72" reactiontime="+96" swimtime="00:02:02.25" resultid="2340" heatid="8979" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="144" reactiontime="+118" swimtime="00:01:58.92" resultid="2341" heatid="9036" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="2342" heatid="9088" lane="5" />
                <RESULT eventid="1664" points="132" reactiontime="+98" swimtime="00:00:56.52" resultid="2343" heatid="9151" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Hanna" gender="F" lastname="Wepa" nation="POL" athleteid="2329">
              <RESULTS>
                <RESULT eventid="1062" points="51" reactiontime="+136" swimtime="00:01:02.42" resultid="2330" heatid="8885" lane="5" />
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="2331" heatid="8936" lane="1" />
                <RESULT eventid="1222" points="97" reactiontime="+134" swimtime="00:04:52.56" resultid="2332" heatid="8966" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.55" />
                    <SPLIT distance="100" swimtime="00:02:22.42" />
                    <SPLIT distance="150" swimtime="00:03:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="48" reactiontime="+138" swimtime="00:02:19.98" resultid="2333" heatid="8979" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="85" reactiontime="+132" swimtime="00:02:21.31" resultid="2334" heatid="9036" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="54" reactiontime="+123" swimtime="00:04:51.91" resultid="2335" heatid="9088" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.28" />
                    <SPLIT distance="100" swimtime="00:02:24.14" />
                    <SPLIT distance="150" swimtime="00:03:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="88" reactiontime="+125" swimtime="00:01:04.71" resultid="2336" heatid="9151" lane="3" />
                <RESULT eventid="1721" points="60" reactiontime="+134" swimtime="00:09:57.76" resultid="2337" heatid="9177" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.43" />
                    <SPLIT distance="100" swimtime="00:02:20.56" />
                    <SPLIT distance="150" swimtime="00:03:36.37" />
                    <SPLIT distance="200" swimtime="00:04:51.61" />
                    <SPLIT distance="250" swimtime="00:06:08.04" />
                    <SPLIT distance="300" swimtime="00:07:25.09" />
                    <SPLIT distance="350" swimtime="00:08:41.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Piotr" gender="M" lastname="Gryciuk" nation="POL" athleteid="2262">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="2263" heatid="8907" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1113" points="332" reactiontime="+84" swimtime="00:02:38.24" resultid="2264" heatid="8928" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:02:02.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2265" heatid="8994" lane="7" entrytime="00:01:04.00" />
                <RESULT eventid="1307" points="395" reactiontime="+81" swimtime="00:01:09.02" resultid="2266" heatid="9017" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="393" reactiontime="+83" swimtime="00:00:29.76" resultid="2267" heatid="9068" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="2268" heatid="9100" lane="3" entrytime="00:02:30.00" />
                <RESULT eventid="1613" points="319" reactiontime="+81" swimtime="00:01:10.86" resultid="2269" heatid="9133" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="2270" heatid="9163" lane="4" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Dorota" gender="F" lastname="Czerniakiewicz" nation="POL" athleteid="2344">
              <RESULTS>
                <RESULT eventid="1187" points="106" reactiontime="+113" swimtime="00:00:54.10" resultid="2345" heatid="8948" lane="7" />
                <RESULT eventid="1222" points="148" reactiontime="+95" swimtime="00:04:14.25" resultid="2346" heatid="8966" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.46" />
                    <SPLIT distance="100" swimtime="00:02:03.65" />
                    <SPLIT distance="150" swimtime="00:03:09.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="144" reactiontime="+89" swimtime="00:01:58.86" resultid="2347" heatid="9037" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="146" reactiontime="+92" swimtime="00:00:54.66" resultid="2348" heatid="9151" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Leszek" gender="M" lastname="Masłowski" nation="POL" athleteid="2271">
              <RESULTS>
                <RESULT eventid="1079" points="65" reactiontime="+105" swimtime="00:00:50.35" resultid="2272" heatid="8895" lane="9" />
                <RESULT comment="Z1 - Nieprawidłowa kolejność stylów pływania (motylkowy, grzbietowy, klasyczny, dowolny) (Time: 17:28)" eventid="1113" reactiontime="+124" status="DSQ" swimtime="00:05:14.85" resultid="2273" heatid="8921" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.82" />
                    <SPLIT distance="100" swimtime="00:02:31.53" />
                    <SPLIT distance="150" swimtime="00:03:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="59" reactiontime="+123" swimtime="00:05:08.90" resultid="2274" heatid="8971" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.10" />
                    <SPLIT distance="100" swimtime="00:02:31.17" />
                    <SPLIT distance="150" swimtime="00:03:51.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="54" reactiontime="+117" swimtime="00:01:58.75" resultid="2275" heatid="8986" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="57" reactiontime="+127" swimtime="00:02:24.02" resultid="2276" heatid="9043" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="46" reactiontime="+107" swimtime="00:04:35.75" resultid="2277" heatid="9094" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.20" />
                    <SPLIT distance="100" swimtime="00:02:06.18" />
                    <SPLIT distance="150" swimtime="00:03:23.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="34" reactiontime="+97" swimtime="00:05:27.52" resultid="2278" heatid="9142" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.35" />
                    <SPLIT distance="100" swimtime="00:02:39.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="72" reactiontime="+120" swimtime="00:01:00.56" resultid="2279" heatid="9159" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Jan" gender="M" lastname="Biskup" nation="POL" athleteid="2284">
              <RESULTS>
                <RESULT eventid="1079" points="115" reactiontime="+103" swimtime="00:00:41.65" resultid="2285" heatid="8894" lane="6" />
                <RESULT eventid="1205" points="37" reactiontime="+112" swimtime="00:01:06.11" resultid="2286" heatid="8954" lane="0" />
                <RESULT eventid="1273" points="90" reactiontime="+113" swimtime="00:01:40.01" resultid="2287" heatid="8985" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="76" reactiontime="+107" swimtime="00:02:10.87" resultid="2288" heatid="9043" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="63" reactiontime="+113" swimtime="00:04:09.36" resultid="2289" heatid="9094" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.91" />
                    <SPLIT distance="100" swimtime="00:01:53.64" />
                    <SPLIT distance="150" swimtime="00:03:03.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="88" reactiontime="+108" swimtime="00:00:56.60" resultid="2290" heatid="9160" lane="9" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2291" heatid="9182" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Wosk" nation="POL" athleteid="2292">
              <RESULTS>
                <RESULT eventid="1079" points="12" reactiontime="+146" swimtime="00:01:28.32" resultid="2293" heatid="8894" lane="5" />
                <RESULT eventid="1205" reactiontime="+80" status="DNS" swimtime="00:00:00.00" resultid="2294" heatid="8954" lane="7" />
                <RESULT eventid="1273" points="12" reactiontime="+135" swimtime="00:03:12.20" resultid="2295" heatid="8985" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="6" reactiontime="+88" swimtime="00:04:17.30" resultid="2296" heatid="9079" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:01.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="13" reactiontime="+148" swimtime="00:01:45.89" resultid="2297" heatid="9159" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="53" reactiontime="+79" swimtime="00:03:59.88" resultid="2360" heatid="9032" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.37" />
                    <SPLIT distance="100" swimtime="00:01:52.54" />
                    <SPLIT distance="150" swimtime="00:02:42.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2305" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2271" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2312" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="2292" number="4" reactiontime="+193" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="51" reactiontime="+126" swimtime="00:03:42.03" resultid="2362" heatid="9109" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.01" />
                    <SPLIT distance="100" swimtime="00:01:40.12" />
                    <SPLIT distance="150" swimtime="00:02:25.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2271" number="1" reactiontime="+126" />
                    <RELAYPOSITION athleteid="2312" number="2" reactiontime="+116" />
                    <RELAYPOSITION athleteid="2305" number="3" reactiontime="+98" />
                    <RELAYPOSITION athleteid="2292" number="4" reactiontime="+116" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="139" reactiontime="+107" swimtime="00:02:54.51" resultid="2358" heatid="9032" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.30" />
                    <SPLIT distance="100" swimtime="00:01:44.41" />
                    <SPLIT distance="150" swimtime="00:02:14.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2298" number="1" reactiontime="+107" />
                    <RELAYPOSITION athleteid="2262" number="2" reactiontime="+106" />
                    <RELAYPOSITION athleteid="2284" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2320" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="2359" heatid="9109" lane="0">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2284" number="1" />
                    <RELAYPOSITION athleteid="2262" number="2" />
                    <RELAYPOSITION athleteid="2298" number="3" />
                    <RELAYPOSITION athleteid="2320" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1525" points="75" reactiontime="+104" swimtime="00:03:43.14" resultid="2356" heatid="9107" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.21" />
                    <SPLIT distance="100" swimtime="00:01:51.74" />
                    <SPLIT distance="150" swimtime="00:02:58.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2349" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="2338" number="2" reactiontime="+15" />
                    <RELAYPOSITION athleteid="2329" number="3" reactiontime="+102" />
                    <RELAYPOSITION athleteid="2344" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="59" reactiontime="+121" swimtime="00:03:31.96" resultid="2357" heatid="8932" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.50" />
                    <SPLIT distance="100" swimtime="00:01:45.27" />
                    <SPLIT distance="150" swimtime="00:02:49.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2349" number="1" reactiontime="+121" />
                    <RELAYPOSITION athleteid="2271" number="2" reactiontime="-34" />
                    <RELAYPOSITION athleteid="2329" number="3" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2320" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="118" reactiontime="+84" swimtime="00:02:48.28" resultid="2361" heatid="8932" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="100" swimtime="00:01:14.37" />
                    <SPLIT distance="150" swimtime="00:01:54.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2262" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="2344" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="2284" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2338" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="RZ" clubid="5956" name="Masters Ikar Mielec">
          <CONTACT city="CHORZELÓW" email="sebastianboicetta@gmail.com" name="SEBASTIAN BOICETTA" phone="501072284" state="PODKA" street="MALINIE 629" zip="39-331" />
          <ATHLETES>
            <ATHLETE birthdate="1975-04-01" firstname="Sebastian" gender="M" lastname="Boicetta" nation="POL" athleteid="5962">
              <RESULTS>
                <RESULT eventid="1079" points="293" reactiontime="+82" swimtime="00:00:30.48" resultid="5963" heatid="8902" lane="6" entrytime="00:00:31.40" entrycourse="SCM" />
                <RESULT eventid="1205" points="219" reactiontime="+64" swimtime="00:00:36.86" resultid="5964" heatid="8958" lane="4" entrytime="00:00:38.13" entrycourse="SCM" />
                <RESULT eventid="1307" points="246" reactiontime="+75" swimtime="00:01:20.84" resultid="5965" heatid="9014" lane="9" entrytime="00:01:19.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="212" reactiontime="+73" swimtime="00:01:21.97" resultid="5966" heatid="9082" lane="6" entrytime="00:01:21.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-18" firstname="Martyna" gender="F" lastname="Radłowska-Lewińska" nation="POL" athleteid="5967">
              <RESULTS>
                <RESULT eventid="1062" points="405" reactiontime="+95" swimtime="00:00:31.41" resultid="5968" heatid="8891" lane="2" entrytime="00:00:31.19" entrycourse="SCM" />
                <RESULT eventid="1256" points="407" reactiontime="+87" swimtime="00:01:08.81" resultid="5969" heatid="8984" lane="0" entrytime="00:01:05.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="374" reactiontime="+87" swimtime="00:01:18.65" resultid="5970" heatid="9006" lane="7" entrytime="00:01:19.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="295" reactiontime="+89" swimtime="00:00:36.62" resultid="5971" heatid="9057" lane="2" entrytime="00:00:35.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KRA" nation="POL" region="MAL" clubid="4306" name="Masters Korona Kraków">
          <CONTACT city="Kraków" email="masterskorona@wp.pl" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="Wysocka" nation="POL" athleteid="7360">
              <RESULTS>
                <RESULT eventid="1222" points="316" reactiontime="+95" swimtime="00:03:17.54" resultid="7361" heatid="8970" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                    <SPLIT distance="150" swimtime="00:02:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="317" reactiontime="+94" swimtime="00:01:31.41" resultid="7362" heatid="9041" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1664" points="345" reactiontime="+92" swimtime="00:00:41.03" resultid="7363" heatid="9156" lane="2" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="Frączek" nation="POL" athleteid="7242">
              <RESULTS>
                <RESULT eventid="1062" points="488" reactiontime="+84" swimtime="00:00:29.51" resultid="7243" heatid="8892" lane="2" entrytime="00:00:29.70" />
                <RESULT comment="Rekord Polski" eventid="1256" points="479" reactiontime="+93" swimtime="00:01:05.15" resultid="7244" heatid="8983" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="405" reactiontime="+82" swimtime="00:00:32.95" resultid="7245" heatid="9058" lane="6" entrytime="00:00:33.60" />
                <RESULT eventid="1491" points="393" reactiontime="+86" swimtime="00:02:31.14" resultid="7246" heatid="9092" lane="2" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:01:52.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-29" firstname="Jolanta" gender="F" lastname="Uczarczyk" nation="POL" athleteid="7377">
              <RESULTS>
                <RESULT eventid="1256" points="199" reactiontime="+85" swimtime="00:01:27.25" resultid="7378" heatid="8980" lane="4" entrytime="00:01:26.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="171" reactiontime="+108" swimtime="00:00:43.91" resultid="7379" heatid="9055" lane="5" entrytime="00:00:44.72" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="7229">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1062" points="502" reactiontime="+73" swimtime="00:00:29.24" resultid="7230" heatid="8892" lane="3" entrytime="00:00:29.60" />
                <RESULT eventid="1187" points="415" reactiontime="+62" swimtime="00:00:34.39" resultid="7231" heatid="8952" lane="4" entrytime="00:00:34.30" />
                <RESULT comment="Rekord Polski" eventid="1290" points="451" reactiontime="+73" swimtime="00:01:13.92" resultid="7232" heatid="9006" lane="5" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="451" reactiontime="+78" swimtime="00:01:21.27" resultid="7233" heatid="9038" lane="7" entrytime="00:01:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="434" reactiontime="+73" swimtime="00:00:32.18" resultid="7234" heatid="9058" lane="5" entrytime="00:00:32.10" />
                <RESULT comment="Rekord Polski" eventid="1664" points="544" reactiontime="+74" swimtime="00:00:35.26" resultid="7235" heatid="9158" lane="5" entrytime="00:00:35.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-16" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="7260">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="7261" heatid="8921" lane="1" />
                <RESULT eventid="1205" points="39" reactiontime="+70" swimtime="00:01:05.00" resultid="7262" heatid="8955" lane="9" entrytime="00:01:10.00" />
                <RESULT eventid="1307" points="32" reactiontime="+87" swimtime="00:02:37.99" resultid="7263" heatid="9009" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="18" reactiontime="+127" swimtime="00:01:22.93" resultid="7264" heatid="9060" lane="1" entrytime="00:01:15.00" />
                <RESULT eventid="1474" points="38" reactiontime="+86" swimtime="00:02:25.20" resultid="7265" heatid="9079" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="7266" heatid="9142" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-10-20" firstname="Janusz" gender="M" lastname="Toporski" nation="POL" athleteid="7324">
              <RESULTS>
                <RESULT eventid="1079" points="143" reactiontime="+83" swimtime="00:00:38.70" resultid="7325" heatid="8898" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1113" points="105" reactiontime="+90" swimtime="00:03:52.30" resultid="7326" heatid="8922" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.20" />
                    <SPLIT distance="100" swimtime="00:02:02.04" />
                    <SPLIT distance="150" swimtime="00:03:02.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="120" reactiontime="+104" swimtime="00:01:31.02" resultid="7327" heatid="8987" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="98" reactiontime="+106" swimtime="00:03:54.88" resultid="7328" heatid="9026" lane="1" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.94" />
                    <SPLIT distance="100" swimtime="00:01:53.13" />
                    <SPLIT distance="150" swimtime="00:02:55.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="103" reactiontime="+93" swimtime="00:00:46.43" resultid="7329" heatid="9060" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1508" points="97" reactiontime="+93" swimtime="00:03:35.63" resultid="7330" heatid="9096" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                    <SPLIT distance="100" swimtime="00:01:42.55" />
                    <SPLIT distance="150" swimtime="00:02:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="104" reactiontime="+113" swimtime="00:01:42.77" resultid="7331" heatid="9129" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="104" reactiontime="+110" swimtime="00:07:30.13" resultid="7332" heatid="9183" lane="3" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                    <SPLIT distance="100" swimtime="00:01:47.61" />
                    <SPLIT distance="150" swimtime="00:02:45.25" />
                    <SPLIT distance="200" swimtime="00:03:42.73" />
                    <SPLIT distance="250" swimtime="00:04:39.92" />
                    <SPLIT distance="300" swimtime="00:05:38.82" />
                    <SPLIT distance="350" swimtime="00:06:35.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-31" firstname="Marek" gender="M" lastname="Juza" nation="POL" athleteid="7380">
              <RESULTS>
                <RESULT eventid="1113" points="287" reactiontime="+91" swimtime="00:02:46.16" resultid="7381" heatid="8928" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:02:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="293" reactiontime="+91" swimtime="00:03:01.38" resultid="7382" heatid="8977" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:27.30" />
                    <SPLIT distance="150" swimtime="00:02:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="359" reactiontime="+94" swimtime="00:00:30.66" resultid="7383" heatid="9068" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1681" points="336" reactiontime="+88" swimtime="00:00:36.32" resultid="7384" heatid="9167" lane="4" entrytime="00:00:37.50" />
                <RESULT eventid="1744" points="233" reactiontime="+87" swimtime="00:05:44.77" resultid="7385" heatid="9191" lane="2" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:57.57" />
                    <SPLIT distance="200" swimtime="00:02:42.13" />
                    <SPLIT distance="250" swimtime="00:03:27.36" />
                    <SPLIT distance="300" swimtime="00:04:13.81" />
                    <SPLIT distance="350" swimtime="00:05:00.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-08-24" firstname="Andrzej" gender="M" lastname="Wygrzywalski" nation="POL" athleteid="7340">
              <RESULTS>
                <RESULT eventid="1079" points="200" reactiontime="+83" swimtime="00:00:34.64" resultid="7341" heatid="8900" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1165" points="181" reactiontime="+84" swimtime="00:25:01.01" resultid="7342" heatid="8942" lane="4" entrytime="00:25:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="100" swimtime="00:01:26.18" />
                    <SPLIT distance="150" swimtime="00:02:15.12" />
                    <SPLIT distance="200" swimtime="00:03:04.35" />
                    <SPLIT distance="250" swimtime="00:03:54.16" />
                    <SPLIT distance="300" swimtime="00:04:44.21" />
                    <SPLIT distance="350" swimtime="00:05:34.49" />
                    <SPLIT distance="400" swimtime="00:06:24.51" />
                    <SPLIT distance="450" swimtime="00:07:15.31" />
                    <SPLIT distance="500" swimtime="00:08:06.12" />
                    <SPLIT distance="550" swimtime="00:08:57.22" />
                    <SPLIT distance="600" swimtime="00:09:48.05" />
                    <SPLIT distance="650" swimtime="00:10:39.34" />
                    <SPLIT distance="700" swimtime="00:11:30.30" />
                    <SPLIT distance="750" swimtime="00:12:21.26" />
                    <SPLIT distance="800" swimtime="00:13:12.53" />
                    <SPLIT distance="850" swimtime="00:14:03.60" />
                    <SPLIT distance="900" swimtime="00:14:55.09" />
                    <SPLIT distance="950" swimtime="00:15:45.99" />
                    <SPLIT distance="1000" swimtime="00:16:37.46" />
                    <SPLIT distance="1050" swimtime="00:17:28.58" />
                    <SPLIT distance="1100" swimtime="00:18:19.67" />
                    <SPLIT distance="1150" swimtime="00:19:10.81" />
                    <SPLIT distance="1200" swimtime="00:20:02.03" />
                    <SPLIT distance="1250" swimtime="00:20:53.42" />
                    <SPLIT distance="1300" swimtime="00:21:43.99" />
                    <SPLIT distance="1350" swimtime="00:22:35.05" />
                    <SPLIT distance="1400" swimtime="00:23:26.15" />
                    <SPLIT distance="1450" swimtime="00:24:15.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="192" reactiontime="+80" swimtime="00:01:17.81" resultid="7343" heatid="8988" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="183" reactiontime="+89" swimtime="00:02:54.87" resultid="7344" heatid="9097" lane="0" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:23.95" />
                    <SPLIT distance="150" swimtime="00:02:10.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="181" reactiontime="+82" swimtime="00:06:15.02" resultid="7345" heatid="9185" lane="7" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:14.35" />
                    <SPLIT distance="200" swimtime="00:03:03.15" />
                    <SPLIT distance="250" swimtime="00:03:52.46" />
                    <SPLIT distance="300" swimtime="00:04:41.77" />
                    <SPLIT distance="350" swimtime="00:05:29.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="7270">
              <RESULTS>
                <RESULT eventid="1062" points="334" reactiontime="+96" swimtime="00:00:33.48" resultid="7271" heatid="8889" lane="3" entrytime="00:00:34.50" />
                <RESULT eventid="1147" points="286" reactiontime="+105" swimtime="00:12:07.38" resultid="7272" heatid="8938" lane="2" entrytime="00:12:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:22.50" />
                    <SPLIT distance="150" swimtime="00:02:07.71" />
                    <SPLIT distance="200" swimtime="00:02:53.31" />
                    <SPLIT distance="250" swimtime="00:03:39.86" />
                    <SPLIT distance="300" swimtime="00:04:27.02" />
                    <SPLIT distance="350" swimtime="00:05:13.95" />
                    <SPLIT distance="400" swimtime="00:06:00.68" />
                    <SPLIT distance="450" swimtime="00:06:47.12" />
                    <SPLIT distance="500" swimtime="00:07:34.04" />
                    <SPLIT distance="550" swimtime="00:08:20.70" />
                    <SPLIT distance="600" swimtime="00:09:07.25" />
                    <SPLIT distance="650" swimtime="00:09:53.52" />
                    <SPLIT distance="700" swimtime="00:10:39.28" />
                    <SPLIT distance="750" swimtime="00:11:25.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="306" reactiontime="+103" swimtime="00:01:15.68" resultid="7273" heatid="8981" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="198" reactiontime="+107" swimtime="00:03:25.20" resultid="7274" heatid="9023" lane="4" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:31.94" />
                    <SPLIT distance="150" swimtime="00:02:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1423" points="256" reactiontime="+94" swimtime="00:00:38.39" resultid="7275" heatid="9054" lane="7" />
                <RESULT eventid="1491" points="295" reactiontime="+88" swimtime="00:02:46.33" resultid="7276" heatid="9091" lane="5" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                    <SPLIT distance="150" swimtime="00:02:04.31" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1595" points="228" reactiontime="+93" swimtime="00:01:29.39" resultid="7277" heatid="9125" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="287" reactiontime="+100" swimtime="00:05:55.43" resultid="7278" heatid="9179" lane="4" entrytime="00:06:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:22.54" />
                    <SPLIT distance="150" swimtime="00:02:07.71" />
                    <SPLIT distance="200" swimtime="00:02:52.58" />
                    <SPLIT distance="250" swimtime="00:03:38.55" />
                    <SPLIT distance="300" swimtime="00:04:25.11" />
                    <SPLIT distance="350" swimtime="00:05:11.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-21" firstname="Adam" gender="M" lastname="Pycia" nation="POL" athleteid="7310">
              <RESULTS>
                <RESULT eventid="1239" points="219" reactiontime="+131" swimtime="00:03:19.82" resultid="7311" heatid="8974" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                    <SPLIT distance="100" swimtime="00:01:37.20" />
                    <SPLIT distance="150" swimtime="00:02:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="262" reactiontime="+95" swimtime="00:01:10.22" resultid="7312" heatid="8991" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K14 - Praca nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie) (Time: 16:34)" eventid="1406" reactiontime="+119" status="DSQ" swimtime="00:01:30.05" resultid="7313" heatid="9047" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="246" reactiontime="+105" swimtime="00:02:38.53" resultid="7314" heatid="9099" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:14.37" />
                    <SPLIT distance="150" swimtime="00:01:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="258" reactiontime="+102" swimtime="00:00:39.63" resultid="7315" heatid="9164" lane="2" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-04-07" firstname="Jacek" gender="M" lastname="Żurek" nation="POL" athleteid="7355">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="7356" heatid="8910" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="7357" heatid="8947" lane="3" entrytime="00:19:00.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="7358" heatid="8996" lane="5" entrytime="00:01:01.00" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="7359" heatid="9018" lane="0" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-12" firstname="Wojciech" gender="M" lastname="Hoffman" nation="POL" athleteid="7247">
              <RESULTS>
                <RESULT eventid="1079" points="330" reactiontime="+76" swimtime="00:00:29.29" resultid="7248" heatid="8904" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1165" points="333" reactiontime="+90" swimtime="00:20:25.73" resultid="7249" heatid="8946" lane="5" entrytime="00:20:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:01:52.59" />
                    <SPLIT distance="200" swimtime="00:02:32.09" />
                    <SPLIT distance="250" swimtime="00:03:12.14" />
                    <SPLIT distance="300" swimtime="00:03:52.40" />
                    <SPLIT distance="350" swimtime="00:04:33.20" />
                    <SPLIT distance="400" swimtime="00:05:13.99" />
                    <SPLIT distance="450" swimtime="00:05:55.14" />
                    <SPLIT distance="500" swimtime="00:06:36.43" />
                    <SPLIT distance="550" swimtime="00:07:17.73" />
                    <SPLIT distance="600" swimtime="00:07:59.31" />
                    <SPLIT distance="650" swimtime="00:08:40.75" />
                    <SPLIT distance="700" swimtime="00:09:22.10" />
                    <SPLIT distance="750" swimtime="00:10:03.54" />
                    <SPLIT distance="800" swimtime="00:10:45.07" />
                    <SPLIT distance="850" swimtime="00:11:26.49" />
                    <SPLIT distance="900" swimtime="00:12:07.95" />
                    <SPLIT distance="950" swimtime="00:12:49.46" />
                    <SPLIT distance="1000" swimtime="00:13:30.60" />
                    <SPLIT distance="1050" swimtime="00:14:12.26" />
                    <SPLIT distance="1100" swimtime="00:14:54.08" />
                    <SPLIT distance="1150" swimtime="00:15:35.94" />
                    <SPLIT distance="1200" swimtime="00:16:17.72" />
                    <SPLIT distance="1250" swimtime="00:16:59.33" />
                    <SPLIT distance="1300" swimtime="00:17:41.57" />
                    <SPLIT distance="1350" swimtime="00:18:23.84" />
                    <SPLIT distance="1400" swimtime="00:19:05.47" />
                    <SPLIT distance="1450" swimtime="00:19:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="332" reactiontime="+80" swimtime="00:01:04.88" resultid="7250" heatid="8993" lane="7" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="336" reactiontime="+78" swimtime="00:02:22.89" resultid="7251" heatid="9101" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="150" swimtime="00:01:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="334" reactiontime="+84" swimtime="00:05:05.89" resultid="7252" heatid="9189" lane="2" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:01:53.02" />
                    <SPLIT distance="200" swimtime="00:02:32.06" />
                    <SPLIT distance="250" swimtime="00:03:10.68" />
                    <SPLIT distance="300" swimtime="00:03:49.64" />
                    <SPLIT distance="350" swimtime="00:04:28.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="7346">
              <RESULTS>
                <RESULT eventid="1096" points="304" reactiontime="+87" swimtime="00:03:01.07" resultid="7347" heatid="8918" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                    <SPLIT distance="150" swimtime="00:02:18.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="313" reactiontime="+92" swimtime="00:01:23.47" resultid="7348" heatid="9004" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="294" reactiontime="+99" swimtime="00:02:46.52" resultid="7349" heatid="9091" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:01:20.15" />
                    <SPLIT distance="150" swimtime="00:02:03.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="285" reactiontime="+92" swimtime="00:06:34.67" resultid="7350" heatid="9114" lane="4" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:28.91" />
                    <SPLIT distance="150" swimtime="00:02:21.58" />
                    <SPLIT distance="200" swimtime="00:03:12.59" />
                    <SPLIT distance="250" swimtime="00:04:08.88" />
                    <SPLIT distance="300" swimtime="00:05:04.27" />
                    <SPLIT distance="350" swimtime="00:05:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="282" reactiontime="+92" swimtime="00:01:23.18" resultid="7351" heatid="9126" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="7253">
              <RESULTS>
                <RESULT eventid="1062" points="285" reactiontime="+95" swimtime="00:00:35.28" resultid="7254" heatid="8889" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1187" points="253" reactiontime="+91" swimtime="00:00:40.57" resultid="7255" heatid="8950" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1256" points="261" reactiontime="+112" swimtime="00:01:19.75" resultid="7256" heatid="8981" lane="1" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="252" reactiontime="+99" swimtime="00:00:38.57" resultid="7257" heatid="9056" lane="4" entrytime="00:00:37.50" />
                <RESULT eventid="1457" points="208" reactiontime="+100" swimtime="00:01:32.86" resultid="7258" heatid="9076" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="201" reactiontime="+98" swimtime="00:03:23.34" resultid="7259" heatid="9139" lane="6" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.33" />
                    <SPLIT distance="100" swimtime="00:01:42.45" />
                    <SPLIT distance="150" swimtime="00:02:35.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-12-07" firstname="Jarosław" gender="M" lastname="Zadrożny" nation="POL" athleteid="7352">
              <RESULTS>
                <RESULT eventid="1079" points="213" reactiontime="+81" swimtime="00:00:33.92" resultid="7353" heatid="8900" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1165" points="207" reactiontime="+94" swimtime="00:23:55.01" resultid="7354" heatid="8943" lane="6" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:23.75" />
                    <SPLIT distance="150" swimtime="00:02:08.87" />
                    <SPLIT distance="200" swimtime="00:02:54.93" />
                    <SPLIT distance="250" swimtime="00:03:41.31" />
                    <SPLIT distance="300" swimtime="00:04:27.69" />
                    <SPLIT distance="350" swimtime="00:05:14.76" />
                    <SPLIT distance="400" swimtime="00:06:03.00" />
                    <SPLIT distance="450" swimtime="00:06:51.26" />
                    <SPLIT distance="500" swimtime="00:07:39.50" />
                    <SPLIT distance="550" swimtime="00:08:28.38" />
                    <SPLIT distance="600" swimtime="00:09:17.04" />
                    <SPLIT distance="650" swimtime="00:10:05.14" />
                    <SPLIT distance="700" swimtime="00:10:54.32" />
                    <SPLIT distance="750" swimtime="00:11:43.15" />
                    <SPLIT distance="800" swimtime="00:12:32.70" />
                    <SPLIT distance="850" swimtime="00:13:21.96" />
                    <SPLIT distance="900" swimtime="00:14:10.69" />
                    <SPLIT distance="950" swimtime="00:14:59.76" />
                    <SPLIT distance="1000" swimtime="00:15:48.40" />
                    <SPLIT distance="1050" swimtime="00:16:38.42" />
                    <SPLIT distance="1100" swimtime="00:17:28.19" />
                    <SPLIT distance="1150" swimtime="00:18:17.54" />
                    <SPLIT distance="1200" swimtime="00:19:06.53" />
                    <SPLIT distance="1250" swimtime="00:19:56.45" />
                    <SPLIT distance="1300" swimtime="00:20:45.05" />
                    <SPLIT distance="1350" swimtime="00:21:33.99" />
                    <SPLIT distance="1400" swimtime="00:22:22.85" />
                    <SPLIT distance="1450" swimtime="00:23:11.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-02" firstname="Wojciech" gender="M" lastname="Kaczmarczyk" nation="POL" athleteid="7370">
              <RESULTS>
                <RESULT eventid="1273" points="47" reactiontime="+108" swimtime="00:02:03.75" resultid="7371" heatid="8985" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="7372" heatid="9043" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-12-18" firstname="Szymon" gender="M" lastname="Pyrć" nation="POL" athleteid="7316">
              <RESULTS>
                <RESULT eventid="1165" points="398" reactiontime="+98" swimtime="00:19:15.39" resultid="7317" heatid="8945" lane="7" entrytime="00:21:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:12.33" />
                    <SPLIT distance="150" swimtime="00:01:50.69" />
                    <SPLIT distance="200" swimtime="00:02:29.19" />
                    <SPLIT distance="250" swimtime="00:03:07.63" />
                    <SPLIT distance="300" swimtime="00:03:46.27" />
                    <SPLIT distance="350" swimtime="00:04:25.08" />
                    <SPLIT distance="400" swimtime="00:05:03.83" />
                    <SPLIT distance="450" swimtime="00:05:42.40" />
                    <SPLIT distance="500" swimtime="00:06:20.99" />
                    <SPLIT distance="550" swimtime="00:07:38.06" />
                    <SPLIT distance="600" swimtime="00:08:16.84" />
                    <SPLIT distance="650" swimtime="00:08:55.53" />
                    <SPLIT distance="700" swimtime="00:09:34.01" />
                    <SPLIT distance="800" swimtime="00:12:08.84" />
                    <SPLIT distance="850" swimtime="00:12:47.74" />
                    <SPLIT distance="900" swimtime="00:13:27.02" />
                    <SPLIT distance="950" swimtime="00:14:06.19" />
                    <SPLIT distance="1050" swimtime="00:15:24.20" />
                    <SPLIT distance="1100" swimtime="00:16:03.11" />
                    <SPLIT distance="1300" swimtime="00:18:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="368" reactiontime="+88" swimtime="00:02:31.47" resultid="7318" heatid="9029" lane="3" entrytime="00:02:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:12.76" />
                    <SPLIT distance="150" swimtime="00:01:53.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="334" reactiontime="+85" swimtime="00:05:39.31" resultid="7319" heatid="9120" lane="7" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:13.26" />
                    <SPLIT distance="200" swimtime="00:02:43.99" />
                    <SPLIT distance="250" swimtime="00:03:34.61" />
                    <SPLIT distance="300" swimtime="00:04:24.29" />
                    <SPLIT distance="350" swimtime="00:05:02.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="7333">
              <RESULTS>
                <RESULT eventid="1079" points="102" reactiontime="+71" swimtime="00:00:43.26" resultid="7334" heatid="8896" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1165" points="104" reactiontime="+114" swimtime="00:30:03.07" resultid="7335" heatid="8941" lane="7" entrytime="00:32:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:30:03.07" />
                    <SPLIT distance="100" swimtime="00:01:56.15" />
                    <SPLIT distance="150" swimtime="00:02:57.70" />
                    <SPLIT distance="200" swimtime="00:03:59.22" />
                    <SPLIT distance="250" swimtime="00:05:01.06" />
                    <SPLIT distance="300" swimtime="00:06:02.50" />
                    <SPLIT distance="350" swimtime="00:07:03.99" />
                    <SPLIT distance="400" swimtime="00:08:04.66" />
                    <SPLIT distance="450" swimtime="00:09:05.40" />
                    <SPLIT distance="500" swimtime="00:10:05.17" />
                    <SPLIT distance="550" swimtime="00:11:05.39" />
                    <SPLIT distance="600" swimtime="00:12:05.47" />
                    <SPLIT distance="650" swimtime="00:13:05.17" />
                    <SPLIT distance="700" swimtime="00:14:05.30" />
                    <SPLIT distance="750" swimtime="00:15:05.79" />
                    <SPLIT distance="800" swimtime="00:16:05.85" />
                    <SPLIT distance="850" swimtime="00:17:05.43" />
                    <SPLIT distance="900" swimtime="00:18:04.55" />
                    <SPLIT distance="950" swimtime="00:19:03.81" />
                    <SPLIT distance="1000" swimtime="00:20:03.65" />
                    <SPLIT distance="1050" swimtime="00:21:02.89" />
                    <SPLIT distance="1100" swimtime="00:22:02.34" />
                    <SPLIT distance="1150" swimtime="00:23:02.46" />
                    <SPLIT distance="1200" swimtime="00:24:02.81" />
                    <SPLIT distance="1250" swimtime="00:25:03.10" />
                    <SPLIT distance="1300" swimtime="00:26:03.61" />
                    <SPLIT distance="1350" swimtime="00:27:03.33" />
                    <SPLIT distance="1400" swimtime="00:28:03.90" />
                    <SPLIT distance="1450" swimtime="00:29:04.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="91" reactiontime="+94" swimtime="00:01:39.73" resultid="7336" heatid="8986" lane="5" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="79" reactiontime="+101" swimtime="00:03:50.67" resultid="7337" heatid="9095" lane="2" entrytime="00:03:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.99" />
                    <SPLIT distance="100" swimtime="00:01:48.67" />
                    <SPLIT distance="150" swimtime="00:02:50.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="65" reactiontime="+112" swimtime="00:01:02.61" resultid="7338" heatid="9159" lane="3" />
                <RESULT eventid="1744" points="82" reactiontime="+115" swimtime="00:08:08.30" resultid="7339" heatid="9182" lane="3" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.81" />
                    <SPLIT distance="100" swimtime="00:01:53.43" />
                    <SPLIT distance="150" swimtime="00:02:55.87" />
                    <SPLIT distance="200" swimtime="00:03:59.11" />
                    <SPLIT distance="250" swimtime="00:05:02.01" />
                    <SPLIT distance="300" swimtime="00:06:05.02" />
                    <SPLIT distance="350" swimtime="00:07:07.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Piotr" gender="M" lastname="Frankiewicz" nation="POL" athleteid="7364">
              <RESULTS>
                <RESULT eventid="1239" points="468" reactiontime="+79" swimtime="00:02:35.07" resultid="7365" heatid="8978" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:53.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="496" reactiontime="+82" swimtime="00:01:03.96" resultid="7366" heatid="9020" lane="7" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="528" reactiontime="+81" swimtime="00:01:08.80" resultid="7367" heatid="9053" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="478" reactiontime="+74" swimtime="00:00:27.87" resultid="7368" heatid="9071" lane="3" entrytime="00:00:27.80" />
                <RESULT eventid="1681" points="552" reactiontime="+74" swimtime="00:00:30.78" resultid="7369" heatid="9172" lane="7" entrytime="00:00:31.42" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="7288">
              <RESULTS>
                <RESULT eventid="1062" points="53" reactiontime="+109" swimtime="00:01:01.56" resultid="7289" heatid="8886" lane="1" entrytime="00:00:58.00" />
                <RESULT eventid="1096" points="39" reactiontime="+105" swimtime="00:05:58.10" resultid="7290" heatid="8916" lane="3" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.75" />
                    <SPLIT distance="100" swimtime="00:02:59.30" />
                    <SPLIT distance="150" swimtime="00:04:39.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="59" reactiontime="+114" swimtime="00:05:44.93" resultid="7291" heatid="8967" lane="8" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.10" />
                    <SPLIT distance="100" swimtime="00:02:41.28" />
                    <SPLIT distance="150" swimtime="00:04:12.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="46" reactiontime="+111" swimtime="00:02:37.81" resultid="7292" heatid="9001" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="70" reactiontime="+112" swimtime="00:02:31.19" resultid="7293" heatid="9037" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="28" reactiontime="+119" swimtime="00:01:19.62" resultid="7294" heatid="9054" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1595" points="27" reactiontime="+107" swimtime="00:03:01.54" resultid="7295" heatid="9123" lane="4" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="74" reactiontime="+105" swimtime="00:01:08.34" resultid="7296" heatid="9152" lane="6" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="7302">
              <RESULTS>
                <RESULT eventid="1079" points="301" reactiontime="+97" swimtime="00:00:30.21" resultid="7303" heatid="8904" lane="2" entrytime="00:00:30.10" />
                <RESULT eventid="1205" points="242" reactiontime="+85" swimtime="00:00:35.62" resultid="7304" heatid="8959" lane="0" entrytime="00:00:37.50" />
                <RESULT eventid="1307" points="298" reactiontime="+90" swimtime="00:01:15.78" resultid="7305" heatid="9014" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="327" reactiontime="+93" swimtime="00:00:31.62" resultid="7306" heatid="9066" lane="5" entrytime="00:00:32.40" />
                <RESULT eventid="1474" points="235" reactiontime="+91" swimtime="00:01:19.21" resultid="7307" heatid="9082" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="263" reactiontime="+98" swimtime="00:01:15.55" resultid="7308" heatid="9133" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="300" reactiontime="+101" swimtime="00:00:37.71" resultid="7309" heatid="9166" lane="6" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-24" firstname="Bogusław" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="7386">
              <RESULTS>
                <RESULT eventid="1079" points="45" reactiontime="+110" swimtime="00:00:56.66" resultid="7387" heatid="8895" lane="5" entrytime="00:00:57.00" />
                <RESULT eventid="1205" points="34" swimtime="00:01:08.20" resultid="7388" heatid="8955" lane="8" entrytime="00:01:07.00" />
                <RESULT eventid="1273" points="41" reactiontime="+120" swimtime="00:02:09.79" resultid="7389" heatid="8986" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="37" reactiontime="+110" swimtime="00:02:45.50" resultid="7390" heatid="9043" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="34" reactiontime="+106" swimtime="00:02:29.84" resultid="7391" heatid="9079" lane="6" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="39" reactiontime="+59" swimtime="00:05:11.10" resultid="7392" heatid="9144" lane="9" entrytime="00:05:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.41" />
                    <SPLIT distance="100" swimtime="00:02:31.02" />
                    <SPLIT distance="150" swimtime="00:03:52.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-17" firstname="Wojciech" gender="M" lastname="Liszkowski" nation="POL" athleteid="7267">
              <RESULTS>
                <RESULT eventid="1440" points="396" reactiontime="+92" swimtime="00:00:29.68" resultid="7268" heatid="9068" lane="7" entrytime="00:00:30.50" />
                <RESULT eventid="1613" points="341" reactiontime="+88" swimtime="00:01:09.33" resultid="7269" heatid="9134" lane="6" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-06" firstname="Matteo" gender="M" lastname="Morlupi" nation="POL" athleteid="7297">
              <RESULTS>
                <RESULT eventid="1079" points="268" reactiontime="+90" swimtime="00:00:31.42" resultid="7298" heatid="8903" lane="5" entrytime="00:00:30.75" />
                <RESULT eventid="1273" points="234" reactiontime="+92" swimtime="00:01:12.83" resultid="7299" heatid="8989" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="253" reactiontime="+96" swimtime="00:01:27.81" resultid="7300" heatid="9048" lane="7" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="281" reactiontime="+94" swimtime="00:00:38.54" resultid="7301" heatid="9167" lane="3" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="7279">
              <RESULTS>
                <RESULT eventid="1079" points="216" reactiontime="+105" swimtime="00:00:33.74" resultid="7280" heatid="8901" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1113" points="112" reactiontime="+119" swimtime="00:03:47.14" resultid="7281" heatid="8923" lane="2" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.86" />
                    <SPLIT distance="100" swimtime="00:01:54.40" />
                    <SPLIT distance="150" swimtime="00:03:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="206" reactiontime="+120" swimtime="00:01:15.99" resultid="7282" heatid="8990" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" reactiontime="+138" status="DNF" swimtime="00:04:41.84" resultid="7283" heatid="9026" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.96" />
                    <SPLIT distance="100" swimtime="00:01:57.82" />
                    <SPLIT distance="150" swimtime="00:03:13.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="119" reactiontime="+129" swimtime="00:00:44.30" resultid="7284" heatid="9062" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1508" points="155" reactiontime="+132" swimtime="00:03:04.92" resultid="7285" heatid="9098" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                    <SPLIT distance="100" swimtime="00:01:30.05" />
                    <SPLIT distance="150" swimtime="00:02:17.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="87" reactiontime="+131" swimtime="00:01:49.15" resultid="7286" heatid="9130" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="129" reactiontime="+124" swimtime="00:06:59.43" resultid="7287" heatid="9185" lane="1" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                    <SPLIT distance="100" swimtime="00:01:36.22" />
                    <SPLIT distance="150" swimtime="00:02:28.69" />
                    <SPLIT distance="200" swimtime="00:03:21.69" />
                    <SPLIT distance="250" swimtime="00:04:16.06" />
                    <SPLIT distance="300" swimtime="00:05:11.68" />
                    <SPLIT distance="350" swimtime="00:06:06.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-08" firstname="Tomasz" gender="M" lastname="Czerniecki" nation="POL" athleteid="7236">
              <RESULTS>
                <RESULT eventid="1079" points="517" reactiontime="+75" swimtime="00:00:25.24" resultid="7237" heatid="8913" lane="5" entrytime="00:00:26.00" />
                <RESULT eventid="1205" points="328" reactiontime="+73" swimtime="00:00:32.19" resultid="7238" heatid="8960" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="7239" heatid="8997" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1307" points="412" reactiontime="+78" swimtime="00:01:08.04" resultid="7240" heatid="9016" lane="0" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="408" reactiontime="+76" swimtime="00:00:29.37" resultid="7241" heatid="9069" lane="9" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-30" firstname="Piotr" gender="M" lastname="Łysiak" nation="POL" athleteid="7373">
              <RESULTS>
                <RESULT eventid="1307" points="290" reactiontime="+89" swimtime="00:01:16.46" resultid="7374" heatid="9015" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="317" reactiontime="+99" swimtime="00:01:21.52" resultid="7375" heatid="9050" lane="5" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="312" reactiontime="+89" swimtime="00:00:37.20" resultid="7376" heatid="9167" lane="5" entrytime="00:00:37.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-26" firstname="Józef" gender="M" lastname="Śmigielski" nation="POL" athleteid="7320">
              <RESULTS>
                <RESULT eventid="1205" points="50" reactiontime="+106" swimtime="00:01:00.08" resultid="7321" heatid="8955" lane="7" entrytime="00:00:59.90" />
                <RESULT eventid="1474" points="61" reactiontime="+106" swimtime="00:02:04.08" resultid="7322" heatid="9080" lane="8" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="58" reactiontime="+107" swimtime="00:04:32.88" resultid="7323" heatid="9144" lane="2" entrytime="00:04:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.81" />
                    <SPLIT distance="100" swimtime="00:02:12.65" />
                    <SPLIT distance="150" swimtime="00:03:24.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Masters Korona C" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="403" reactiontime="+83" swimtime="00:01:51.78" resultid="7401" heatid="9109" lane="4" entrytime="00:02:15.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="100" swimtime="00:00:58.08" />
                    <SPLIT distance="150" swimtime="00:01:26.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7267" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="7316" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="7373" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="7236" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="357" reactiontime="+91" swimtime="00:02:07.50" resultid="7402" heatid="9034" lane="2" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                    <SPLIT distance="100" swimtime="00:01:10.39" />
                    <SPLIT distance="150" swimtime="00:01:42.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7267" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="7373" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="7316" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="7236" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Masters Korona B" number="2">
              <RESULTS>
                <RESULT eventid="1548" points="363" reactiontime="+90" swimtime="00:01:55.73" resultid="7403" heatid="9111" lane="3" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:00.87" />
                    <SPLIT distance="150" swimtime="00:01:30.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7380" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="7297" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="7247" number="3" />
                    <RELAYPOSITION athleteid="7364" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="355" reactiontime="+68" swimtime="00:02:07.79" resultid="7404" heatid="9034" lane="5" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:05.61" />
                    <SPLIT distance="150" swimtime="00:01:36.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7247" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="7364" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="7380" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="7297" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Masters Korona E" number="3">
              <RESULTS>
                <RESULT eventid="1381" points="160" reactiontime="+85" swimtime="00:02:46.41" resultid="7405" heatid="9033" lane="8" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.57" />
                    <SPLIT distance="100" swimtime="00:01:30.36" />
                    <SPLIT distance="150" swimtime="00:02:01.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7279" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="7310" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="7302" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="7333" number="4" reactiontime="+77" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" name="Masters Korona F" number="3">
              <RESULTS>
                <RESULT eventid="1548" points="88" swimtime="00:03:05.70" resultid="7406" heatid="9109" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.10" />
                    <SPLIT distance="100" swimtime="00:01:44.54" />
                    <SPLIT distance="150" swimtime="00:02:31.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7320" number="1" />
                    <RELAYPOSITION athleteid="7333" number="2" reactiontime="+82" />
                    <RELAYPOSITION athleteid="7260" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="7279" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Masters Korona D" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1525" points="397" reactiontime="+84" swimtime="00:02:08.21" resultid="7399" heatid="9108" lane="3" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                    <SPLIT distance="100" swimtime="00:01:03.31" />
                    <SPLIT distance="150" swimtime="00:01:32.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7242" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="7270" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="7229" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="7360" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Masters KoronaD" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1358" points="386" reactiontime="+66" swimtime="00:02:22.82" resultid="7400" heatid="9031" lane="6" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:16.04" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7229" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="7360" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="7242" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="7270" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Masters Korona C" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1130" points="402" reactiontime="+76" swimtime="00:01:51.87" resultid="7393" heatid="8935" lane="6" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                    <SPLIT distance="100" swimtime="00:00:57.94" />
                    <SPLIT distance="150" swimtime="00:01:27.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7229" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="7380" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="7242" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="7236" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="390" reactiontime="+67" swimtime="00:02:03.81" resultid="7394" heatid="9176" lane="2" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:05.59" />
                    <SPLIT distance="150" swimtime="00:01:34.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7229" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="7364" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="7267" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="7242" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Masters Korona D" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="260" reactiontime="+90" swimtime="00:02:09.41" resultid="7395" heatid="8934" lane="7" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                    <SPLIT distance="150" swimtime="00:01:39.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7302" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="7360" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="7346" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="7316" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="253" reactiontime="+76" swimtime="00:02:23.10" resultid="7396" heatid="9175" lane="7" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:16.63" />
                    <SPLIT distance="150" swimtime="00:01:53.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7302" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="7360" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="7346" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="7373" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Masters Korona E" number="3">
              <RESULTS>
                <RESULT eventid="1130" points="183" reactiontime="+97" swimtime="00:02:25.30" resultid="7397" heatid="8933" lane="2" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:17.89" />
                    <SPLIT distance="150" swimtime="00:01:41.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7253" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="7333" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="7270" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="7279" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="138" reactiontime="+90" swimtime="00:02:55.06" resultid="7398" heatid="9174" lane="8" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:42.89" />
                    <SPLIT distance="150" swimtime="00:02:20.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7253" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="7333" number="2" reactiontime="+98" />
                    <RELAYPOSITION athleteid="7270" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="7279" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MASKRAS" nation="POL" region="LU" clubid="2556" name="Masters Kraśnik">
          <CONTACT city="Kraśnik" email="jurek@krasnik.info" internet="www.masterskrasnik.za.pl" name="Michalczyk Jerzy" phone="601 69 89 77" street="Żwirki i Wigury 2" zip="23-210" />
          <ATHLETES>
            <ATHLETE birthdate="1960-09-07" firstname="Andrzej" gender="M" lastname="Cis" nation="POL" athleteid="2562">
              <RESULTS>
                <RESULT eventid="1079" points="272" reactiontime="+74" swimtime="00:00:31.24" resultid="2563" heatid="8899" lane="7" entrytime="00:00:35.80" />
                <RESULT eventid="1205" points="188" reactiontime="+56" swimtime="00:00:38.73" resultid="2564" heatid="8958" lane="5" entrytime="00:00:38.60" />
                <RESULT eventid="1273" points="252" reactiontime="+75" swimtime="00:01:11.10" resultid="2565" heatid="8989" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="169" reactiontime="+63" swimtime="00:01:28.35" resultid="2566" heatid="9082" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="142" reactiontime="+77" swimtime="00:03:23.00" resultid="2567" heatid="9146" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.06" />
                    <SPLIT distance="100" swimtime="00:01:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2568" heatid="9184" lane="5" entrytime="00:06:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-27" firstname="Janusz" gender="M" lastname="Wasiuk" nation="POL" athleteid="2588">
              <RESULTS>
                <RESULT eventid="1165" points="90" reactiontime="+155" swimtime="00:31:33.13" resultid="2589" heatid="8940" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.78" />
                    <SPLIT distance="100" swimtime="00:02:00.11" />
                    <SPLIT distance="150" swimtime="00:03:04.68" />
                    <SPLIT distance="200" swimtime="00:04:09.61" />
                    <SPLIT distance="250" swimtime="00:05:16.44" />
                    <SPLIT distance="300" swimtime="00:06:20.32" />
                    <SPLIT distance="350" swimtime="00:07:24.89" />
                    <SPLIT distance="400" swimtime="00:08:30.54" />
                    <SPLIT distance="450" swimtime="00:09:34.97" />
                    <SPLIT distance="500" swimtime="00:10:40.78" />
                    <SPLIT distance="550" swimtime="00:11:48.09" />
                    <SPLIT distance="600" swimtime="00:12:54.42" />
                    <SPLIT distance="650" swimtime="00:13:59.76" />
                    <SPLIT distance="700" swimtime="00:15:05.94" />
                    <SPLIT distance="750" swimtime="00:16:10.17" />
                    <SPLIT distance="800" swimtime="00:17:14.36" />
                    <SPLIT distance="850" swimtime="00:18:16.38" />
                    <SPLIT distance="900" swimtime="00:19:20.75" />
                    <SPLIT distance="950" swimtime="00:20:22.05" />
                    <SPLIT distance="1000" swimtime="00:21:25.33" />
                    <SPLIT distance="1050" swimtime="00:22:26.86" />
                    <SPLIT distance="1100" swimtime="00:23:27.66" />
                    <SPLIT distance="1150" swimtime="00:24:28.80" />
                    <SPLIT distance="1200" swimtime="00:25:29.40" />
                    <SPLIT distance="1250" swimtime="00:26:31.57" />
                    <SPLIT distance="1300" swimtime="00:27:35.57" />
                    <SPLIT distance="1350" swimtime="00:28:37.75" />
                    <SPLIT distance="1400" swimtime="00:29:38.89" />
                    <SPLIT distance="1450" swimtime="00:30:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="98" reactiontime="+97" swimtime="00:00:48.15" resultid="2590" heatid="8955" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1239" points="152" reactiontime="+109" swimtime="00:03:45.31" resultid="2591" heatid="8972" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                    <SPLIT distance="100" swimtime="00:01:47.91" />
                    <SPLIT distance="150" swimtime="00:02:47.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="160" reactiontime="+112" swimtime="00:01:42.33" resultid="2592" heatid="9045" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="91" reactiontime="+144" swimtime="00:08:42.45" resultid="2593" heatid="9117" lane="9" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.12" />
                    <SPLIT distance="100" swimtime="00:02:07.61" />
                    <SPLIT distance="150" swimtime="00:03:19.73" />
                    <SPLIT distance="200" swimtime="00:04:29.80" />
                    <SPLIT distance="250" swimtime="00:05:38.62" />
                    <SPLIT distance="300" swimtime="00:06:45.73" />
                    <SPLIT distance="350" swimtime="00:07:45.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="112" reactiontime="+122" swimtime="00:01:40.31" resultid="2594" heatid="9128" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="192" reactiontime="+107" swimtime="00:00:43.71" resultid="2595" heatid="9161" lane="7" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-12-19" firstname="Waldemar" gender="M" lastname="Rusowicz" nation="POL" athleteid="2575">
              <RESULTS>
                <RESULT eventid="1113" points="120" reactiontime="+99" swimtime="00:03:42.17" resultid="2576" heatid="8922" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.84" />
                    <SPLIT distance="100" swimtime="00:01:52.66" />
                    <SPLIT distance="150" swimtime="00:02:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="178" reactiontime="+103" swimtime="00:03:34.00" resultid="2577" heatid="8973" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.17" />
                    <SPLIT distance="100" swimtime="00:01:43.82" />
                    <SPLIT distance="150" swimtime="00:02:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="127" reactiontime="+101" swimtime="00:01:40.60" resultid="2578" heatid="9009" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="171" reactiontime="+98" swimtime="00:01:40.03" resultid="2579" heatid="9045" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="2580" heatid="9060" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1474" points="69" reactiontime="+96" swimtime="00:01:58.82" resultid="2581" heatid="9080" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="168" reactiontime="+109" swimtime="00:00:45.76" resultid="2582" heatid="9162" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="2569">
              <RESULTS>
                <RESULT eventid="1079" points="109" reactiontime="+102" swimtime="00:00:42.39" resultid="2570" heatid="8898" lane="0" entrytime="00:00:38.40" />
                <RESULT eventid="1307" points="110" reactiontime="+96" swimtime="00:01:45.73" resultid="2571" heatid="9009" lane="7" entrytime="00:01:55.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K5 - Brak wynurzenia części głowy w czasie każdego pełnego cykluruchu (ramion i nóg), za wyjątkim pierwszego cyklu postarciei nawrocie (Time: 16:29)" eventid="1406" reactiontime="+101" status="DSQ" swimtime="00:01:55.56" resultid="2572" heatid="9044" lane="3" entrytime="00:01:54.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="92" reactiontime="+93" swimtime="00:00:48.14" resultid="2573" heatid="9061" lane="9" entrytime="00:00:49.20" />
                <RESULT eventid="1681" points="117" reactiontime="+96" swimtime="00:00:51.58" resultid="2574" heatid="9161" lane="8" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="2583">
              <RESULTS>
                <RESULT eventid="1113" points="118" reactiontime="+109" swimtime="00:03:43.16" resultid="2584" heatid="8922" lane="1" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.95" />
                    <SPLIT distance="100" swimtime="00:01:44.86" />
                    <SPLIT distance="150" swimtime="00:02:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="75" reactiontime="+99" swimtime="00:04:16.66" resultid="2585" heatid="9025" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.69" />
                    <SPLIT distance="100" swimtime="00:01:59.46" />
                    <SPLIT distance="150" swimtime="00:03:08.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="113" reactiontime="+93" swimtime="00:08:06.70" resultid="2586" heatid="9117" lane="3" entrytime="00:07:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.26" />
                    <SPLIT distance="100" swimtime="00:01:57.42" />
                    <SPLIT distance="150" swimtime="00:03:00.16" />
                    <SPLIT distance="200" swimtime="00:04:00.58" />
                    <SPLIT distance="250" swimtime="00:05:10.67" />
                    <SPLIT distance="300" swimtime="00:06:20.21" />
                    <SPLIT distance="350" swimtime="00:07:14.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="107" reactiontime="+89" swimtime="00:03:43.50" resultid="2587" heatid="9144" lane="4" entrytime="00:03:54.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.81" />
                    <SPLIT distance="100" swimtime="00:01:48.36" />
                    <SPLIT distance="150" swimtime="00:02:46.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" nation="POL" clubid="2754" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Tomasz Doniec" phone="693703490" />
          <ATHLETES>
            <ATHLETE birthdate="1973-11-06" firstname="Małgorzata" gender="F" lastname="Wach" nation="POL" athleteid="2774">
              <RESULTS>
                <RESULT eventid="1187" points="272" reactiontime="+60" swimtime="00:00:39.60" resultid="2775" heatid="8951" lane="9" entrytime="00:00:39.50" entrycourse="SCM" />
                <RESULT eventid="1256" points="255" reactiontime="+87" swimtime="00:01:20.42" resultid="2776" heatid="8981" lane="8" entrytime="00:01:21.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="241" reactiontime="+84" swimtime="00:02:57.97" resultid="2777" heatid="9090" lane="5" entrytime="00:03:01.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:27.09" />
                    <SPLIT distance="150" swimtime="00:02:14.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="245" reactiontime="+89" swimtime="00:00:45.97" resultid="2778" heatid="9155" lane="9" entrytime="00:00:45.57" entrycourse="SCM" />
                <RESULT eventid="1062" points="286" reactiontime="+83" swimtime="00:00:35.25" resultid="3140" heatid="8888" lane="4" entrytime="00:00:37.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-02-07" firstname="Bogdan" gender="M" lastname="Szczurek" nation="POL" athleteid="2817">
              <RESULTS>
                <RESULT eventid="1079" points="76" reactiontime="+113" swimtime="00:00:47.76" resultid="2818" heatid="8896" lane="9" entrytime="00:00:49.42" entrycourse="SCM" />
                <RESULT eventid="1165" reactiontime="+131" status="OTL" swimtime="00:37:26.56" resultid="2819" heatid="8941" lane="0" entrytime="00:35:32.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.61" />
                    <SPLIT distance="100" swimtime="00:01:58.21" />
                    <SPLIT distance="150" swimtime="00:03:09.45" />
                    <SPLIT distance="200" swimtime="00:04:20.88" />
                    <SPLIT distance="250" swimtime="00:05:33.94" />
                    <SPLIT distance="300" swimtime="00:07:59.39" />
                    <SPLIT distance="350" swimtime="00:09:13.22" />
                    <SPLIT distance="400" swimtime="00:10:28.75" />
                    <SPLIT distance="450" swimtime="00:11:41.28" />
                    <SPLIT distance="500" swimtime="00:12:58.06" />
                    <SPLIT distance="550" swimtime="00:14:18.66" />
                    <SPLIT distance="600" swimtime="00:15:39.97" />
                    <SPLIT distance="650" swimtime="00:16:48.65" />
                    <SPLIT distance="700" swimtime="00:18:06.25" />
                    <SPLIT distance="750" swimtime="00:19:26.86" />
                    <SPLIT distance="800" swimtime="00:20:42.25" />
                    <SPLIT distance="850" swimtime="00:21:58.67" />
                    <SPLIT distance="900" swimtime="00:23:08.30" />
                    <SPLIT distance="950" swimtime="00:24:25.39" />
                    <SPLIT distance="1000" swimtime="00:25:44.38" />
                    <SPLIT distance="1050" swimtime="00:27:02.01" />
                    <SPLIT distance="1100" swimtime="00:30:53.43" />
                    <SPLIT distance="1150" swimtime="00:32:16.71" />
                    <SPLIT distance="1200" swimtime="00:33:33.30" />
                    <SPLIT distance="1250" swimtime="00:34:52.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="55" reactiontime="+106" swimtime="00:00:58.39" resultid="2820" heatid="8954" lane="2" />
                <RESULT eventid="1273" points="56" reactiontime="+127" swimtime="00:01:56.96" resultid="2821" heatid="8986" lane="6" entrytime="00:01:55.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="59" reactiontime="+92" swimtime="00:02:05.30" resultid="2822" heatid="9080" lane="9" entrytime="00:02:07.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="2823" heatid="9095" lane="8" entrytime="00:04:16.09" entrycourse="SCM" />
                <RESULT eventid="1647" points="58" reactiontime="+88" swimtime="00:04:32.67" resultid="2824" heatid="9143" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.29" />
                    <SPLIT distance="100" swimtime="00:02:13.13" />
                    <SPLIT distance="150" swimtime="00:03:23.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2825" heatid="9182" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-16" firstname="Tomasz" gender="M" lastname="Doniec" nation="POL" athleteid="2810">
              <RESULTS>
                <RESULT eventid="1079" points="209" reactiontime="+89" swimtime="00:00:34.12" resultid="2811" heatid="8901" lane="9" entrytime="00:00:32.44" entrycourse="SCM" />
                <RESULT eventid="1239" points="201" reactiontime="+98" swimtime="00:03:25.50" resultid="2812" heatid="8973" lane="4" entrytime="00:03:26.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:36.76" />
                    <SPLIT distance="150" swimtime="00:02:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="245" reactiontime="+103" swimtime="00:01:28.86" resultid="2813" heatid="9048" lane="2" entrytime="00:01:29.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="2814" heatid="9062" lane="6" entrytime="00:00:39.95" entrycourse="SCM" />
                <RESULT comment="M4 - Obrót na plecy w czasie wyścigu (za wyjątkiem wykonania nawrotu, po dotknięciu dłońmi, a przed opuszczeniem ściany) (Time: 9:22)" eventid="1613" reactiontime="+113" status="DSQ" swimtime="00:01:50.42" resultid="2815" heatid="9128" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="281" reactiontime="+94" swimtime="00:00:38.51" resultid="2816" heatid="9165" lane="3" entrytime="00:00:39.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-22" firstname="Mateusz" gender="M" lastname="Dybek" nation="POL" athleteid="2803">
              <RESULTS>
                <RESULT eventid="1079" points="468" reactiontime="+93" swimtime="00:00:26.08" resultid="2804" heatid="8912" lane="7" entrytime="00:00:26.40" entrycourse="SCM" />
                <RESULT eventid="1273" points="492" reactiontime="+82" swimtime="00:00:56.90" resultid="2805" heatid="8999" lane="4" entrytime="00:00:56.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="431" reactiontime="+83" swimtime="00:01:07.06" resultid="2806" heatid="9018" lane="7" entrytime="00:01:09.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="495" reactiontime="+78" swimtime="00:00:27.54" resultid="2807" heatid="9070" lane="5" entrytime="00:00:28.50" entrycourse="SCM" />
                <RESULT eventid="1508" points="411" reactiontime="+84" swimtime="00:02:13.58" resultid="2808" heatid="9103" lane="4" entrytime="00:02:12.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:03.73" />
                    <SPLIT distance="150" swimtime="00:01:39.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="397" reactiontime="+84" swimtime="00:01:05.89" resultid="2809" heatid="9133" lane="4" entrytime="00:01:10.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="2826">
              <RESULTS>
                <RESULT eventid="1079" points="106" reactiontime="+116" swimtime="00:00:42.71" resultid="2827" heatid="8897" lane="6" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT comment="Rekord Polski" eventid="1113" points="74" reactiontime="+118" swimtime="00:04:20.52" resultid="2828" heatid="8922" lane="8" entrytime="00:04:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.51" />
                    <SPLIT distance="100" swimtime="00:02:15.40" />
                    <SPLIT distance="150" swimtime="00:03:26.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1205" points="69" reactiontime="+85" swimtime="00:00:54.15" resultid="2829" heatid="8956" lane="9" entrytime="00:00:54.00" entrycourse="SCM" />
                <RESULT comment="Rekord Polski" eventid="1273" points="101" reactiontime="+136" swimtime="00:01:36.21" resultid="2830" heatid="8987" lane="1" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1440" points="45" reactiontime="+116" swimtime="00:01:01.08" resultid="2831" heatid="9060" lane="7" entrytime="00:01:02.00" entrycourse="SCM" />
                <RESULT comment="Rekord Polski" eventid="1508" points="97" reactiontime="+125" swimtime="00:03:35.62" resultid="2832" heatid="9095" lane="5" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                    <SPLIT distance="100" swimtime="00:01:40.97" />
                    <SPLIT distance="150" swimtime="00:02:37.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="94" reactiontime="+113" swimtime="00:00:55.45" resultid="2833" heatid="9160" lane="6" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2834" heatid="9183" lane="6" entrytime="00:07:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-04" firstname="Małgorzata" gender="F" lastname="Skalska" nation="POL" athleteid="2768">
              <RESULTS>
                <RESULT eventid="1222" points="230" reactiontime="+86" swimtime="00:03:39.44" resultid="2769" heatid="8969" lane="0" entrytime="00:03:35.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                    <SPLIT distance="100" swimtime="00:01:44.85" />
                    <SPLIT distance="150" swimtime="00:02:42.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="194" reactiontime="+87" swimtime="00:01:37.87" resultid="2770" heatid="9003" lane="1" entrytime="00:01:39.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="232" reactiontime="+82" swimtime="00:01:41.41" resultid="2771" heatid="9040" lane="0" entrytime="00:01:38.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="179" reactiontime="+81" swimtime="00:03:16.56" resultid="2772" heatid="9090" lane="8" entrytime="00:03:20.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                    <SPLIT distance="100" swimtime="00:01:35.87" />
                    <SPLIT distance="150" swimtime="00:02:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="226" reactiontime="+76" swimtime="00:00:47.28" resultid="2773" heatid="9154" lane="5" entrytime="00:00:46.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="2861">
              <RESULTS>
                <RESULT eventid="1222" points="91" reactiontime="+117" swimtime="00:04:59.17" resultid="2862" heatid="8967" lane="2" entrytime="00:04:30.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.48" />
                    <SPLIT distance="100" swimtime="00:02:20.10" />
                    <SPLIT distance="150" swimtime="00:03:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="79" reactiontime="+77" swimtime="00:02:07.72" resultid="2863" heatid="9075" lane="9" entrytime="00:02:02.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="80" reactiontime="+91" swimtime="00:04:35.63" resultid="2864" heatid="9139" lane="9" entrytime="00:04:16.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.69" />
                    <SPLIT distance="100" swimtime="00:02:09.73" />
                    <SPLIT distance="150" swimtime="00:03:22.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-25" firstname="Jerzy" gender="M" lastname="Korba" nation="POL" athleteid="2794">
              <RESULTS>
                <RESULT eventid="1079" points="400" reactiontime="+77" swimtime="00:00:27.49" resultid="2795" heatid="8909" lane="3" entrytime="00:00:27.90" entrycourse="SCM" />
                <RESULT eventid="1165" points="342" reactiontime="+98" swimtime="00:20:14.76" resultid="2796" heatid="8945" lane="5" entrytime="00:21:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                    <SPLIT distance="100" swimtime="00:01:13.07" />
                    <SPLIT distance="150" swimtime="00:01:52.27" />
                    <SPLIT distance="200" swimtime="00:02:32.00" />
                    <SPLIT distance="250" swimtime="00:03:12.21" />
                    <SPLIT distance="300" swimtime="00:03:52.36" />
                    <SPLIT distance="350" swimtime="00:04:33.11" />
                    <SPLIT distance="400" swimtime="00:05:13.16" />
                    <SPLIT distance="450" swimtime="00:05:53.44" />
                    <SPLIT distance="500" swimtime="00:06:34.05" />
                    <SPLIT distance="550" swimtime="00:07:14.60" />
                    <SPLIT distance="600" swimtime="00:07:55.93" />
                    <SPLIT distance="650" swimtime="00:08:36.46" />
                    <SPLIT distance="700" swimtime="00:09:17.70" />
                    <SPLIT distance="750" swimtime="00:09:58.53" />
                    <SPLIT distance="800" swimtime="00:10:39.46" />
                    <SPLIT distance="850" swimtime="00:11:20.49" />
                    <SPLIT distance="900" swimtime="00:12:01.80" />
                    <SPLIT distance="950" swimtime="00:12:43.29" />
                    <SPLIT distance="1000" swimtime="00:13:24.31" />
                    <SPLIT distance="1050" swimtime="00:14:05.30" />
                    <SPLIT distance="1150" swimtime="00:16:09.80" />
                    <SPLIT distance="1200" swimtime="00:16:51.20" />
                    <SPLIT distance="1250" swimtime="00:17:33.38" />
                    <SPLIT distance="1300" swimtime="00:18:15.41" />
                    <SPLIT distance="1400" swimtime="00:19:38.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="324" reactiontime="+87" swimtime="00:02:55.40" resultid="2797" heatid="8976" lane="0" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:01:24.00" />
                    <SPLIT distance="150" swimtime="00:02:10.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2798" heatid="8996" lane="9" entrytime="00:01:01.50" entrycourse="SCM" />
                <RESULT eventid="1406" points="355" reactiontime="+91" swimtime="00:01:18.53" resultid="2799" heatid="9051" lane="0" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="281" reactiontime="+101" swimtime="00:05:59.15" resultid="2800" heatid="9120" lane="2" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:25.21" />
                    <SPLIT distance="150" swimtime="00:02:12.75" />
                    <SPLIT distance="200" swimtime="00:02:58.28" />
                    <SPLIT distance="250" swimtime="00:03:50.15" />
                    <SPLIT distance="300" swimtime="00:04:41.90" />
                    <SPLIT distance="350" swimtime="00:05:22.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="379" reactiontime="+81" swimtime="00:00:34.89" resultid="2801" heatid="9169" lane="7" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-28" firstname="Wojciech" gender="M" lastname="Wolski" nation="POL" athleteid="2865">
              <RESULTS>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="2866" heatid="9028" lane="7" entrytime="00:03:09.76" entrycourse="SCM" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="2867" heatid="9119" lane="9" entrytime="00:06:50.54" entrycourse="SCM" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="2868" heatid="9132" lane="0" entrytime="00:01:22.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="2779">
              <RESULTS>
                <RESULT eventid="1062" points="587" reactiontime="+88" swimtime="00:00:27.75" resultid="2780" heatid="8893" lane="7" entrytime="00:00:28.30" entrycourse="SCM" />
                <RESULT eventid="1096" points="584" reactiontime="+81" swimtime="00:02:25.71" resultid="2781" heatid="8920" lane="4" entrytime="00:02:28.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:09.83" />
                    <SPLIT distance="150" swimtime="00:01:51.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="609" reactiontime="+79" swimtime="00:01:00.17" resultid="2782" heatid="8984" lane="5" entrytime="00:00:59.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="581" reactiontime="+83" swimtime="00:01:07.92" resultid="2783" heatid="9007" lane="3" entrytime="00:01:08.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="529" reactiontime="+84" swimtime="00:01:17.10" resultid="2784" heatid="9042" lane="4" entrytime="00:01:14.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="630" reactiontime="+82" swimtime="00:02:09.17" resultid="2785" heatid="9093" lane="4" entrytime="00:02:12.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:02.23" />
                    <SPLIT distance="150" swimtime="00:01:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="490" reactiontime="+80" swimtime="00:01:09.25" resultid="2786" heatid="9127" lane="6" entrytime="00:01:09.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="577" reactiontime="+81" swimtime="00:00:34.58" resultid="2787" heatid="9158" lane="4" entrytime="00:00:34.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-03-22" firstname="Sandra" gender="F" lastname="Wolska" nation="POL" athleteid="2835">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="2836" heatid="8919" lane="9" entrytime="00:03:05.00" entrycourse="SCM" />
                <RESULT eventid="1222" points="277" reactiontime="+88" swimtime="00:03:26.22" resultid="2837" heatid="8970" lane="3" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:01:32.63" />
                    <SPLIT distance="150" swimtime="00:02:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="134" reactiontime="+92" swimtime="00:03:53.72" resultid="2838" heatid="9022" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                    <SPLIT distance="100" swimtime="00:01:44.77" />
                    <SPLIT distance="150" swimtime="00:02:47.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="307" reactiontime="+87" swimtime="00:01:32.36" resultid="2839" heatid="9036" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="223" reactiontime="+92" swimtime="00:07:08.38" resultid="2840" heatid="9113" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="100" swimtime="00:01:45.05" />
                    <SPLIT distance="150" swimtime="00:02:41.23" />
                    <SPLIT distance="200" swimtime="00:03:37.34" />
                    <SPLIT distance="250" swimtime="00:04:31.17" />
                    <SPLIT distance="300" swimtime="00:05:27.47" />
                    <SPLIT distance="350" swimtime="00:06:18.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="149" reactiontime="+96" swimtime="00:01:42.97" resultid="2841" heatid="9123" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="334" reactiontime="+87" swimtime="00:00:41.49" resultid="2842" heatid="9152" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-27" firstname="Michał" gender="M" lastname="Klupa" nation="POL" athleteid="2849">
              <RESULTS>
                <RESULT eventid="1113" points="464" reactiontime="+76" swimtime="00:02:21.55" resultid="2850" heatid="8931" lane="1" entrytime="00:02:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="100" swimtime="00:01:04.20" />
                    <SPLIT distance="150" swimtime="00:01:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="474" reactiontime="+61" swimtime="00:00:28.48" resultid="2851" heatid="8964" lane="5" entrytime="00:00:28.50" entrycourse="SCM" />
                <RESULT eventid="1307" points="505" reactiontime="+79" swimtime="00:01:03.61" resultid="2852" heatid="9020" lane="1" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="498" reactiontime="+66" swimtime="00:01:01.73" resultid="2853" heatid="9087" lane="0" entrytime="00:01:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="496" reactiontime="+77" swimtime="00:02:05.50" resultid="2854" heatid="9105" lane="7" entrytime="00:02:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                    <SPLIT distance="100" swimtime="00:00:59.91" />
                    <SPLIT distance="150" swimtime="00:01:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="460" reactiontime="+69" swimtime="00:02:17.37" resultid="2855" heatid="9150" lane="2" entrytime="00:02:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:06.72" />
                    <SPLIT distance="150" swimtime="00:01:41.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-08-12" firstname="Konrad" gender="M" lastname="Plutecki" nation="POL" athleteid="2856">
              <RESULTS>
                <RESULT eventid="1079" points="438" reactiontime="+79" swimtime="00:00:26.66" resultid="2857" heatid="8911" lane="0" entrytime="00:00:26.80" entrycourse="SCM" />
                <RESULT eventid="1273" points="470" reactiontime="+78" swimtime="00:00:57.80" resultid="2858" heatid="8998" lane="8" entrytime="00:00:59.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="465" reactiontime="+79" swimtime="00:02:08.21" resultid="2859" heatid="9102" lane="3" entrytime="00:02:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="100" swimtime="00:01:01.61" />
                    <SPLIT distance="150" swimtime="00:01:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="398" reactiontime="+75" swimtime="00:04:48.34" resultid="2860" heatid="9189" lane="5" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                    <SPLIT distance="200" swimtime="00:02:24.73" />
                    <SPLIT distance="250" swimtime="00:03:01.24" />
                    <SPLIT distance="300" swimtime="00:03:36.25" />
                    <SPLIT distance="350" swimtime="00:04:09.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-06" firstname="Sebastian" gender="M" lastname="Buzowski" nation="POL" athleteid="2843">
              <RESULTS>
                <RESULT eventid="1079" points="441" reactiontime="+80" swimtime="00:00:26.61" resultid="2844" heatid="8910" lane="2" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1205" points="299" reactiontime="+73" swimtime="00:00:33.22" resultid="2845" heatid="8961" lane="2" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="422" reactiontime="+77" swimtime="00:00:59.89" resultid="2846" heatid="8996" lane="4" entrytime="00:01:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="392" reactiontime="+85" swimtime="00:00:29.77" resultid="2847" heatid="9069" lane="1" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1508" points="308" reactiontime="+79" swimtime="00:02:27.06" resultid="2848" heatid="9101" lane="7" entrytime="00:02:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:07.00" />
                    <SPLIT distance="150" swimtime="00:01:46.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-16" firstname="Kamil" gender="M" lastname="Latuszek" nation="POL" athleteid="2788">
              <RESULTS>
                <RESULT eventid="1079" points="467" reactiontime="+76" swimtime="00:00:26.11" resultid="2789" heatid="8911" lane="3" entrytime="00:00:26.50" entrycourse="SCM" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2790" heatid="8946" lane="9" entrytime="00:21:14.99" entrycourse="SCM" />
                <RESULT eventid="1273" points="473" reactiontime="+81" swimtime="00:00:57.65" resultid="2791" heatid="8999" lane="0" entrytime="00:00:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="422" reactiontime="+79" swimtime="00:00:29.06" resultid="2792" heatid="9071" lane="0" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1508" points="384" reactiontime="+80" swimtime="00:02:16.61" resultid="2793" heatid="9103" lane="1" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                    <SPLIT distance="150" swimtime="00:01:41.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="Palmowska" nation="POL" athleteid="2760">
              <RESULTS>
                <RESULT eventid="1096" points="431" reactiontime="+70" swimtime="00:02:41.29" resultid="2761" heatid="8920" lane="3" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:02:02.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="445" reactiontime="+66" swimtime="00:00:33.60" resultid="2762" heatid="8953" lane="0" entrytime="00:00:33.50" entrycourse="SCM" />
                <RESULT eventid="1290" points="449" reactiontime="+69" swimtime="00:01:14.04" resultid="2763" heatid="9007" lane="2" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="437" reactiontime="+63" swimtime="00:01:12.49" resultid="2764" heatid="9078" lane="7" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="395" reactiontime="+74" swimtime="00:02:30.86" resultid="2765" heatid="9093" lane="0" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                    <SPLIT distance="150" swimtime="00:01:52.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="437" reactiontime="+67" swimtime="00:02:37.04" resultid="2766" heatid="9141" lane="2" entrytime="00:02:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:16.35" />
                    <SPLIT distance="150" swimtime="00:01:56.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="419" reactiontime="+65" swimtime="00:05:13.17" resultid="2767" heatid="9181" lane="7" entrytime="00:05:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:54.04" />
                    <SPLIT distance="200" swimtime="00:02:34.15" />
                    <SPLIT distance="250" swimtime="00:03:14.23" />
                    <SPLIT distance="300" swimtime="00:03:55.01" />
                    <SPLIT distance="350" swimtime="00:04:35.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="3663" heatid="8938" lane="5" entrytime="00:12:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-19" firstname="Paulina" gender="F" lastname="Palka" nation="POL" athleteid="2755">
              <RESULTS>
                <RESULT eventid="1187" points="424" reactiontime="+56" swimtime="00:00:34.16" resultid="2756" heatid="8952" lane="8" entrytime="00:00:35.60" entrycourse="SCM" />
                <RESULT eventid="1457" points="429" reactiontime="+58" swimtime="00:01:12.93" resultid="2757" heatid="9077" lane="5" entrytime="00:01:18.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="345" reactiontime="+73" swimtime="00:06:10.45" resultid="2758" heatid="9114" lane="3" entrytime="00:06:30.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:31.95" />
                    <SPLIT distance="150" swimtime="00:02:18.02" />
                    <SPLIT distance="200" swimtime="00:03:04.49" />
                    <SPLIT distance="250" swimtime="00:03:57.81" />
                    <SPLIT distance="300" swimtime="00:04:49.05" />
                    <SPLIT distance="350" swimtime="00:05:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="397" reactiontime="+57" swimtime="00:02:42.22" resultid="2759" heatid="9140" lane="7" entrytime="00:02:58.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:19.53" />
                    <SPLIT distance="150" swimtime="00:02:01.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="455" reactiontime="+67" swimtime="00:01:57.60" resultid="2873" heatid="9034" lane="1" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="100" swimtime="00:01:03.70" />
                    <SPLIT distance="150" swimtime="00:01:32.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2849" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="2794" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="2788" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2803" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="502" reactiontime="+80" swimtime="00:01:43.91" resultid="2874" heatid="9111" lane="4" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                    <SPLIT distance="100" swimtime="00:00:51.19" />
                    <SPLIT distance="150" swimtime="00:01:17.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2803" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2849" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="2788" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="2843" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT comment="G7 - Brak pozycji na plecach przy opuszczaniu ściany nawrotowej (Time: 13:25)" eventid="1381" reactiontime="+134" status="DSQ" swimtime="00:02:36.79" resultid="2875" heatid="9032" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.95" />
                    <SPLIT distance="100" swimtime="00:01:34.81" />
                    <SPLIT distance="150" swimtime="00:02:09.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2826" number="1" reactiontime="+134" status="DSQ" />
                    <RELAYPOSITION athleteid="2810" number="2" reactiontime="+40" status="DSQ" />
                    <RELAYPOSITION athleteid="2865" number="3" reactiontime="+33" status="DSQ" />
                    <RELAYPOSITION athleteid="2843" number="4" reactiontime="+58" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="215" reactiontime="+87" swimtime="00:02:17.86" resultid="2876" heatid="9109" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                    <SPLIT distance="150" swimtime="00:01:49.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2865" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="2826" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2810" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="2794" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="213" reactiontime="+73" swimtime="00:02:53.99" resultid="2871" heatid="9031" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:34.65" />
                    <SPLIT distance="150" swimtime="00:02:18.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2760" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="2861" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2768" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2774" number="4" reactiontime="+85" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="208" reactiontime="+67" swimtime="00:02:39.03" resultid="2872" heatid="9107" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:22.79" />
                    <SPLIT distance="150" swimtime="00:02:02.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2760" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="2861" number="2" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2768" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2774" number="4" reactiontime="+84" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="353" swimtime="00:01:56.81" resultid="2869" heatid="8932" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="100" swimtime="00:01:05.12" />
                    <SPLIT distance="150" swimtime="00:01:31.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2760" number="1" />
                    <RELAYPOSITION athleteid="2774" number="2" />
                    <RELAYPOSITION athleteid="2849" number="3" />
                    <RELAYPOSITION athleteid="2788" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="304" reactiontime="+61" swimtime="00:02:14.58" resultid="2870" heatid="9173" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:08.91" />
                    <SPLIT distance="150" swimtime="00:01:36.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2760" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2794" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="2849" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="2768" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1698" points="115" reactiontime="+74" swimtime="00:03:05.70" resultid="2877" heatid="9173" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.61" />
                    <SPLIT distance="100" swimtime="00:01:54.37" />
                    <SPLIT distance="150" swimtime="00:02:29.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2861" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2826" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="2865" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2774" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4892" name="Masters Zdzieszowice">
          <CONTACT name="Jajuga" />
          <ATHLETES>
            <ATHLETE birthdate="1967-01-21" firstname="Andrzej" gender="M" lastname="Rola" nation="POL" athleteid="4924">
              <RESULTS>
                <RESULT eventid="1079" points="275" reactiontime="+84" swimtime="00:00:31.15" resultid="4925" heatid="8909" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="1205" points="207" reactiontime="+72" swimtime="00:00:37.56" resultid="4926" heatid="8960" lane="8" entrytime="00:00:34.50" />
                <RESULT eventid="1307" points="262" reactiontime="+101" swimtime="00:01:19.10" resultid="4927" heatid="9014" lane="1" entrytime="00:01:17.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="4928" heatid="9083" lane="3" entrytime="00:01:15.34" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-08" firstname="Jacek" gender="M" lastname="Zalejski" nation="POL" athleteid="4920">
              <RESULTS>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="4921" heatid="8989" lane="8" entrytime="00:01:15.45" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="4922" heatid="9012" lane="8" entrytime="00:01:25.34" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="4923" heatid="9063" lane="5" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-23" firstname="Katarzyna" gender="F" lastname="Gniot" nation="POL" athleteid="4899">
              <RESULTS>
                <RESULT eventid="1062" points="173" reactiontime="+100" swimtime="00:00:41.70" resultid="4900" heatid="8888" lane="5" entrytime="00:00:37.33" />
                <RESULT eventid="1664" points="178" reactiontime="+101" swimtime="00:00:51.15" resultid="4901" heatid="9155" lane="8" entrytime="00:00:45.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Grzegorz" gender="M" lastname="Sierka" nation="POL" athleteid="4912">
              <RESULTS>
                <RESULT eventid="1205" points="460" reactiontime="+62" swimtime="00:00:28.78" resultid="4913" heatid="8964" lane="4" entrytime="00:00:28.45" />
                <RESULT eventid="1307" points="487" reactiontime="+78" swimtime="00:01:04.39" resultid="4914" heatid="9020" lane="4" entrytime="00:01:02.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="489" swimtime="00:01:02.08" resultid="4915" heatid="9087" lane="2" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="413" reactiontime="+78" swimtime="00:02:13.35" resultid="4916" heatid="9105" lane="9" entrytime="00:02:09.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:04.93" />
                    <SPLIT distance="150" swimtime="00:01:39.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-05" firstname="Szymon" gender="M" lastname="Paciej" nation="POL" athleteid="4917">
              <RESULTS>
                <RESULT eventid="1307" points="362" reactiontime="+85" swimtime="00:01:11.08" resultid="4918" heatid="9014" lane="5" entrytime="00:01:15.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="332" reactiontime="+90" swimtime="00:00:31.46" resultid="4919" heatid="9068" lane="6" entrytime="00:00:30.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="4907">
              <RESULTS>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="4908" heatid="8946" lane="8" entrytime="00:21:00.13" />
                <RESULT eventid="1341" points="373" reactiontime="+74" swimtime="00:02:30.81" resultid="4909" heatid="9030" lane="9" entrytime="00:02:40.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:50.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="388" reactiontime="+86" swimtime="00:05:22.66" resultid="4910" heatid="9121" lane="1" entrytime="00:05:40.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:56.39" />
                    <SPLIT distance="200" swimtime="00:02:38.49" />
                    <SPLIT distance="250" swimtime="00:03:24.90" />
                    <SPLIT distance="300" swimtime="00:04:11.01" />
                    <SPLIT distance="350" swimtime="00:04:48.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="408" reactiontime="+79" swimtime="00:04:46.15" resultid="4911" heatid="9191" lane="7" entrytime="00:04:45.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:09.22" />
                    <SPLIT distance="150" swimtime="00:01:45.48" />
                    <SPLIT distance="200" swimtime="00:02:21.94" />
                    <SPLIT distance="250" swimtime="00:02:58.36" />
                    <SPLIT distance="300" swimtime="00:03:34.77" />
                    <SPLIT distance="350" swimtime="00:04:11.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-18" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="4902">
              <RESULTS>
                <RESULT eventid="1096" points="309" reactiontime="+105" swimtime="00:03:00.19" resultid="4903" heatid="8919" lane="1" entrytime="00:03:03.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:24.64" />
                    <SPLIT distance="150" swimtime="00:02:17.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="302" reactiontime="+97" swimtime="00:01:24.48" resultid="4904" heatid="9005" lane="0" entrytime="00:01:23.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="287" reactiontime="+77" swimtime="00:01:23.37" resultid="4905" heatid="9076" lane="5" entrytime="00:01:23.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="291" reactiontime="+79" swimtime="00:02:59.92" resultid="4906" heatid="9140" lane="0" entrytime="00:03:03.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="100" swimtime="00:01:26.60" />
                    <SPLIT distance="150" swimtime="00:02:13.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-08" firstname="Przemysław" gender="M" lastname="Osiwała" nation="POL" athleteid="4893">
              <RESULTS>
                <RESULT eventid="1113" points="335" reactiontime="+88" swimtime="00:02:37.70" resultid="4894" heatid="8927" lane="6" entrytime="00:02:45.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:02:01.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="317" reactiontime="+88" swimtime="00:02:39.05" resultid="4895" heatid="9029" lane="6" entrytime="00:02:42.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:15.51" />
                    <SPLIT distance="150" swimtime="00:01:56.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="357" reactiontime="+81" swimtime="00:00:30.71" resultid="4896" heatid="9068" lane="3" entrytime="00:00:30.25" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="4897" heatid="9121" lane="0" entrytime="00:05:40.22" />
                <RESULT eventid="1613" points="352" reactiontime="+79" swimtime="00:01:08.55" resultid="4898" heatid="9133" lane="5" entrytime="00:01:10.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="431" reactiontime="+85" swimtime="00:01:49.31" resultid="4931" heatid="9110" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:00:55.19" />
                    <SPLIT distance="150" swimtime="00:01:23.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4917" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="4907" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4893" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4912" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="417" reactiontime="+62" swimtime="00:02:01.12" resultid="4932" heatid="9033" lane="4" entrytime="00:02:15.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                    <SPLIT distance="150" swimtime="00:01:32.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4912" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4907" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="4893" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4917" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="235" reactiontime="+96" swimtime="00:02:13.76" resultid="4929" heatid="8933" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:01:45.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4902" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="4899" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="4924" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4893" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="210" swimtime="00:02:32.23" resultid="4930" heatid="9174" lane="5" entrytime="00:02:30.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:30.92" />
                    <SPLIT distance="150" swimtime="00:02:01.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4902" number="1" />
                    <RELAYPOSITION athleteid="4899" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4893" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4924" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3685" name="Masters Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos Rafał" phone="604184311" />
          <ATHLETES>
            <ATHLETE birthdate="1979-06-12" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" athleteid="3698">
              <RESULTS>
                <RESULT eventid="1079" points="444" reactiontime="+76" swimtime="00:00:26.54" resultid="3699" heatid="8913" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1273" points="426" reactiontime="+79" swimtime="00:00:59.70" resultid="3700" heatid="8997" lane="9" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="209" reactiontime="+93" swimtime="00:01:25.33" resultid="3701" heatid="9013" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="409" reactiontime="+79" swimtime="00:00:29.35" resultid="3702" heatid="9071" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="1613" points="379" reactiontime="+74" swimtime="00:01:06.91" resultid="3703" heatid="9135" lane="8" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-08-19" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" athleteid="3704">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="3705" heatid="8905" lane="3" entrytime="00:00:29.97" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="3706" heatid="9013" lane="9" entrytime="00:01:20.14" />
                <RESULT eventid="1406" points="266" reactiontime="+82" swimtime="00:01:26.46" resultid="3707" heatid="9047" lane="9" entrytime="00:01:31.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="3708" heatid="9120" lane="4" entrytime="00:05:53.36" />
                <RESULT eventid="1681" points="415" reactiontime="+84" swimtime="00:00:33.83" resultid="3709" heatid="9165" lane="5" entrytime="00:00:39.13" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-28" firstname="Artur" gender="M" lastname="Frąckowiak" nation="POL" athleteid="3686">
              <RESULTS>
                <RESULT eventid="1079" points="429" reactiontime="+84" swimtime="00:00:26.86" resultid="3687" heatid="8908" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1165" reactiontime="+82" status="DNF" swimtime="00:00:00.00" resultid="3688" heatid="8945" lane="3" entrytime="00:21:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:01:07.90" />
                    <SPLIT distance="150" swimtime="00:01:45.06" />
                    <SPLIT distance="200" swimtime="00:02:23.44" />
                    <SPLIT distance="250" swimtime="00:03:02.01" />
                    <SPLIT distance="300" swimtime="00:03:41.20" />
                    <SPLIT distance="350" swimtime="00:04:20.74" />
                    <SPLIT distance="400" swimtime="00:05:00.42" />
                    <SPLIT distance="450" swimtime="00:05:39.93" />
                    <SPLIT distance="500" swimtime="00:06:19.45" />
                    <SPLIT distance="550" swimtime="00:06:59.28" />
                    <SPLIT distance="600" swimtime="00:07:39.25" />
                    <SPLIT distance="650" swimtime="00:08:18.98" />
                    <SPLIT distance="700" swimtime="00:08:59.39" />
                    <SPLIT distance="750" swimtime="00:09:40.34" />
                    <SPLIT distance="800" swimtime="00:10:21.02" />
                    <SPLIT distance="850" swimtime="00:11:02.09" />
                    <SPLIT distance="900" swimtime="00:11:43.49" />
                    <SPLIT distance="950" swimtime="00:12:25.45" />
                    <SPLIT distance="1000" swimtime="00:12:46.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="445" reactiontime="+86" swimtime="00:00:58.84" resultid="3689" heatid="8995" lane="7" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="416" reactiontime="+90" swimtime="00:01:07.86" resultid="3690" heatid="9018" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="404" reactiontime="+82" swimtime="00:00:29.47" resultid="3691" heatid="9067" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1508" points="420" reactiontime="+85" swimtime="00:02:12.60" resultid="3692" heatid="9102" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                    <SPLIT distance="100" swimtime="00:01:03.04" />
                    <SPLIT distance="150" swimtime="00:01:37.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="379" reactiontime="+86" swimtime="00:04:53.16" resultid="3693" heatid="9188" lane="6" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:06.74" />
                    <SPLIT distance="150" swimtime="00:01:43.01" />
                    <SPLIT distance="200" swimtime="00:02:20.72" />
                    <SPLIT distance="250" swimtime="00:02:58.87" />
                    <SPLIT distance="300" swimtime="00:03:37.71" />
                    <SPLIT distance="350" swimtime="00:04:16.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-09" firstname="Marcin" gender="M" lastname="Strąkowski" nation="POL" athleteid="3694">
              <RESULTS>
                <RESULT eventid="1079" points="355" reactiontime="+83" swimtime="00:00:28.60" resultid="3695" heatid="8907" lane="1" entrytime="00:00:28.99" />
                <RESULT eventid="1273" points="291" reactiontime="+84" swimtime="00:01:07.80" resultid="3696" heatid="8992" lane="9" entrytime="00:01:08.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="300" reactiontime="+84" swimtime="00:00:37.70" resultid="3697" heatid="9168" lane="9" entrytime="00:00:37.27" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-31" firstname="Anna" gender="F" lastname="Jakóbczyk" nation="POL" athleteid="3747">
              <RESULTS>
                <RESULT eventid="1062" points="209" reactiontime="+98" swimtime="00:00:39.14" resultid="3748" heatid="8889" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1187" points="171" reactiontime="+87" swimtime="00:00:46.23" resultid="3749" heatid="8950" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1222" points="186" reactiontime="+98" swimtime="00:03:55.41" resultid="3750" heatid="8969" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.55" />
                    <SPLIT distance="100" swimtime="00:01:52.47" />
                    <SPLIT distance="150" swimtime="00:02:54.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="187" reactiontime="+95" swimtime="00:01:48.96" resultid="3751" heatid="9039" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="3752" heatid="9076" lane="3" entrytime="00:01:25.00" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="3753" heatid="9140" lane="1" entrytime="00:03:00.00" />
                <RESULT eventid="1664" points="206" reactiontime="+97" swimtime="00:00:48.71" resultid="3754" heatid="9155" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-18" firstname="Konrad" gender="M" lastname="Hasik" nation="POL" athleteid="3716">
              <RESULTS>
                <RESULT eventid="1079" points="421" reactiontime="+84" swimtime="00:00:27.02" resultid="3717" heatid="8915" lane="8" entrytime="00:00:24.00" />
                <RESULT eventid="1113" points="377" reactiontime="+87" swimtime="00:02:31.69" resultid="3718" heatid="8928" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                    <SPLIT distance="150" swimtime="00:01:55.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="383" reactiontime="+66" swimtime="00:00:30.59" resultid="3719" heatid="8965" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1307" points="434" reactiontime="+85" swimtime="00:01:06.88" resultid="3720" heatid="9021" lane="9" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="380" reactiontime="+89" swimtime="00:01:16.77" resultid="3721" heatid="9052" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="352" reactiontime="+67" swimtime="00:01:09.25" resultid="3722" heatid="9086" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="324" reactiontime="+72" swimtime="00:02:34.40" resultid="3723" heatid="9149" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:15.30" />
                    <SPLIT distance="150" swimtime="00:01:55.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="3740">
              <RESULTS>
                <RESULT eventid="1079" points="349" reactiontime="+81" swimtime="00:00:28.75" resultid="3741" heatid="8904" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1165" points="344" reactiontime="+89" swimtime="00:20:13.10" resultid="3742" heatid="8945" lane="4" entrytime="00:21:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:14.80" />
                    <SPLIT distance="150" swimtime="00:01:54.48" />
                    <SPLIT distance="200" swimtime="00:02:34.27" />
                    <SPLIT distance="250" swimtime="00:03:14.45" />
                    <SPLIT distance="300" swimtime="00:03:54.53" />
                    <SPLIT distance="350" swimtime="00:04:34.51" />
                    <SPLIT distance="400" swimtime="00:05:15.30" />
                    <SPLIT distance="450" swimtime="00:05:55.21" />
                    <SPLIT distance="500" swimtime="00:06:35.55" />
                    <SPLIT distance="550" swimtime="00:07:15.40" />
                    <SPLIT distance="600" swimtime="00:07:55.38" />
                    <SPLIT distance="650" swimtime="00:08:35.17" />
                    <SPLIT distance="700" swimtime="00:09:15.28" />
                    <SPLIT distance="750" swimtime="00:09:55.27" />
                    <SPLIT distance="800" swimtime="00:10:35.34" />
                    <SPLIT distance="850" swimtime="00:11:16.50" />
                    <SPLIT distance="900" swimtime="00:11:56.63" />
                    <SPLIT distance="950" swimtime="00:12:36.72" />
                    <SPLIT distance="1000" swimtime="00:13:17.77" />
                    <SPLIT distance="1050" swimtime="00:13:58.35" />
                    <SPLIT distance="1100" swimtime="00:14:38.78" />
                    <SPLIT distance="1150" swimtime="00:15:19.56" />
                    <SPLIT distance="1200" swimtime="00:16:00.70" />
                    <SPLIT distance="1250" swimtime="00:16:42.59" />
                    <SPLIT distance="1300" swimtime="00:17:25.32" />
                    <SPLIT distance="1350" swimtime="00:18:08.96" />
                    <SPLIT distance="1400" swimtime="00:18:52.49" />
                    <SPLIT distance="1450" swimtime="00:19:34.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3743" heatid="8996" lane="2" entrytime="00:01:01.01" />
                <RESULT eventid="1440" points="291" reactiontime="+86" swimtime="00:00:32.88" resultid="3744" heatid="9069" lane="6" entrytime="00:00:29.99" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="3745" heatid="9104" lane="1" entrytime="00:02:10.01" />
                <RESULT eventid="1744" points="297" reactiontime="+82" swimtime="00:05:17.96" resultid="3746" heatid="9189" lane="6" entrytime="00:05:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:11.13" />
                    <SPLIT distance="150" swimtime="00:01:50.09" />
                    <SPLIT distance="200" swimtime="00:02:29.11" />
                    <SPLIT distance="250" swimtime="00:03:09.87" />
                    <SPLIT distance="300" swimtime="00:03:52.28" />
                    <SPLIT distance="350" swimtime="00:04:35.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="3728">
              <RESULTS>
                <RESULT eventid="1079" points="356" reactiontime="+91" swimtime="00:00:28.57" resultid="3729" heatid="8899" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1113" points="261" reactiontime="+94" swimtime="00:02:51.48" resultid="3730" heatid="8924" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:19.01" />
                    <SPLIT distance="150" swimtime="00:02:09.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="3731" heatid="8974" lane="3" entrytime="00:03:20.00" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="3732" heatid="9011" lane="7" entrytime="00:01:30.00" />
                <RESULT eventid="1406" points="247" reactiontime="+98" swimtime="00:01:28.52" resultid="3733" heatid="9048" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="229" reactiontime="+93" swimtime="00:00:41.27" resultid="3734" heatid="9162" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-08" firstname="Marcin" gender="M" lastname="Babuchowski" nation="POL" athleteid="3710">
              <RESULTS>
                <RESULT eventid="1079" points="573" reactiontime="+72" swimtime="00:00:24.39" resultid="3711" heatid="8915" lane="7" entrytime="00:00:24.00" />
                <RESULT comment="Rekord Polski" eventid="1273" points="614" reactiontime="+79" swimtime="00:00:52.86" resultid="3712" heatid="9000" lane="6" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.69" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1440" points="648" reactiontime="+72" swimtime="00:00:25.18" resultid="3713" heatid="9073" lane="4" entrytime="00:00:24.50" />
                <RESULT eventid="1508" points="589" reactiontime="+75" swimtime="00:01:58.51" resultid="3714" heatid="9106" lane="3" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                    <SPLIT distance="100" swimtime="00:00:58.82" />
                    <SPLIT distance="150" swimtime="00:01:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1613" points="643" reactiontime="+73" swimtime="00:00:56.12" resultid="3715" heatid="9137" lane="4" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-02" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="3755">
              <RESULTS>
                <RESULT eventid="1079" points="443" reactiontime="+91" swimtime="00:00:26.56" resultid="3756" heatid="8913" lane="0" entrytime="00:00:26.00" />
                <RESULT eventid="1273" points="392" reactiontime="+88" swimtime="00:01:01.40" resultid="3757" heatid="8995" lane="1" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="3758" heatid="9067" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1681" points="375" reactiontime="+87" swimtime="00:00:34.99" resultid="3759" heatid="9170" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-14" firstname="Jakub" gender="M" lastname="Gryczyński" nation="POL" athleteid="3724">
              <RESULTS>
                <RESULT eventid="1079" points="324" reactiontime="+85" swimtime="00:00:29.49" resultid="3725" heatid="8902" lane="5" entrytime="00:00:31.10" />
                <RESULT eventid="1406" points="260" reactiontime="+91" swimtime="00:01:27.11" resultid="3726" heatid="9047" lane="0" entrytime="00:01:31.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="286" reactiontime="+88" swimtime="00:00:38.28" resultid="3727" heatid="9166" lane="4" entrytime="00:00:38.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-14" firstname="Damian" gender="M" lastname="Karkusiński" nation="POL" athleteid="3735">
              <RESULTS>
                <RESULT eventid="1079" points="304" reactiontime="+117" swimtime="00:00:30.12" resultid="3736" heatid="8905" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1205" points="255" reactiontime="+66" swimtime="00:00:35.03" resultid="3737" heatid="8960" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="3738" heatid="9084" lane="8" entrytime="00:01:14.00" />
                <RESULT eventid="1681" points="241" reactiontime="+86" swimtime="00:00:40.53" resultid="3739" heatid="9162" lane="7" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="468" reactiontime="+65" swimtime="00:01:56.50" resultid="3760" heatid="9035" lane="7" entrytime="00:01:53.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="150" swimtime="00:01:29.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3710" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="3716" number="2" />
                    <RELAYPOSITION athleteid="3698" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3686" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="305" reactiontime="+66" swimtime="00:02:14.43" resultid="3761" heatid="9034" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:12.97" />
                    <SPLIT distance="150" swimtime="00:01:44.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3735" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3704" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="3755" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3740" number="4" reactiontime="+95" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1548" points="500" reactiontime="+103" swimtime="00:01:44.04" resultid="3762" heatid="9112" lane="4" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="100" swimtime="00:00:53.18" />
                    <SPLIT distance="150" swimtime="00:01:20.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3755" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="3698" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3716" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3710" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1548" points="299" reactiontime="+85" swimtime="00:02:03.47" resultid="3763" heatid="9112" lane="6" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                    <SPLIT distance="100" swimtime="00:01:03.28" />
                    <SPLIT distance="150" swimtime="00:01:32.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3694" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="3728" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3740" number="3" reactiontime="+10" />
                    <RELAYPOSITION athleteid="3686" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MKS AQUATI" nation="POL" clubid="3160" name="Międzyszkolny Klub Sportowy AQUATIC" shortname="Międzyszkolny Klub Sportowy AQ">
          <CONTACT city="Gubin" email="mks@gubin.com.pl" name="Patek Ziemowit" phone="693323270" state="LUBUS" street="Piastowska 26" zip="66-620" />
          <ATHLETES>
            <ATHLETE birthdate="1953-05-24" firstname="Anna" gender="F" lastname="Krupińska" nation="POL" athleteid="3161">
              <RESULTS>
                <RESULT eventid="1222" points="182" reactiontime="+113" swimtime="00:03:57.31" resultid="3162" heatid="8968" lane="0" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.70" />
                    <SPLIT distance="100" swimtime="00:01:55.28" />
                    <SPLIT distance="150" swimtime="00:02:57.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="181" reactiontime="+102" swimtime="00:01:50.10" resultid="3163" heatid="9039" lane="9" entrytime="00:01:49.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="201" reactiontime="+113" swimtime="00:00:49.15" resultid="3164" heatid="9153" lane="4" entrytime="00:00:49.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-29" firstname="Sylwia" gender="F" lastname="Gorockiewicz" nation="POL" athleteid="3456">
              <RESULTS>
                <RESULT eventid="1222" points="109" reactiontime="+110" swimtime="00:04:41.51" resultid="3457" heatid="8967" lane="6" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.96" />
                    <SPLIT distance="100" swimtime="00:02:13.99" />
                    <SPLIT distance="150" swimtime="00:03:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="112" reactiontime="+106" swimtime="00:02:09.04" resultid="3458" heatid="9037" lane="4" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="108" reactiontime="+120" swimtime="00:01:00.38" resultid="3459" heatid="9153" lane="9" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="5601" name="MKP PD">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1968-02-22" firstname="Nina" gender="F" lastname="Hlatká" nation="SVK" athleteid="5613">
              <RESULTS>
                <RESULT eventid="1062" points="360" reactiontime="+96" swimtime="00:00:32.66" resultid="5614" heatid="8890" lane="1" entrytime="00:00:32.90" />
                <RESULT eventid="1256" points="349" reactiontime="+89" swimtime="00:01:12.41" resultid="5615" heatid="8982" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="283" reactiontime="+93" swimtime="00:00:43.86" resultid="5616" heatid="9155" lane="0" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-04-12" firstname="Mária" gender="F" lastname="Hausnerová" nation="SVK" athleteid="5607">
              <RESULTS>
                <RESULT eventid="1062" points="248" reactiontime="+85" swimtime="00:00:36.99" resultid="5608" heatid="8888" lane="2" entrytime="00:00:38.50" />
                <RESULT eventid="1187" points="193" reactiontime="+85" swimtime="00:00:44.39" resultid="5609" heatid="8950" lane="0" entrytime="00:00:46.20" />
                <RESULT eventid="1290" points="198" reactiontime="+90" swimtime="00:01:37.12" resultid="5610" heatid="9002" lane="6" entrytime="00:01:44.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="187" reactiontime="+69" swimtime="00:01:36.10" resultid="5611" heatid="9075" lane="4" entrytime="00:01:39.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="163" reactiontime="+93" swimtime="00:00:52.71" resultid="5612" heatid="9153" lane="2" entrytime="00:00:52.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" region="ZAC" clubid="2710" name="MKP Szczecin">
          <CONTACT name="Grzeszewski Sławomir" />
          <ATHLETES>
            <ATHLETE birthdate="1984-07-26" firstname="Marcin" gender="M" lastname="Gargas" nation="POL" athleteid="2724">
              <RESULTS>
                <RESULT eventid="1079" points="197" reactiontime="+111" swimtime="00:00:34.77" resultid="2725" heatid="8899" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2726" heatid="8988" lane="0" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="2718" />
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DZDZE" nation="POL" region="DOLNOSLĄSK" clubid="4731" name="MKS DZIEWIĄTKA Dzierżoniów">
          <CONTACT email="serhetabat@wp.pl" name="Piotr Kuszka" phone="604226649" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-18" firstname="Artur" gender="M" lastname="Kiraga" nation="POL" athleteid="4757">
              <RESULTS>
                <RESULT eventid="1079" points="288" reactiontime="+90" swimtime="00:00:30.65" resultid="4758" heatid="8902" lane="3" entrytime="00:00:31.18" />
                <RESULT eventid="1205" points="171" reactiontime="+68" swimtime="00:00:39.99" resultid="4759" heatid="8958" lane="8" entrytime="00:00:41.00" />
                <RESULT eventid="1273" points="261" reactiontime="+75" swimtime="00:01:10.32" resultid="4760" heatid="8990" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="250" reactiontime="+93" swimtime="00:00:34.58" resultid="4761" heatid="9064" lane="7" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-27" firstname="Ewelina" gender="F" lastname="Gutkowska" nation="POL" athleteid="4750">
              <RESULTS>
                <RESULT eventid="1062" points="412" reactiontime="+80" swimtime="00:00:31.22" resultid="4751" heatid="8891" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1096" points="311" reactiontime="+86" swimtime="00:02:59.75" resultid="4752" heatid="8920" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:22.11" />
                    <SPLIT distance="150" swimtime="00:02:14.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="399" reactiontime="+83" swimtime="00:01:09.27" resultid="4753" heatid="8982" lane="4" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="356" reactiontime="+85" swimtime="00:01:19.96" resultid="4754" heatid="9006" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="309" reactiontime="+85" swimtime="00:00:36.06" resultid="4755" heatid="9058" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1491" points="362" reactiontime="+85" swimtime="00:02:35.32" resultid="4756" heatid="9093" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="150" swimtime="00:01:53.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-05-03" firstname="Krzysztof" gender="M" lastname="Pawlaczek" nation="POL" athleteid="4762">
              <RESULTS>
                <RESULT eventid="1079" points="386" reactiontime="+78" swimtime="00:00:27.81" resultid="4763" heatid="8907" lane="4" entrytime="00:00:28.46" />
                <RESULT eventid="1239" points="357" reactiontime="+87" swimtime="00:02:49.72" resultid="4764" heatid="8977" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:22.11" />
                    <SPLIT distance="150" swimtime="00:02:06.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="388" reactiontime="+84" swimtime="00:01:09.41" resultid="4765" heatid="9017" lane="3" entrytime="00:01:10.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="4766" heatid="9051" lane="4" entrytime="00:01:17.67" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="4767" heatid="9069" lane="3" entrytime="00:00:29.96" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="4768" heatid="9170" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-04-14" firstname="Piotr" gender="M" lastname="Kuszka" nation="POL" athleteid="4769">
              <RESULTS>
                <RESULT eventid="1079" points="228" reactiontime="+74" swimtime="00:00:33.15" resultid="4770" heatid="8900" lane="9" entrytime="00:00:34.01" />
                <RESULT eventid="1239" points="201" reactiontime="+101" swimtime="00:03:25.66" resultid="4771" heatid="8974" lane="2" entrytime="00:03:21.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                    <SPLIT distance="100" swimtime="00:01:37.33" />
                    <SPLIT distance="150" swimtime="00:02:31.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="163" reactiontime="+97" swimtime="00:01:32.62" resultid="4772" heatid="9011" lane="9" entrytime="00:01:34.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="227" reactiontime="+94" swimtime="00:01:31.04" resultid="4773" heatid="9046" lane="4" entrytime="00:01:31.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="164" reactiontime="+98" swimtime="00:00:39.79" resultid="4774" heatid="9062" lane="5" entrytime="00:00:39.14" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="4775" heatid="9165" lane="2" entrytime="00:00:39.64" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00816" nation="POL" region="SZ" clubid="4485" name="MKS Neptun Stargard">
          <CONTACT city="Stargard Szcz." email="prezes@mksneptun.pl" internet="www.mksneptun.pl" name="Miedzyszkolny Klub Sportowy &quot;Neptun&quot;" phone="602731410" state="ZACHO" street="Os. Zachód B 15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1994-09-30" firstname="Mateusz" gender="M" lastname="Drozd" nation="POL" license="100816700109" athleteid="5630">
              <RESULTS>
                <RESULT eventid="1079" points="568" reactiontime="+73" swimtime="00:00:24.45" resultid="5631" heatid="8915" lane="6" entrytime="00:00:23.82" />
                <RESULT eventid="1113" points="531" reactiontime="+74" swimtime="00:02:15.35" resultid="5632" heatid="8931" lane="3" entrytime="00:02:12.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="100" swimtime="00:01:02.84" />
                    <SPLIT distance="150" swimtime="00:01:42.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="468" reactiontime="+80" swimtime="00:00:28.60" resultid="5633" heatid="8964" lane="3" entrytime="00:00:28.62" />
                <RESULT eventid="1307" points="567" reactiontime="+74" swimtime="00:01:01.19" resultid="5634" heatid="9021" lane="1" entrytime="00:01:00.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="526" reactiontime="+78" swimtime="00:00:27.00" resultid="5635" heatid="9073" lane="0" entrytime="00:00:26.60" />
                <RESULT eventid="1508" points="581" reactiontime="+73" swimtime="00:01:59.07" resultid="5636" heatid="9106" lane="5" entrytime="00:01:55.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                    <SPLIT distance="100" swimtime="00:00:57.79" />
                    <SPLIT distance="150" swimtime="00:01:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="527" reactiontime="+72" swimtime="00:00:59.95" resultid="5637" heatid="9137" lane="7" entrytime="00:00:57.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="5638" heatid="9150" lane="1" entrytime="00:02:18.44" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00811" nation="POL" region="SLA" clubid="4608" name="MKS Pałac Młodzieży Katowice">
          <CONTACT city="Katowice" email="r.puchalski@duosport.pl" name="Puchalski Robert" phone="503-684-584" state="ŚLĄSK" street="Mikołowska 26" zip="40-066" />
          <ATHLETES>
            <ATHLETE birthdate="1986-09-01" firstname="Błażej" gender="M" lastname="Kornaga" nation="POL" athleteid="4615">
              <RESULTS>
                <RESULT eventid="1079" points="363" reactiontime="+90" swimtime="00:00:28.38" resultid="4616" heatid="8906" lane="2" entrytime="00:00:29.09" />
                <RESULT eventid="1273" points="330" reactiontime="+86" swimtime="00:01:04.97" resultid="4617" heatid="8992" lane="6" entrytime="00:01:07.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-08-16" firstname="Jacek" gender="M" lastname="Syska" nation="POL" athleteid="4612">
              <RESULTS>
                <RESULT eventid="1079" points="209" reactiontime="+93" swimtime="00:00:34.13" resultid="4613" heatid="8900" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1440" points="210" reactiontime="+83" swimtime="00:00:36.67" resultid="4614" heatid="9063" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1782" name="MOSiR KSZO Ostrowiec Św.">
          <CONTACT name="Różalski" phone="510600865" street="Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" license="M01012200001" athleteid="1783">
              <RESULTS>
                <RESULT eventid="1079" points="236" reactiontime="+97" swimtime="00:00:32.74" resultid="1784" heatid="8899" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1113" points="145" reactiontime="+98" swimtime="00:03:28.22" resultid="1785" heatid="8922" lane="5" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.10" />
                    <SPLIT distance="100" swimtime="00:01:42.43" />
                    <SPLIT distance="150" swimtime="00:02:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="146" reactiontime="+108" swimtime="00:03:48.35" resultid="1786" heatid="8972" lane="1" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.90" />
                    <SPLIT distance="100" swimtime="00:01:47.44" />
                    <SPLIT distance="150" swimtime="00:02:49.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="202" reactiontime="+104" swimtime="00:01:26.27" resultid="1787" heatid="9010" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="213" reactiontime="+100" swimtime="00:00:36.47" resultid="1788" heatid="9061" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1508" points="134" reactiontime="+105" swimtime="00:03:13.76" resultid="1789" heatid="9095" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                    <SPLIT distance="100" swimtime="00:01:31.39" />
                    <SPLIT distance="150" swimtime="00:02:23.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="113" reactiontime="+104" swimtime="00:01:39.99" resultid="1790" heatid="9129" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="202" reactiontime="+100" swimtime="00:00:42.99" resultid="1791" heatid="9161" lane="4" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" region="PDK" clubid="2639" name="MOTYL -SENIOR MOSiR Stalowa Wola" shortname="MOTYL -SENIOR MOSiR Stalowa Wo">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" phone="600831914" state="PODK" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="2640">
              <RESULTS>
                <RESULT eventid="1062" points="285" reactiontime="+95" swimtime="00:00:35.29" resultid="2641" heatid="8889" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1096" points="281" reactiontime="+90" swimtime="00:03:05.89" resultid="2642" heatid="8918" lane="3" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:01:30.32" />
                    <SPLIT distance="150" swimtime="00:02:23.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="268" reactiontime="+98" swimtime="00:03:28.60" resultid="2643" heatid="8969" lane="7" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                    <SPLIT distance="100" swimtime="00:01:42.25" />
                    <SPLIT distance="150" swimtime="00:02:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="293" reactiontime="+93" swimtime="00:01:25.32" resultid="2644" heatid="9004" lane="7" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="237" swimtime="00:01:40.67" resultid="2645" heatid="9040" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="259" reactiontime="+97" swimtime="00:06:47.32" resultid="2646" heatid="9114" lane="2" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                    <SPLIT distance="100" swimtime="00:01:37.09" />
                    <SPLIT distance="150" swimtime="00:02:32.57" />
                    <SPLIT distance="200" swimtime="00:03:25.42" />
                    <SPLIT distance="250" swimtime="00:04:20.00" />
                    <SPLIT distance="300" swimtime="00:05:15.44" />
                    <SPLIT distance="350" swimtime="00:06:02.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="196" reactiontime="+95" swimtime="00:01:33.99" resultid="2647" heatid="9125" lane="8" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="288" reactiontime="+93" swimtime="00:00:43.61" resultid="2648" heatid="9155" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="2690">
              <RESULTS>
                <RESULT eventid="1079" points="284" reactiontime="+96" swimtime="00:00:30.79" resultid="2691" heatid="8904" lane="7" entrytime="00:00:30.20" />
                <RESULT eventid="1113" points="267" reactiontime="+97" swimtime="00:02:50.14" resultid="2692" heatid="8927" lane="0" entrytime="00:02:49.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:10.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="257" reactiontime="+76" swimtime="00:00:34.91" resultid="2693" heatid="8959" lane="4" entrytime="00:00:35.05" />
                <RESULT eventid="1273" points="309" reactiontime="+88" swimtime="00:01:06.43" resultid="2694" heatid="8992" lane="4" entrytime="00:01:06.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="233" reactiontime="+80" swimtime="00:01:19.46" resultid="2695" heatid="9083" lane="1" entrytime="00:01:18.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="248" reactiontime="+90" swimtime="00:06:14.53" resultid="2696" heatid="9120" lane="0" entrytime="00:06:04.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:01:27.92" />
                    <SPLIT distance="150" swimtime="00:02:15.84" />
                    <SPLIT distance="200" swimtime="00:03:01.79" />
                    <SPLIT distance="250" swimtime="00:03:56.54" />
                    <SPLIT distance="300" swimtime="00:04:51.46" />
                    <SPLIT distance="350" swimtime="00:05:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="250" reactiontime="+81" swimtime="00:02:48.36" resultid="2697" heatid="9147" lane="1" entrytime="00:02:51.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                    <SPLIT distance="100" swimtime="00:01:21.70" />
                    <SPLIT distance="150" swimtime="00:02:05.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2698" heatid="9187" lane="1" entrytime="00:05:31.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-07" firstname="Paweł" gender="M" lastname="Ciurko" nation="POL" athleteid="2649">
              <RESULTS>
                <RESULT eventid="1113" points="292" reactiontime="+96" swimtime="00:02:45.17" resultid="2650" heatid="8925" lane="7" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:22.38" />
                    <SPLIT distance="150" swimtime="00:02:06.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="323" reactiontime="+90" swimtime="00:02:55.45" resultid="2651" heatid="8975" lane="5" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:22.96" />
                    <SPLIT distance="150" swimtime="00:02:08.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="211" reactiontime="+99" swimtime="00:03:02.12" resultid="2652" heatid="9027" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:15.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="354" reactiontime="+83" swimtime="00:01:18.55" resultid="2653" heatid="9048" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="260" reactiontime="+108" swimtime="00:06:08.69" resultid="2654" heatid="9119" lane="4" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:28.69" />
                    <SPLIT distance="150" swimtime="00:02:20.10" />
                    <SPLIT distance="200" swimtime="00:03:08.74" />
                    <SPLIT distance="250" swimtime="00:03:58.38" />
                    <SPLIT distance="300" swimtime="00:04:47.47" />
                    <SPLIT distance="350" swimtime="00:05:29.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="264" reactiontime="+97" swimtime="00:01:15.47" resultid="2655" heatid="9131" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" reactiontime="+69" status="DNF" swimtime="00:00:00.00" resultid="2656" heatid="9146" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzimierz" gender="M" lastname="Jarzyna" nation="POL" athleteid="2675">
              <RESULTS>
                <RESULT eventid="1113" points="172" reactiontime="+102" swimtime="00:03:17.00" resultid="2676" heatid="8923" lane="6" entrytime="00:03:31.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                    <SPLIT distance="100" swimtime="00:01:35.04" />
                    <SPLIT distance="150" swimtime="00:02:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="153" reactiontime="+78" swimtime="00:00:41.49" resultid="2677" heatid="8957" lane="0" entrytime="00:00:43.88" />
                <RESULT eventid="1307" points="191" reactiontime="+88" swimtime="00:01:27.93" resultid="2678" heatid="9010" lane="4" entrytime="00:01:34.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="170" swimtime="00:01:28.26" resultid="2679" heatid="9081" lane="2" entrytime="00:01:33.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="177" reactiontime="+110" swimtime="00:06:58.97" resultid="2680" heatid="9118" lane="0" entrytime="00:07:20.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.03" />
                    <SPLIT distance="100" swimtime="00:01:46.79" />
                    <SPLIT distance="150" swimtime="00:02:40.77" />
                    <SPLIT distance="200" swimtime="00:03:32.47" />
                    <SPLIT distance="250" swimtime="00:04:33.19" />
                    <SPLIT distance="300" swimtime="00:05:31.40" />
                    <SPLIT distance="350" swimtime="00:06:17.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1647" points="164" reactiontime="+83" swimtime="00:03:13.63" resultid="2681" heatid="9145" lane="3" entrytime="00:03:33.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                    <SPLIT distance="100" swimtime="00:01:36.13" />
                    <SPLIT distance="150" swimtime="00:02:27.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="191" reactiontime="+99" swimtime="00:06:08.12" resultid="2682" heatid="9185" lane="9" entrytime="00:06:28.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:28.19" />
                    <SPLIT distance="150" swimtime="00:02:16.21" />
                    <SPLIT distance="200" swimtime="00:03:04.28" />
                    <SPLIT distance="250" swimtime="00:03:52.49" />
                    <SPLIT distance="300" swimtime="00:04:38.70" />
                    <SPLIT distance="350" swimtime="00:05:23.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Paweł" gender="M" lastname="Cieśliński" nation="POL" athleteid="2683">
              <RESULTS>
                <RESULT eventid="1113" points="235" reactiontime="+97" swimtime="00:02:57.42" resultid="2684" heatid="8925" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:27.92" />
                    <SPLIT distance="150" swimtime="00:02:17.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="284" reactiontime="+104" swimtime="00:03:03.16" resultid="2685" heatid="8975" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.92" />
                    <SPLIT distance="100" swimtime="00:01:29.26" />
                    <SPLIT distance="150" swimtime="00:02:16.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="208" reactiontime="+115" swimtime="00:03:03.06" resultid="2686" heatid="9028" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:29.40" />
                    <SPLIT distance="150" swimtime="00:02:17.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="286" reactiontime="+96" swimtime="00:01:24.36" resultid="2687" heatid="9050" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="2688" heatid="9132" lane="6" entrytime="00:01:20.00" />
                <RESULT eventid="1681" points="319" reactiontime="+100" swimtime="00:00:36.92" resultid="2689" heatid="9167" lane="8" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="2657">
              <RESULTS>
                <RESULT eventid="1113" points="303" reactiontime="+83" swimtime="00:02:43.09" resultid="2658" heatid="8927" lane="4" entrytime="00:02:42.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                    <SPLIT distance="150" swimtime="00:02:04.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2659" heatid="8945" lane="0" entrytime="00:21:50.30" />
                <RESULT eventid="1205" points="300" reactiontime="+75" swimtime="00:00:33.18" resultid="2660" heatid="8961" lane="3" entrytime="00:00:32.53" />
                <RESULT eventid="1307" points="335" reactiontime="+88" swimtime="00:01:12.92" resultid="2661" heatid="9016" lane="2" entrytime="00:01:12.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="282" reactiontime="+69" swimtime="00:01:14.62" resultid="2662" heatid="9084" lane="7" entrytime="00:01:12.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="270" reactiontime="+101" swimtime="00:06:04.29" resultid="2663" heatid="9120" lane="8" entrytime="00:06:03.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:26.47" />
                    <SPLIT distance="150" swimtime="00:02:14.07" />
                    <SPLIT distance="200" swimtime="00:03:00.31" />
                    <SPLIT distance="250" swimtime="00:03:51.89" />
                    <SPLIT distance="300" swimtime="00:04:43.91" />
                    <SPLIT distance="350" swimtime="00:05:25.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="237" reactiontime="+71" swimtime="00:02:51.37" resultid="2664" heatid="9148" lane="9" entrytime="00:02:41.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:23.27" />
                    <SPLIT distance="150" swimtime="00:02:07.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="300" reactiontime="+90" swimtime="00:05:16.93" resultid="2665" heatid="9187" lane="5" entrytime="00:05:27.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:52.19" />
                    <SPLIT distance="200" swimtime="00:02:33.41" />
                    <SPLIT distance="250" swimtime="00:03:15.23" />
                    <SPLIT distance="300" swimtime="00:03:56.99" />
                    <SPLIT distance="350" swimtime="00:04:37.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="2699">
              <RESULTS>
                <RESULT eventid="1079" points="476" reactiontime="+76" swimtime="00:00:25.93" resultid="2700" heatid="8914" lane="1" entrytime="00:00:25.89" />
                <RESULT eventid="1113" points="508" reactiontime="+76" swimtime="00:02:17.32" resultid="2701" heatid="8931" lane="7" entrytime="00:02:17.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                    <SPLIT distance="100" swimtime="00:01:04.69" />
                    <SPLIT distance="150" swimtime="00:01:44.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="506" reactiontime="+76" swimtime="00:00:56.37" resultid="2702" heatid="9000" lane="8" entrytime="00:00:55.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="522" reactiontime="+80" swimtime="00:01:02.89" resultid="2703" heatid="9020" lane="2" entrytime="00:01:03.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="509" reactiontime="+75" swimtime="00:00:27.29" resultid="2704" heatid="9072" lane="6" entrytime="00:00:27.19" />
                <RESULT eventid="1508" points="514" reactiontime="+77" swimtime="00:02:04.02" resultid="2705" heatid="9105" lane="5" entrytime="00:02:05.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                    <SPLIT distance="100" swimtime="00:01:01.26" />
                    <SPLIT distance="150" swimtime="00:01:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="540" reactiontime="+71" swimtime="00:00:59.47" resultid="2706" heatid="9137" lane="9" entrytime="00:00:59.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="458" reactiontime="+82" swimtime="00:00:32.74" resultid="2707" heatid="9172" lane="0" entrytime="00:00:32.59" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="2666">
              <RESULTS>
                <RESULT eventid="1079" points="448" reactiontime="+93" swimtime="00:00:26.47" resultid="2667" heatid="8912" lane="8" entrytime="00:00:26.47" />
                <RESULT eventid="1113" points="385" reactiontime="+85" swimtime="00:02:30.57" resultid="2668" heatid="8930" lane="9" entrytime="00:02:28.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:10.17" />
                    <SPLIT distance="150" swimtime="00:01:55.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="438" reactiontime="+74" swimtime="00:00:29.24" resultid="2669" heatid="8964" lane="8" entrytime="00:00:29.96" />
                <RESULT eventid="1273" points="445" reactiontime="+90" swimtime="00:00:58.82" resultid="2670" heatid="8998" lane="6" entrytime="00:00:58.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="358" reactiontime="+91" swimtime="00:00:30.69" resultid="2671" heatid="9068" lane="4" entrytime="00:00:30.03" />
                <RESULT eventid="1474" points="435" reactiontime="+77" swimtime="00:01:04.58" resultid="2672" heatid="9086" lane="6" entrytime="00:01:05.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="389" reactiontime="+79" swimtime="00:02:25.34" resultid="2673" heatid="9149" lane="3" entrytime="00:02:26.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:11.70" />
                    <SPLIT distance="150" swimtime="00:01:49.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="337" reactiontime="+85" swimtime="00:00:36.27" resultid="2674" heatid="9168" lane="4" entrytime="00:00:36.49" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="377" reactiontime="+75" swimtime="00:01:54.32" resultid="2708" heatid="9111" lane="2" entrytime="00:01:53.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                    <SPLIT distance="100" swimtime="00:00:58.05" />
                    <SPLIT distance="150" swimtime="00:01:28.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2699" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="2675" number="2" />
                    <RELAYPOSITION athleteid="2690" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2666" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="339" reactiontime="+60" swimtime="00:02:09.74" resultid="2709" heatid="9034" lane="9" entrytime="00:02:11.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                    <SPLIT distance="150" swimtime="00:01:37.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2666" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="2690" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="2699" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="2675" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="5639" name="MSC &quot;Euro-Lviv&quot;">
          <CONTACT city="Lviv" email="riff@mail.lviv.ua" fax="+380322430304" name="Ruslan Friauf" phone="+380676734796" street="Karpincya 18A/3" zip="79012" />
          <ATHLETES>
            <ATHLETE birthdate="1932-06-01" firstname="Serhiy" gender="M" lastname="Simankov" nation="UKR" athleteid="5733">
              <RESULTS>
                <RESULT eventid="1079" points="110" reactiontime="+122" swimtime="00:00:42.20" resultid="5734" heatid="8897" lane="0" entrytime="00:00:40.30" />
                <RESULT eventid="1341" points="57" reactiontime="+135" swimtime="00:04:40.84" resultid="5735" heatid="9025" lane="4" entrytime="00:04:47.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.02" />
                    <SPLIT distance="100" swimtime="00:02:11.46" />
                    <SPLIT distance="150" swimtime="00:03:28.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="97" reactiontime="+115" swimtime="00:00:47.43" resultid="5736" heatid="9061" lane="1" entrytime="00:00:47.10" />
                <RESULT eventid="1613" points="63" reactiontime="+123" swimtime="00:02:01.56" resultid="5737" heatid="9129" lane="2" entrytime="00:02:04.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="105" reactiontime="+112" swimtime="00:00:53.41" resultid="5738" heatid="9160" lane="4" entrytime="00:00:54.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-28" firstname="Valentyna" gender="F" lastname="Kvita" nation="UKR" athleteid="5654">
              <RESULTS>
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="5655" heatid="8939" lane="6" entrytime="00:10:35.00" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="5656" heatid="8984" lane="7" entrytime="00:01:02.90" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="5657" heatid="9093" lane="2" entrytime="00:02:21.00" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="5658" heatid="9181" lane="6" entrytime="00:04:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-06" firstname="Mariya" gender="F" lastname="Vasylko" nation="UKR" athleteid="5674">
              <RESULTS>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="5675" heatid="8949" lane="7" entrytime="00:00:52.00" />
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="5676" heatid="9055" lane="4" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-18" firstname="Dmytro" gender="M" lastname="Melnyk" nation="UKR" athleteid="5710">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="5711" heatid="8911" lane="6" entrytime="00:00:26.55" />
                <RESULT eventid="1406" points="403" reactiontime="+77" swimtime="00:01:15.28" resultid="5712" heatid="9052" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="382" reactiontime="+80" swimtime="00:00:30.02" resultid="5713" heatid="9069" lane="5" entrytime="00:00:29.80" />
                <RESULT eventid="1681" points="443" reactiontime="+74" swimtime="00:00:33.10" resultid="5714" heatid="9171" lane="7" entrytime="00:00:33.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-18" firstname="Vladyslav" gender="M" lastname="Horovoy" nation="UKR" athleteid="5685">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5686" heatid="8963" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="5687" heatid="8999" lane="3" entrytime="00:00:57.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="5688" heatid="9105" lane="1" entrytime="00:02:08.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="5689" heatid="9192" lane="2" entrytime="00:04:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-02-27" firstname="Olena" gender="F" lastname="Pereyaslova" nation="UKR" athleteid="5667">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="5668" heatid="8918" lane="2" entrytime="00:03:15.00" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="5669" heatid="8981" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="5670" heatid="9091" lane="6" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-31" firstname="Roman" gender="M" lastname="Koretskyy" nation="UKR" athleteid="5702" />
            <ATHLETE birthdate="1976-02-03" firstname="Romana" gender="F" lastname="Sirenko" nation="UKR" athleteid="5671">
              <RESULTS>
                <RESULT eventid="1187" points="299" reactiontime="+78" swimtime="00:00:38.38" resultid="5672" heatid="8951" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1423" points="293" swimtime="00:00:36.70" resultid="5673" heatid="9057" lane="7" entrytime="00:00:35.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-05-09" firstname="Lidiya" gender="F" lastname="Tymoshenko" nation="UKR" athleteid="5662">
              <RESULTS>
                <RESULT eventid="1062" points="113" reactiontime="+134" swimtime="00:00:47.93" resultid="5663" heatid="8886" lane="3" entrytime="00:00:49.09" />
                <RESULT eventid="1388" points="116" reactiontime="+109" swimtime="00:02:07.72" resultid="5664" heatid="9038" lane="9" entrytime="00:02:06.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="87" reactiontime="+121" swimtime="00:01:55.08" resultid="5665" heatid="8979" lane="1" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="144" reactiontime="+101" swimtime="00:00:54.88" resultid="5666" heatid="9152" lane="5" entrytime="00:00:58.34" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-22" firstname="Volodymyr" gender="M" lastname="Rybko" nation="UKR" athleteid="5717">
              <RESULTS>
                <RESULT eventid="1165" points="347" reactiontime="+91" swimtime="00:20:08.60" resultid="5718" heatid="8946" lane="4" entrytime="00:20:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:01:53.22" />
                    <SPLIT distance="200" swimtime="00:02:33.23" />
                    <SPLIT distance="250" swimtime="00:03:12.66" />
                    <SPLIT distance="300" swimtime="00:03:52.62" />
                    <SPLIT distance="350" swimtime="00:04:32.88" />
                    <SPLIT distance="400" swimtime="00:05:12.97" />
                    <SPLIT distance="450" swimtime="00:05:52.34" />
                    <SPLIT distance="500" swimtime="00:06:31.70" />
                    <SPLIT distance="550" swimtime="00:07:11.58" />
                    <SPLIT distance="600" swimtime="00:07:51.93" />
                    <SPLIT distance="650" swimtime="00:08:32.07" />
                    <SPLIT distance="700" swimtime="00:09:12.62" />
                    <SPLIT distance="750" swimtime="00:09:54.72" />
                    <SPLIT distance="800" swimtime="00:10:35.29" />
                    <SPLIT distance="850" swimtime="00:11:15.13" />
                    <SPLIT distance="900" swimtime="00:11:55.21" />
                    <SPLIT distance="950" swimtime="00:12:35.06" />
                    <SPLIT distance="1000" swimtime="00:13:16.29" />
                    <SPLIT distance="1050" swimtime="00:13:56.53" />
                    <SPLIT distance="1100" swimtime="00:14:36.19" />
                    <SPLIT distance="1150" swimtime="00:15:17.47" />
                    <SPLIT distance="1200" swimtime="00:15:58.70" />
                    <SPLIT distance="1250" swimtime="00:16:40.01" />
                    <SPLIT distance="1300" swimtime="00:17:20.61" />
                    <SPLIT distance="1350" swimtime="00:18:00.36" />
                    <SPLIT distance="1400" swimtime="00:18:41.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="347" reactiontime="+83" swimtime="00:01:12.04" resultid="5719" heatid="9018" lane="6" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="296" reactiontime="+81" swimtime="00:05:53.28" resultid="5720" heatid="9120" lane="5" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:01:22.75" />
                    <SPLIT distance="150" swimtime="00:02:07.99" />
                    <SPLIT distance="200" swimtime="00:02:53.76" />
                    <SPLIT distance="250" swimtime="00:03:46.17" />
                    <SPLIT distance="300" swimtime="00:04:39.42" />
                    <SPLIT distance="350" swimtime="00:05:17.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="268" reactiontime="+77" swimtime="00:01:15.06" resultid="5721" heatid="9135" lane="7" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="358" reactiontime="+82" swimtime="00:04:58.87" resultid="5722" heatid="9189" lane="7" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:50.78" />
                    <SPLIT distance="200" swimtime="00:02:29.64" />
                    <SPLIT distance="250" swimtime="00:03:07.95" />
                    <SPLIT distance="300" swimtime="00:03:46.76" />
                    <SPLIT distance="350" swimtime="00:04:25.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-04-06" firstname="Sergiy" gender="M" lastname="Mashkin" nation="UKR" athleteid="5705">
              <RESULTS>
                <RESULT eventid="1079" points="243" reactiontime="+96" swimtime="00:00:32.45" resultid="5706" heatid="8906" lane="8" entrytime="00:00:29.50" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="5707" heatid="8992" lane="7" entrytime="00:01:07.50" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="5708" heatid="9066" lane="9" entrytime="00:00:33.20" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="5709" heatid="9147" lane="7" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-27" firstname="Oleh" gender="M" lastname="Biront" nation="UKR" athleteid="5677">
              <RESULTS>
                <RESULT eventid="1079" points="229" reactiontime="+110" swimtime="00:00:33.08" resultid="5678" heatid="8901" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1239" points="198" reactiontime="+106" swimtime="00:03:26.62" resultid="5679" heatid="8973" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                    <SPLIT distance="100" swimtime="00:01:37.57" />
                    <SPLIT distance="150" swimtime="00:02:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="210" reactiontime="+93" swimtime="00:01:33.54" resultid="5680" heatid="9048" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="251" reactiontime="+106" swimtime="00:00:39.99" resultid="5681" heatid="9164" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-06" firstname="Lyudmyla" gender="F" lastname="Khiresh" nation="UKR" athleteid="5649" />
            <ATHLETE birthdate="1954-06-05" firstname="Mykhailo" gender="M" lastname="Shelest" nation="UKR" athleteid="5723">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5724" heatid="8959" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="5725" heatid="8974" lane="6" entrytime="00:03:20.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="5726" heatid="9049" lane="0" entrytime="00:01:27.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="5727" heatid="9167" lane="7" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-02" firstname="Serhiy" gender="M" lastname="Zhykh" nation="UKR" athleteid="5739" />
            <ATHLETE birthdate="1972-09-13" firstname="Oleksandr" gender="M" lastname="Syrbu" nation="UKR" athleteid="5728">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="5729" heatid="8914" lane="9" entrytime="00:00:25.95" />
                <RESULT eventid="1273" points="475" reactiontime="+80" swimtime="00:00:57.57" resultid="5730" heatid="8999" lane="5" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="519" reactiontime="+79" swimtime="00:00:27.12" resultid="5731" heatid="9072" lane="2" entrytime="00:00:27.20" />
                <RESULT eventid="1613" points="441" reactiontime="+91" swimtime="00:01:03.62" resultid="5732" heatid="9136" lane="0" entrytime="00:01:03.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-13" firstname="Bohdan" gender="M" lastname="Osidach" nation="UKR" athleteid="5715" />
            <ATHLETE birthdate="1949-03-31" firstname="Myron" gender="M" lastname="Kolodko" nation="UKR" athleteid="5696">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="5697" heatid="8923" lane="7" entrytime="00:03:39.00" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="5698" heatid="9026" lane="7" entrytime="00:04:15.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="5699" heatid="9062" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="5700" heatid="9117" lane="5" entrytime="00:07:45.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="5701" heatid="9130" lane="1" entrytime="00:01:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-11-30" firstname="Tetiana" gender="F" lastname="Kozakova" nation="UKR" athleteid="5659" />
            <ATHLETE birthdate="1952-07-12" firstname="Petro" gender="M" lastname="Gemba" nation="UKR" athleteid="5644">
              <RESULTS>
                <RESULT eventid="1165" points="249" reactiontime="+96" swimtime="00:22:30.50" resultid="5645" heatid="8943" lane="5" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:09.45" />
                    <SPLIT distance="200" swimtime="00:02:54.58" />
                    <SPLIT distance="250" swimtime="00:03:40.12" />
                    <SPLIT distance="300" swimtime="00:04:25.73" />
                    <SPLIT distance="350" swimtime="00:05:11.05" />
                    <SPLIT distance="400" swimtime="00:05:56.33" />
                    <SPLIT distance="450" swimtime="00:06:40.87" />
                    <SPLIT distance="500" swimtime="00:07:25.51" />
                    <SPLIT distance="550" swimtime="00:08:10.53" />
                    <SPLIT distance="600" swimtime="00:08:55.74" />
                    <SPLIT distance="650" swimtime="00:09:41.36" />
                    <SPLIT distance="700" swimtime="00:10:26.48" />
                    <SPLIT distance="750" swimtime="00:11:11.25" />
                    <SPLIT distance="800" swimtime="00:11:56.54" />
                    <SPLIT distance="850" swimtime="00:12:42.01" />
                    <SPLIT distance="900" swimtime="00:13:27.26" />
                    <SPLIT distance="950" swimtime="00:14:12.29" />
                    <SPLIT distance="1000" swimtime="00:14:57.41" />
                    <SPLIT distance="1050" swimtime="00:15:42.30" />
                    <SPLIT distance="1100" swimtime="00:16:27.97" />
                    <SPLIT distance="1150" swimtime="00:17:13.47" />
                    <SPLIT distance="1200" swimtime="00:17:59.41" />
                    <SPLIT distance="1250" swimtime="00:18:45.03" />
                    <SPLIT distance="1300" swimtime="00:19:30.69" />
                    <SPLIT distance="1350" swimtime="00:20:16.73" />
                    <SPLIT distance="1400" swimtime="00:21:02.49" />
                    <SPLIT distance="1450" swimtime="00:21:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="191" reactiontime="+89" swimtime="00:01:27.83" resultid="5646" heatid="9011" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="215" reactiontime="+93" swimtime="00:02:45.75" resultid="5647" heatid="9098" lane="8" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:19.75" />
                    <SPLIT distance="150" swimtime="00:02:02.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="233" reactiontime="+97" swimtime="00:05:44.78" resultid="5648" heatid="9186" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                    <SPLIT distance="150" swimtime="00:02:09.53" />
                    <SPLIT distance="200" swimtime="00:02:53.56" />
                    <SPLIT distance="250" swimtime="00:03:37.27" />
                    <SPLIT distance="300" swimtime="00:04:19.84" />
                    <SPLIT distance="350" swimtime="00:05:02.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-05-31" firstname="Zenoviy" gender="M" lastname="Kushnir" nation="UKR" athleteid="5640">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5641" heatid="8955" lane="6" entrytime="00:00:58.80" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="5642" heatid="9044" lane="2" entrytime="00:02:08.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="5643" heatid="9144" lane="8" entrytime="00:04:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yuriy" gender="M" lastname="Denisov" nation="UKR" athleteid="5682" />
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="Friauf" nation="UKR" athleteid="5690" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="5743" heatid="9035" lane="1" entrytime="00:01:58.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5728" number="1" />
                    <RELAYPOSITION athleteid="5710" number="2" />
                    <RELAYPOSITION athleteid="5677" number="3" />
                    <RELAYPOSITION athleteid="5717" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1548" points="394" reactiontime="+80" swimtime="00:01:52.60" resultid="5744" heatid="9112" lane="0" entrytime="00:01:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.02" />
                    <SPLIT distance="100" swimtime="00:00:52.76" />
                    <SPLIT distance="150" swimtime="00:01:25.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5685" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5710" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="5717" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="5728" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="5742" heatid="8935" lane="2" entrytime="00:01:56.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5728" number="1" />
                    <RELAYPOSITION athleteid="5710" number="2" />
                    <RELAYPOSITION athleteid="5667" number="3" />
                    <RELAYPOSITION athleteid="5654" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+71" status="DNS" swimtime="00:00:00.00" resultid="5745" heatid="8934" lane="3" entrytime="00:02:06.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:31.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5654" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5710" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="5728" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5667" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2969" name="MSwim Szczecin">
          <CONTACT city="Wołczkowo" email="m@mswim.pl" internet="www.mswim.pl" name="Kaczanowski Miłosz" phone="888 18 1234" street="Słoneczna 5" zip="72-003" />
          <ATHLETES>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="2986">
              <RESULTS>
                <RESULT eventid="1187" points="237" reactiontime="+82" swimtime="00:00:41.45" resultid="2987" heatid="8950" lane="7" entrytime="00:00:42.50" />
                <RESULT eventid="1457" points="244" reactiontime="+82" swimtime="00:01:28.03" resultid="2988" heatid="9076" lane="8" entrytime="00:01:30.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="245" reactiontime="+89" swimtime="00:03:10.50" resultid="2989" heatid="9139" lane="5" entrytime="00:03:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:32.08" />
                    <SPLIT distance="150" swimtime="00:02:21.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-10-12" firstname="Zbigniew" gender="M" lastname="Szozda" nation="POL" athleteid="2977">
              <RESULTS>
                <RESULT eventid="1205" points="233" reactiontime="+135" swimtime="00:00:36.08" resultid="2980" heatid="8959" lane="1" entrytime="00:00:36.50" />
                <RESULT eventid="1239" points="238" reactiontime="+105" swimtime="00:03:14.30" resultid="2981" heatid="8975" lane="9" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                    <SPLIT distance="100" swimtime="00:01:31.82" />
                    <SPLIT distance="150" swimtime="00:02:22.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="2982" heatid="9048" lane="6" entrytime="00:01:29.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="2983" heatid="9083" lane="9" entrytime="00:01:20.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="2984" heatid="9131" lane="4" entrytime="00:01:25.00" />
                <RESULT eventid="1647" points="195" reactiontime="+81" swimtime="00:03:02.81" resultid="2985" heatid="9146" lane="5" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="150" swimtime="00:02:13.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01511" nation="POL" region="SLA" clubid="2229" name="MTP Delfin Cieszyn">
          <CONTACT city="Cieszyn" email="k.widzik@delfincieszyn.pl" name="Widzik Katarzyna" phone="735951829" state="11" street="Plac Wolności  7a" zip="43-400" />
          <ATHLETES>
            <ATHLETE birthdate="1990-06-12" firstname="Katarzyna" gender="F" lastname="Widzik" nation="POL" athleteid="2230">
              <RESULTS>
                <RESULT eventid="1147" points="431" reactiontime="+84" swimtime="00:10:34.30" resultid="2231" heatid="8936" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:14.30" />
                    <SPLIT distance="150" swimtime="00:01:53.74" />
                    <SPLIT distance="200" swimtime="00:02:32.72" />
                    <SPLIT distance="250" swimtime="00:03:12.63" />
                    <SPLIT distance="300" swimtime="00:03:52.69" />
                    <SPLIT distance="350" swimtime="00:04:33.06" />
                    <SPLIT distance="400" swimtime="00:05:13.63" />
                    <SPLIT distance="450" swimtime="00:05:54.11" />
                    <SPLIT distance="500" swimtime="00:06:34.68" />
                    <SPLIT distance="550" swimtime="00:07:15.24" />
                    <SPLIT distance="600" swimtime="00:07:55.74" />
                    <SPLIT distance="650" swimtime="00:08:35.56" />
                    <SPLIT distance="700" swimtime="00:09:16.10" />
                    <SPLIT distance="750" swimtime="00:09:55.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="374" reactiontime="+79" swimtime="00:03:06.71" resultid="2232" heatid="8969" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:29.23" />
                    <SPLIT distance="150" swimtime="00:02:17.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="319" reactiontime="+81" swimtime="00:02:54.88" resultid="2233" heatid="9023" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:23.40" />
                    <SPLIT distance="150" swimtime="00:02:08.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="407" reactiontime="+66" swimtime="00:01:14.24" resultid="2234" heatid="9078" lane="2" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" status="DNS" swimtime="00:00:00.00" resultid="2235" heatid="9114" lane="6" entrytime="00:06:45.00" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="2236" heatid="9141" lane="1" entrytime="00:02:45.00" />
                <RESULT eventid="1721" points="436" reactiontime="+76" swimtime="00:05:09.17" resultid="2237" heatid="9181" lane="5" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:51.89" />
                    <SPLIT distance="200" swimtime="00:02:31.58" />
                    <SPLIT distance="250" swimtime="00:03:11.27" />
                    <SPLIT distance="300" swimtime="00:03:51.21" />
                    <SPLIT distance="350" swimtime="00:04:30.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1776" name="Neptun Team Tarnów">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1986-06-23" firstname="Mateusz" gender="M" lastname="Dymiter" nation="POL" athleteid="1777">
              <RESULTS>
                <RESULT eventid="1239" points="366" reactiontime="+94" swimtime="00:02:48.32" resultid="1778" heatid="8975" lane="3" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:03.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="392" reactiontime="+90" swimtime="00:01:09.19" resultid="1779" heatid="9016" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="1780" heatid="9083" lane="0" entrytime="00:01:19.00" />
                <RESULT eventid="1578" points="340" reactiontime="+101" swimtime="00:05:37.14" resultid="1781" heatid="9120" lane="1" entrytime="00:06:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="150" swimtime="00:01:56.08" />
                    <SPLIT distance="200" swimtime="00:02:40.15" />
                    <SPLIT distance="250" swimtime="00:03:27.86" />
                    <SPLIT distance="300" swimtime="00:04:15.78" />
                    <SPLIT distance="350" swimtime="00:04:58.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" clubid="1761" name="Niezrzeszeni">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1986-08-06" firstname="Oleksandr" gender="M" lastname="Broshevan" nation="POL" athleteid="1931">
              <RESULTS>
                <RESULT eventid="1079" points="382" reactiontime="+99" swimtime="00:00:27.91" resultid="1932" heatid="8911" lane="7" entrytime="00:00:26.66" />
                <RESULT eventid="1273" points="309" reactiontime="+87" swimtime="00:01:06.43" resultid="1933" heatid="8994" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="339" reactiontime="+101" swimtime="00:01:12.63" resultid="1934" heatid="9015" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M12 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 17:15)" eventid="1440" reactiontime="+99" status="DSQ" swimtime="00:00:29.58" resultid="1935" heatid="9071" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1681" points="295" reactiontime="+89" swimtime="00:00:37.89" resultid="1936" heatid="9165" lane="9" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-03-15" firstname="Jiří" gender="M" lastname="Janovský " nation="CZE" athleteid="8879">
              <RESULTS>
                <RESULT eventid="1165" points="316" reactiontime="+103" swimtime="00:20:47.80" resultid="8880" heatid="8944" lane="7" entrytime="00:22:11.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:16.36" />
                    <SPLIT distance="150" swimtime="00:01:56.87" />
                    <SPLIT distance="200" swimtime="00:03:18.37" />
                    <SPLIT distance="250" swimtime="00:04:00.12" />
                    <SPLIT distance="300" swimtime="00:04:40.81" />
                    <SPLIT distance="350" swimtime="00:05:22.10" />
                    <SPLIT distance="400" swimtime="00:06:04.09" />
                    <SPLIT distance="450" swimtime="00:06:45.71" />
                    <SPLIT distance="500" swimtime="00:07:27.72" />
                    <SPLIT distance="550" swimtime="00:08:09.58" />
                    <SPLIT distance="600" swimtime="00:08:51.83" />
                    <SPLIT distance="650" swimtime="00:09:34.29" />
                    <SPLIT distance="700" swimtime="00:10:16.12" />
                    <SPLIT distance="750" swimtime="00:10:58.33" />
                    <SPLIT distance="800" swimtime="00:11:41.21" />
                    <SPLIT distance="850" swimtime="00:12:23.53" />
                    <SPLIT distance="900" swimtime="00:13:05.92" />
                    <SPLIT distance="950" swimtime="00:13:48.59" />
                    <SPLIT distance="1000" swimtime="00:15:13.35" />
                    <SPLIT distance="1050" swimtime="00:16:38.32" />
                    <SPLIT distance="1100" swimtime="00:19:26.65" />
                    <SPLIT distance="1150" swimtime="00:20:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="196" swimtime="00:00:38.20" resultid="8881" heatid="8959" lane="7" entrytime="00:00:36.50" />
                <RESULT eventid="1440" points="259" reactiontime="+95" swimtime="00:00:34.16" resultid="8882" heatid="9065" lane="4" entrytime="00:00:33.50" />
                <RESULT eventid="1578" points="262" reactiontime="+107" swimtime="00:06:07.90" resultid="8883" heatid="9119" lane="7" entrytime="00:06:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:22.51" />
                    <SPLIT distance="150" swimtime="00:02:09.89" />
                    <SPLIT distance="200" swimtime="00:02:56.01" />
                    <SPLIT distance="250" swimtime="00:03:51.90" />
                    <SPLIT distance="300" swimtime="00:04:48.89" />
                    <SPLIT distance="350" swimtime="00:05:29.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="321" reactiontime="+106" swimtime="00:05:09.97" resultid="8884" heatid="9188" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:52.25" />
                    <SPLIT distance="200" swimtime="00:02:31.60" />
                    <SPLIT distance="250" swimtime="00:03:50.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-23" firstname="Staravoitau" gender="M" lastname="Aliaksei" nation="BLR" athleteid="1923">
              <RESULTS>
                <RESULT eventid="1079" points="224" reactiontime="+113" swimtime="00:00:33.32" resultid="1924" heatid="8900" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1681" points="229" reactiontime="+108" swimtime="00:00:41.25" resultid="1925" heatid="9163" lane="2" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-10-01" firstname="Jozef" gender="M" lastname="Král" nation="SVK" athleteid="1926">
              <RESULTS>
                <RESULT eventid="1113" points="138" reactiontime="+107" swimtime="00:03:31.67" resultid="1927" heatid="8923" lane="4" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                    <SPLIT distance="100" swimtime="00:01:44.33" />
                    <SPLIT distance="150" swimtime="00:02:43.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="117" reactiontime="+104" swimtime="00:03:41.49" resultid="1928" heatid="9027" lane="2" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                    <SPLIT distance="100" swimtime="00:01:44.96" />
                    <SPLIT distance="150" swimtime="00:02:45.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="164" reactiontime="+100" swimtime="00:00:39.76" resultid="1929" heatid="9063" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1613" points="160" reactiontime="+101" swimtime="00:01:29.18" resultid="1930" heatid="9131" lane="8" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-26" firstname="Alshevich" gender="M" lastname="Andrei" nation="BLR" athleteid="1920">
              <RESULTS>
                <RESULT eventid="1079" points="439" reactiontime="+96" swimtime="00:00:26.65" resultid="1921" heatid="8912" lane="3" entrytime="00:00:26.30" />
                <RESULT eventid="1440" points="441" reactiontime="+93" swimtime="00:00:28.63" resultid="1922" heatid="9070" lane="4" entrytime="00:00:28.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3046" name="Niezrzeszeni ">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1985-09-25" firstname="Sandro" gender="M" lastname="Surwiło" nation="POL" athleteid="4199">
              <RESULTS>
                <RESULT eventid="1079" points="338" reactiontime="+101" swimtime="00:00:29.07" resultid="4200" heatid="8901" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1273" points="278" reactiontime="+100" swimtime="00:01:08.81" resultid="4201" heatid="8990" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="250" reactiontime="+108" swimtime="00:02:37.57" resultid="4202" heatid="9099" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:53.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-03-17" firstname="Przemysław" gender="M" lastname="Pobóg-Zarzecki" nation="POL" athleteid="6350">
              <RESULTS>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="6351" heatid="8991" lane="2" entrytime="00:01:10.00" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="6352" heatid="9013" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="6353" heatid="9165" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-10-29" firstname="Mateusz" gender="M" lastname="Czarnota" nation="POL" athleteid="2256">
              <RESULTS>
                <RESULT eventid="1113" points="608" reactiontime="+75" swimtime="00:02:09.39" resultid="2257" heatid="8921" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="100" swimtime="00:01:00.65" />
                    <SPLIT distance="150" swimtime="00:01:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" reactiontime="+73" status="DNF" swimtime="00:00:00.00" resultid="2258" heatid="8940" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.74" />
                    <SPLIT distance="100" swimtime="00:00:56.00" />
                    <SPLIT distance="150" swimtime="00:01:25.74" />
                    <SPLIT distance="200" swimtime="00:01:55.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="638" reactiontime="+75" swimtime="00:01:55.37" resultid="2259" heatid="9094" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                    <SPLIT distance="100" swimtime="00:00:55.68" />
                    <SPLIT distance="150" swimtime="00:01:25.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="636" reactiontime="+72" swimtime="00:04:33.74" resultid="2260" heatid="9116" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:03.93" />
                    <SPLIT distance="150" swimtime="00:01:39.82" />
                    <SPLIT distance="200" swimtime="00:02:15.09" />
                    <SPLIT distance="250" swimtime="00:02:53.74" />
                    <SPLIT distance="300" swimtime="00:03:32.47" />
                    <SPLIT distance="350" swimtime="00:04:03.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-30" firstname="Arkadiusz" gender="M" lastname="Kawalec" nation="POL" athleteid="6181">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="6182" heatid="8913" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="6183" heatid="9071" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="6184" heatid="9171" lane="9" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-27" firstname="Weronika" gender="F" lastname="Kabut" nation="POL" athleteid="4182">
              <RESULTS>
                <RESULT eventid="1062" points="458" reactiontime="+79" swimtime="00:00:30.14" resultid="4183" heatid="8891" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1256" points="433" reactiontime="+79" swimtime="00:01:07.39" resultid="4184" heatid="8983" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="372" reactiontime="+79" swimtime="00:01:18.77" resultid="4185" heatid="9005" lane="8" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="301" reactiontime="+86" swimtime="00:01:33.04" resultid="4186" heatid="9040" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="342" reactiontime="+83" swimtime="00:00:34.85" resultid="4187" heatid="9057" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-03-28" firstname="Katarzyna" gender="F" lastname="Wnęk" nation="POL" athleteid="4175">
              <RESULTS>
                <RESULT eventid="1222" points="349" reactiontime="+93" swimtime="00:03:10.96" resultid="4176" heatid="8970" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                    <SPLIT distance="100" swimtime="00:01:30.39" />
                    <SPLIT distance="150" swimtime="00:02:19.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="391" reactiontime="+101" swimtime="00:01:09.74" resultid="4177" heatid="8982" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="357" reactiontime="+83" swimtime="00:01:27.90" resultid="4178" heatid="9041" lane="9" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="360" reactiontime="+87" swimtime="00:02:35.71" resultid="4179" heatid="9092" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:14.61" />
                    <SPLIT distance="150" swimtime="00:01:55.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="353" reactiontime="+92" swimtime="00:00:40.72" resultid="4180" heatid="9157" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1721" points="318" reactiontime="+101" swimtime="00:05:43.55" resultid="4181" heatid="9180" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                    <SPLIT distance="100" swimtime="00:01:21.70" />
                    <SPLIT distance="150" swimtime="00:02:04.83" />
                    <SPLIT distance="200" swimtime="00:02:48.84" />
                    <SPLIT distance="250" swimtime="00:03:33.39" />
                    <SPLIT distance="300" swimtime="00:04:17.98" />
                    <SPLIT distance="350" swimtime="00:05:03.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-09-24" firstname="Daria" gender="F" lastname="Radczuk" nation="POL" athleteid="3375">
              <RESULTS>
                <RESULT eventid="1062" points="409" reactiontime="+91" swimtime="00:00:31.30" resultid="3376" heatid="8891" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1147" points="450" reactiontime="+91" swimtime="00:10:25.48" resultid="3377" heatid="8939" lane="7" entrytime="00:11:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:13.65" />
                    <SPLIT distance="150" swimtime="00:01:52.85" />
                    <SPLIT distance="200" swimtime="00:02:32.69" />
                    <SPLIT distance="250" swimtime="00:03:12.65" />
                    <SPLIT distance="300" swimtime="00:03:52.96" />
                    <SPLIT distance="350" swimtime="00:04:33.18" />
                    <SPLIT distance="400" swimtime="00:05:13.46" />
                    <SPLIT distance="450" swimtime="00:05:52.75" />
                    <SPLIT distance="500" swimtime="00:06:32.34" />
                    <SPLIT distance="550" swimtime="00:07:11.63" />
                    <SPLIT distance="600" swimtime="00:07:51.14" />
                    <SPLIT distance="650" swimtime="00:08:30.56" />
                    <SPLIT distance="700" swimtime="00:09:09.43" />
                    <SPLIT distance="750" swimtime="00:09:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="445" reactiontime="+84" swimtime="00:01:06.81" resultid="3378" heatid="8984" lane="9" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="381" reactiontime="+88" swimtime="00:02:44.92" resultid="3379" heatid="9024" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:18.57" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="466" reactiontime="+90" swimtime="00:05:02.44" resultid="3380" heatid="9181" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:50.94" />
                    <SPLIT distance="200" swimtime="00:02:29.81" />
                    <SPLIT distance="250" swimtime="00:03:08.83" />
                    <SPLIT distance="300" swimtime="00:03:47.93" />
                    <SPLIT distance="350" swimtime="00:04:26.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-11-21" firstname="Zbigniew" gender="M" lastname="Dymecki" nation="POL" athleteid="1878">
              <RESULTS>
                <RESULT eventid="1079" points="84" reactiontime="+95" swimtime="00:00:46.23" resultid="1879" heatid="8896" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1113" points="60" reactiontime="+108" swimtime="00:04:39.25" resultid="1880" heatid="8921" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.80" />
                    <SPLIT distance="100" swimtime="00:02:21.21" />
                    <SPLIT distance="150" swimtime="00:03:37.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="74" reactiontime="+96" swimtime="00:01:46.73" resultid="1881" heatid="8986" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="67" reactiontime="+106" swimtime="00:02:04.19" resultid="1882" heatid="9009" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="54" reactiontime="+98" swimtime="00:00:57.53" resultid="1883" heatid="9060" lane="6" entrytime="00:00:55.00" />
                <RESULT comment="Z1 - Nieprawidłowa kolejność stylów pływania (motylkowy, grzbietowy, klasyczny, dowolny) (Time: 20:23)" eventid="1578" reactiontime="+116" status="DSQ" swimtime="00:09:47.11" resultid="1884" heatid="9116" lane="3" entrytime="00:10:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.80" />
                    <SPLIT distance="100" swimtime="00:02:24.59" />
                    <SPLIT distance="150" swimtime="00:03:47.34" />
                    <SPLIT distance="200" swimtime="00:05:04.09" />
                    <SPLIT distance="250" swimtime="00:06:25.10" />
                    <SPLIT distance="300" swimtime="00:07:42.61" />
                    <SPLIT distance="350" swimtime="00:08:44.35" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M2 - Wykonanie więcej niż jednego ruchu ramionami pod wodą po starcie lub nawrocie (Time: 9:22)" eventid="1613" reactiontime="+106" status="DSQ" swimtime="00:02:22.53" resultid="1885" heatid="9128" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="42" reactiontime="+114" swimtime="00:05:04.50" resultid="1886" heatid="9144" lane="0" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.73" />
                    <SPLIT distance="100" swimtime="00:02:29.14" />
                    <SPLIT distance="150" swimtime="00:03:47.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-11-14" firstname="Aleksandra" gender="F" lastname="Matraszek" nation="POL" athleteid="1809">
              <RESULTS>
                <RESULT eventid="1062" points="417" reactiontime="+92" swimtime="00:00:31.09" resultid="1810" heatid="8892" lane="8" entrytime="00:00:30.30" />
                <RESULT eventid="1096" points="321" reactiontime="+90" swimtime="00:02:57.97" resultid="1811" heatid="8919" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="150" swimtime="00:02:16.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="386" reactiontime="+89" swimtime="00:01:10.02" resultid="1812" heatid="8983" lane="8" entrytime="00:01:09.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="356" reactiontime="+90" swimtime="00:01:20.00" resultid="1813" heatid="9004" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="365" reactiontime="+92" swimtime="00:01:27.22" resultid="1814" heatid="9042" lane="7" entrytime="00:01:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="320" reactiontime="+95" swimtime="00:02:41.96" resultid="1815" heatid="9092" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:01:58.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="398" reactiontime="+90" swimtime="00:00:39.15" resultid="1816" heatid="9158" lane="7" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-09" firstname="Alina" gender="F" lastname="Wieczorkiewicz" nation="POL" athleteid="1764">
              <RESULTS>
                <RESULT eventid="1062" points="14" reactiontime="+133" swimtime="00:01:34.90" resultid="1793" heatid="8886" lane="0" entrytime="00:01:35.25" />
                <RESULT eventid="1664" points="27" reactiontime="+125" swimtime="00:01:35.42" resultid="1794" heatid="9152" lane="8" entrytime="00:01:35.25" />
                <RESULT eventid="1187" points="23" reactiontime="+94" swimtime="00:01:29.38" resultid="1832" heatid="8948" lane="3" entrytime="00:01:24.35" />
                <RESULT eventid="1290" reactiontime="+129" status="DNF" swimtime="00:00:00.00" resultid="1833" heatid="9001" lane="6" entrytime="00:03:19.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:12.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="26" reactiontime="+121" swimtime="00:03:29.11" resultid="1834" heatid="9037" lane="7" entrytime="00:03:23.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:03:24.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="23" reactiontime="+102" swimtime="00:03:10.93" resultid="1835" heatid="9074" lane="6" entrytime="00:03:00.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="22" reactiontime="+108" swimtime="00:07:00.16" resultid="1836" heatid="9138" lane="7" entrytime="00:06:54.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.44" />
                    <SPLIT distance="100" swimtime="00:03:23.03" />
                    <SPLIT distance="150" swimtime="00:05:13.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-16" firstname="Michalina" gender="F" lastname="Bąk" nation="POL" athleteid="1937">
              <RESULTS>
                <RESULT eventid="1062" points="538" reactiontime="+85" swimtime="00:00:28.57" resultid="1938" heatid="8893" lane="3" entrytime="00:00:27.50" />
                <RESULT eventid="1256" points="537" reactiontime="+86" swimtime="00:01:02.75" resultid="1939" heatid="8984" lane="6" entrytime="00:01:01.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="448" reactiontime="+88" swimtime="00:00:31.84" resultid="1940" heatid="9059" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1595" points="387" reactiontime="+84" swimtime="00:01:14.91" resultid="1941" heatid="9127" lane="8" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-29" firstname="Piotr" gender="M" lastname="Krzekotowski" nation="POL" athleteid="1899">
              <RESULTS>
                <RESULT eventid="1273" points="124" reactiontime="+94" swimtime="00:01:30.05" resultid="1900" heatid="8987" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="96" reactiontime="+94" swimtime="00:01:50.26" resultid="1901" heatid="9009" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="127" reactiontime="+97" swimtime="00:01:50.43" resultid="1902" heatid="9045" lane="9" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="121" reactiontime="+100" swimtime="00:03:20.58" resultid="1903" heatid="9096" lane="1" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:35.44" />
                    <SPLIT distance="150" swimtime="00:02:28.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-11-19" firstname="Judyta" gender="F" lastname="Sołtyk" nation="POL" athleteid="1762">
              <RESULTS>
                <RESULT eventid="1147" points="452" reactiontime="+88" swimtime="00:10:24.49" resultid="1792" heatid="8939" lane="2" entrytime="00:10:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:11.98" />
                    <SPLIT distance="150" swimtime="00:01:50.16" />
                    <SPLIT distance="200" swimtime="00:02:28.99" />
                    <SPLIT distance="250" swimtime="00:03:08.25" />
                    <SPLIT distance="300" swimtime="00:03:47.63" />
                    <SPLIT distance="350" swimtime="00:04:26.87" />
                    <SPLIT distance="400" swimtime="00:05:06.51" />
                    <SPLIT distance="450" swimtime="00:05:46.24" />
                    <SPLIT distance="500" swimtime="00:06:26.05" />
                    <SPLIT distance="550" swimtime="00:07:05.97" />
                    <SPLIT distance="600" swimtime="00:07:46.01" />
                    <SPLIT distance="650" swimtime="00:08:25.93" />
                    <SPLIT distance="700" swimtime="00:09:05.94" />
                    <SPLIT distance="750" swimtime="00:09:45.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-21" firstname="Mateusz" gender="M" lastname="Dudek" nation="POL" athleteid="4163">
              <RESULTS>
                <RESULT eventid="1165" reactiontime="+90" status="DNF" swimtime="00:00:00.00" resultid="4164" heatid="8947" lane="1" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:11.98" />
                    <SPLIT distance="150" swimtime="00:01:50.18" />
                    <SPLIT distance="200" swimtime="00:02:29.08" />
                    <SPLIT distance="250" swimtime="00:03:08.43" />
                    <SPLIT distance="300" swimtime="00:03:47.88" />
                    <SPLIT distance="350" swimtime="00:04:27.81" />
                    <SPLIT distance="400" swimtime="00:05:08.27" />
                    <SPLIT distance="450" swimtime="00:05:48.56" />
                    <SPLIT distance="500" swimtime="00:06:28.61" />
                    <SPLIT distance="550" swimtime="00:07:09.14" />
                    <SPLIT distance="600" swimtime="00:07:50.34" />
                    <SPLIT distance="650" swimtime="00:08:31.44" />
                    <SPLIT distance="700" swimtime="00:09:12.47" />
                    <SPLIT distance="750" swimtime="00:09:54.27" />
                    <SPLIT distance="800" swimtime="00:10:36.14" />
                    <SPLIT distance="850" swimtime="00:11:17.94" />
                    <SPLIT distance="900" swimtime="00:12:00.25" />
                    <SPLIT distance="950" swimtime="00:12:42.05" />
                    <SPLIT distance="1000" swimtime="00:13:24.06" />
                    <SPLIT distance="1050" swimtime="00:14:06.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="484" reactiontime="+79" swimtime="00:02:33.41" resultid="4165" heatid="8978" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:13.65" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="518" reactiontime="+80" swimtime="00:01:09.24" resultid="4166" heatid="9053" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="4167" heatid="9104" lane="2" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" athleteid="2384">
              <RESULTS>
                <RESULT eventid="1165" points="146" reactiontime="+125" swimtime="00:26:51.40" resultid="2385" heatid="8942" lane="0" entrytime="00:28:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:36.00" />
                    <SPLIT distance="150" swimtime="00:02:29.83" />
                    <SPLIT distance="200" swimtime="00:03:23.25" />
                    <SPLIT distance="250" swimtime="00:05:10.95" />
                    <SPLIT distance="350" swimtime="00:07:51.82" />
                    <SPLIT distance="400" swimtime="00:08:45.69" />
                    <SPLIT distance="450" swimtime="00:09:39.80" />
                    <SPLIT distance="500" swimtime="00:10:33.86" />
                    <SPLIT distance="550" swimtime="00:11:28.81" />
                    <SPLIT distance="600" swimtime="00:12:23.24" />
                    <SPLIT distance="650" swimtime="00:13:17.80" />
                    <SPLIT distance="700" swimtime="00:14:12.60" />
                    <SPLIT distance="900" swimtime="00:17:50.65" />
                    <SPLIT distance="950" swimtime="00:18:45.10" />
                    <SPLIT distance="1000" swimtime="00:19:39.72" />
                    <SPLIT distance="1050" swimtime="00:20:33.90" />
                    <SPLIT distance="1100" swimtime="00:21:28.37" />
                    <SPLIT distance="1200" swimtime="00:23:17.61" />
                    <SPLIT distance="1350" swimtime="00:25:07.14" />
                    <SPLIT distance="1400" swimtime="00:26:01.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="143" reactiontime="+113" swimtime="00:01:25.76" resultid="2386" heatid="8987" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="116" reactiontime="+128" swimtime="00:01:53.97" resultid="2387" heatid="9044" lane="5" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="136" reactiontime="+118" swimtime="00:03:12.99" resultid="2388" heatid="9096" lane="7" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.98" />
                    <SPLIT distance="100" swimtime="00:01:33.28" />
                    <SPLIT distance="150" swimtime="00:02:26.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="145" reactiontime="+111" swimtime="00:06:43.31" resultid="2389" heatid="9184" lane="9" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:01:33.90" />
                    <SPLIT distance="150" swimtime="00:02:25.09" />
                    <SPLIT distance="200" swimtime="00:03:17.58" />
                    <SPLIT distance="250" swimtime="00:04:09.87" />
                    <SPLIT distance="350" swimtime="00:05:54.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-10" firstname="Jolanta" gender="F" lastname="Płatek" nation="POL" athleteid="4209">
              <RESULTS>
                <RESULT eventid="1187" points="305" reactiontime="+81" swimtime="00:00:38.12" resultid="4210" heatid="8951" lane="0" entrytime="00:00:39.00" />
                <RESULT eventid="1457" points="301" reactiontime="+77" swimtime="00:01:22.03" resultid="4211" heatid="9076" lane="2" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="287" reactiontime="+76" swimtime="00:03:00.75" resultid="4212" heatid="9140" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                    <SPLIT distance="100" swimtime="00:01:27.15" />
                    <SPLIT distance="150" swimtime="00:02:13.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="274" reactiontime="+98" swimtime="00:06:00.94" resultid="4213" heatid="9180" lane="0" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                    <SPLIT distance="150" swimtime="00:02:09.37" />
                    <SPLIT distance="200" swimtime="00:02:55.07" />
                    <SPLIT distance="250" swimtime="00:03:41.50" />
                    <SPLIT distance="300" swimtime="00:04:28.06" />
                    <SPLIT distance="350" swimtime="00:05:14.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-31" firstname="Piotr" gender="M" lastname="Krogulec" nation="POL" athleteid="5530">
              <RESULTS>
                <RESULT eventid="1079" points="426" reactiontime="+87" swimtime="00:00:26.91" resultid="5531" heatid="8909" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1205" points="377" reactiontime="+67" swimtime="00:00:30.75" resultid="5532" heatid="8962" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1307" points="429" reactiontime="+84" swimtime="00:01:07.16" resultid="5533" heatid="9015" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="421" reactiontime="+82" swimtime="00:00:29.07" resultid="5534" heatid="9069" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1474" points="381" reactiontime="+70" swimtime="00:01:07.46" resultid="5535" heatid="9083" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="382" reactiontime="+86" swimtime="00:01:06.72" resultid="5536" heatid="9135" lane="0" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="367" reactiontime="+77" swimtime="00:00:35.26" resultid="5537" heatid="9169" lane="6" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="2059">
              <RESULTS>
                <RESULT eventid="1079" points="230" reactiontime="+93" swimtime="00:00:33.04" resultid="2060" heatid="8901" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1165" points="163" reactiontime="+106" swimtime="00:25:54.31" resultid="2061" heatid="8942" lane="6" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                    <SPLIT distance="100" swimtime="00:01:29.42" />
                    <SPLIT distance="150" swimtime="00:02:18.73" />
                    <SPLIT distance="200" swimtime="00:03:09.25" />
                    <SPLIT distance="250" swimtime="00:04:00.84" />
                    <SPLIT distance="300" swimtime="00:04:53.99" />
                    <SPLIT distance="350" swimtime="00:05:44.84" />
                    <SPLIT distance="400" swimtime="00:06:39.22" />
                    <SPLIT distance="450" swimtime="00:07:31.47" />
                    <SPLIT distance="500" swimtime="00:08:22.86" />
                    <SPLIT distance="550" swimtime="00:09:14.35" />
                    <SPLIT distance="600" swimtime="00:10:06.62" />
                    <SPLIT distance="650" swimtime="00:10:59.50" />
                    <SPLIT distance="700" swimtime="00:11:52.04" />
                    <SPLIT distance="750" swimtime="00:12:44.47" />
                    <SPLIT distance="800" swimtime="00:13:38.30" />
                    <SPLIT distance="850" swimtime="00:14:30.39" />
                    <SPLIT distance="900" swimtime="00:15:23.74" />
                    <SPLIT distance="950" swimtime="00:16:14.68" />
                    <SPLIT distance="1000" swimtime="00:17:08.56" />
                    <SPLIT distance="1050" swimtime="00:17:59.16" />
                    <SPLIT distance="1100" swimtime="00:18:54.66" />
                    <SPLIT distance="1150" swimtime="00:19:46.58" />
                    <SPLIT distance="1200" swimtime="00:20:39.06" />
                    <SPLIT distance="1250" swimtime="00:21:33.38" />
                    <SPLIT distance="1300" swimtime="00:22:25.07" />
                    <SPLIT distance="1350" swimtime="00:23:17.71" />
                    <SPLIT distance="1400" swimtime="00:24:10.49" />
                    <SPLIT distance="1450" swimtime="00:25:05.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="166" reactiontime="+80" swimtime="00:00:40.40" resultid="2062" heatid="8958" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1341" points="84" reactiontime="+98" swimtime="00:04:07.70" resultid="2063" heatid="9026" lane="6" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                    <SPLIT distance="100" swimtime="00:01:55.07" />
                    <SPLIT distance="150" swimtime="00:03:02.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="163" reactiontime="+81" swimtime="00:01:29.49" resultid="2064" heatid="9081" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="182" reactiontime="+96" swimtime="00:02:55.28" resultid="2065" heatid="9098" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:23.59" />
                    <SPLIT distance="150" swimtime="00:02:10.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="124" reactiontime="+97" swimtime="00:01:37.07" resultid="2066" heatid="9130" lane="9" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="155" reactiontime="+99" swimtime="00:06:34.51" resultid="2067" heatid="9185" lane="5" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                    <SPLIT distance="100" swimtime="00:01:27.31" />
                    <SPLIT distance="150" swimtime="00:02:18.34" />
                    <SPLIT distance="200" swimtime="00:03:09.45" />
                    <SPLIT distance="250" swimtime="00:04:02.46" />
                    <SPLIT distance="300" swimtime="00:04:52.61" />
                    <SPLIT distance="350" swimtime="00:05:45.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-01" firstname="Jolanta" gender="F" lastname="Zawadzka" nation="POL" athleteid="2390">
              <RESULTS>
                <RESULT eventid="1290" points="202" reactiontime="+100" swimtime="00:01:36.57" resultid="2391" heatid="9003" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="185" reactiontime="+84" swimtime="00:00:42.77" resultid="2392" heatid="9056" lane="9" entrytime="00:00:43.00" />
                <RESULT eventid="1664" points="236" reactiontime="+92" swimtime="00:00:46.57" resultid="2393" heatid="9155" lane="6" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-12-07" firstname="Ewelina" gender="F" lastname="Kot" nation="POL" athleteid="5617">
              <RESULTS>
                <RESULT eventid="1096" points="281" reactiontime="+91" swimtime="00:03:06.03" resultid="5618" heatid="8918" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:25.81" />
                    <SPLIT distance="150" swimtime="00:02:22.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="268" reactiontime="+95" swimtime="00:12:22.80" resultid="5619" heatid="8938" lane="1" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:25.29" />
                    <SPLIT distance="150" swimtime="00:02:10.58" />
                    <SPLIT distance="200" swimtime="00:02:56.68" />
                    <SPLIT distance="250" swimtime="00:03:43.46" />
                    <SPLIT distance="300" swimtime="00:04:30.19" />
                    <SPLIT distance="350" swimtime="00:05:17.18" />
                    <SPLIT distance="400" swimtime="00:06:04.54" />
                    <SPLIT distance="450" swimtime="00:06:51.75" />
                    <SPLIT distance="500" swimtime="00:07:39.15" />
                    <SPLIT distance="550" swimtime="00:08:26.64" />
                    <SPLIT distance="600" swimtime="00:09:14.37" />
                    <SPLIT distance="650" swimtime="00:10:01.86" />
                    <SPLIT distance="700" swimtime="00:10:49.57" />
                    <SPLIT distance="750" swimtime="00:11:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="5620" heatid="9180" lane="7" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-02" firstname="Bernard" gender="M" lastname="Wierzbik" nation="POL" athleteid="6176">
              <RESULTS>
                <RESULT eventid="1307" points="224" reactiontime="+85" swimtime="00:01:23.37" resultid="6177" heatid="9012" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="170" reactiontime="+106" swimtime="00:03:15.73" resultid="6178" heatid="9028" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="100" swimtime="00:01:29.76" />
                    <SPLIT distance="150" swimtime="00:02:23.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="249" reactiontime="+85" swimtime="00:00:34.64" resultid="6179" heatid="9065" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1613" points="220" reactiontime="+93" swimtime="00:01:20.21" resultid="6180" heatid="9132" lane="7" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-03" firstname="Patryk" gender="M" lastname="Dzwonek" nation="POL" athleteid="6332">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="6333" heatid="8895" lane="0" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="6334" heatid="8954" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-06-28" firstname="Bolesław" gender="M" lastname="Czyż" nation="POL" athleteid="6173" />
            <ATHLETE birthdate="1994-09-27" firstname="Aleksandra" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="6340">
              <RESULTS>
                <RESULT eventid="1187" points="480" reactiontime="+63" swimtime="00:00:32.77" resultid="6341" heatid="8953" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1256" points="465" reactiontime="+75" swimtime="00:01:05.80" resultid="6342" heatid="8983" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="412" reactiontime="+73" swimtime="00:01:13.93" resultid="6343" heatid="9078" lane="1" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-04-23" firstname="Marek" gender="M" lastname="Pisulak" nation="POL" athleteid="2041">
              <RESULTS>
                <RESULT eventid="1079" points="72" reactiontime="+103" swimtime="00:00:48.50" resultid="2042" heatid="8896" lane="4" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-30" firstname="Patryk" gender="M" lastname="Suchodolski" nation="POL" athleteid="6335">
              <RESULTS>
                <RESULT eventid="1205" points="403" reactiontime="+68" swimtime="00:00:30.08" resultid="6336" heatid="8964" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1239" points="397" reactiontime="+82" swimtime="00:02:43.80" resultid="6337" heatid="8978" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:01:58.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="486" reactiontime="+77" swimtime="00:01:10.72" resultid="6338" heatid="9053" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="438" reactiontime="+73" swimtime="00:00:28.69" resultid="6339" heatid="9072" lane="9" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Michał" gender="M" lastname="Gawroński" nation="POL" athleteid="4168">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="4169" heatid="8929" lane="4" entrytime="00:02:30.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="4170" heatid="8963" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="4171" heatid="8977" lane="6" entrytime="00:02:50.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="4172" heatid="9104" lane="0" entrytime="00:02:12.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="4173" heatid="9122" lane="2" entrytime="00:05:15.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="4174" heatid="9149" lane="5" entrytime="00:02:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-03" firstname="Ilona" gender="F" lastname="Szkudlarz" nation="POL" athleteid="4203">
              <RESULTS>
                <RESULT eventid="1187" points="214" reactiontime="+79" swimtime="00:00:42.87" resultid="4204" heatid="8950" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1290" points="257" reactiontime="+92" swimtime="00:01:29.12" resultid="4205" heatid="9002" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="259" reactiontime="+96" swimtime="00:01:37.79" resultid="4206" heatid="9039" lane="3" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="273" reactiontime="+94" swimtime="00:02:50.67" resultid="4207" heatid="9091" lane="0" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:22.79" />
                    <SPLIT distance="150" swimtime="00:02:06.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="267" reactiontime="+93" swimtime="00:00:44.71" resultid="4208" heatid="9155" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-11-29" firstname="Edward" gender="M" lastname="Dziekoński" nation="POL" athleteid="3360">
              <RESULTS>
                <RESULT eventid="1079" points="137" reactiontime="+109" swimtime="00:00:39.26" resultid="3361" heatid="8897" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1165" points="122" reactiontime="+130" swimtime="00:28:31.33" resultid="3362" heatid="8942" lane="8" entrytime="00:28:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.34" />
                    <SPLIT distance="100" swimtime="00:01:45.53" />
                    <SPLIT distance="150" swimtime="00:02:42.95" />
                    <SPLIT distance="200" swimtime="00:03:40.64" />
                    <SPLIT distance="250" swimtime="00:04:37.25" />
                    <SPLIT distance="300" swimtime="00:05:34.65" />
                    <SPLIT distance="350" swimtime="00:06:33.12" />
                    <SPLIT distance="400" swimtime="00:07:31.15" />
                    <SPLIT distance="450" swimtime="00:08:28.68" />
                    <SPLIT distance="500" swimtime="00:09:25.11" />
                    <SPLIT distance="550" swimtime="00:10:21.28" />
                    <SPLIT distance="600" swimtime="00:11:17.45" />
                    <SPLIT distance="650" swimtime="00:12:14.69" />
                    <SPLIT distance="700" swimtime="00:13:11.95" />
                    <SPLIT distance="750" swimtime="00:14:09.87" />
                    <SPLIT distance="800" swimtime="00:15:07.02" />
                    <SPLIT distance="850" swimtime="00:16:04.31" />
                    <SPLIT distance="900" swimtime="00:17:02.73" />
                    <SPLIT distance="950" swimtime="00:17:59.96" />
                    <SPLIT distance="1000" swimtime="00:18:57.23" />
                    <SPLIT distance="1050" swimtime="00:19:54.91" />
                    <SPLIT distance="1100" swimtime="00:20:52.39" />
                    <SPLIT distance="1150" swimtime="00:21:49.85" />
                    <SPLIT distance="1200" swimtime="00:22:48.22" />
                    <SPLIT distance="1250" swimtime="00:23:47.10" />
                    <SPLIT distance="1300" swimtime="00:24:45.51" />
                    <SPLIT distance="1350" swimtime="00:25:43.81" />
                    <SPLIT distance="1400" swimtime="00:26:40.97" />
                    <SPLIT distance="1450" swimtime="00:27:38.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="84" reactiontime="+99" swimtime="00:00:50.66" resultid="3363" heatid="8956" lane="3" entrytime="00:00:48.00" />
                <RESULT eventid="1307" points="102" reactiontime="+104" swimtime="00:01:48.27" resultid="3364" heatid="9009" lane="5" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="126" reactiontime="+106" swimtime="00:00:43.41" resultid="3365" heatid="9062" lane="0" entrytime="00:00:41.50" />
                <RESULT eventid="1508" points="106" reactiontime="+110" swimtime="00:03:29.57" resultid="3366" heatid="9096" lane="3" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:36.98" />
                    <SPLIT distance="150" swimtime="00:02:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="69" reactiontime="+126" swimtime="00:04:17.73" resultid="3367" heatid="9144" lane="3" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.47" />
                    <SPLIT distance="100" swimtime="00:02:03.62" />
                    <SPLIT distance="150" swimtime="00:03:11.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="111" reactiontime="+126" swimtime="00:07:21.58" resultid="3368" heatid="9183" lane="4" entrytime="00:07:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.20" />
                    <SPLIT distance="100" swimtime="00:01:38.62" />
                    <SPLIT distance="150" swimtime="00:02:33.79" />
                    <SPLIT distance="200" swimtime="00:03:32.23" />
                    <SPLIT distance="250" swimtime="00:04:31.25" />
                    <SPLIT distance="300" swimtime="00:05:29.81" />
                    <SPLIT distance="350" swimtime="00:06:27.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-24" firstname="Igor" gender="M" lastname="Okarmus" nation="POL" athleteid="2038">
              <RESULTS>
                <RESULT eventid="1165" points="332" reactiontime="+106" swimtime="00:20:26.98" resultid="2039" heatid="8947" lane="9" entrytime="00:20:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:14.34" />
                    <SPLIT distance="150" swimtime="00:01:53.58" />
                    <SPLIT distance="200" swimtime="00:02:33.41" />
                    <SPLIT distance="250" swimtime="00:03:13.21" />
                    <SPLIT distance="300" swimtime="00:03:54.04" />
                    <SPLIT distance="350" swimtime="00:04:34.56" />
                    <SPLIT distance="400" swimtime="00:05:15.32" />
                    <SPLIT distance="450" swimtime="00:05:56.08" />
                    <SPLIT distance="500" swimtime="00:06:37.00" />
                    <SPLIT distance="550" swimtime="00:07:17.49" />
                    <SPLIT distance="600" swimtime="00:07:58.33" />
                    <SPLIT distance="650" swimtime="00:08:39.30" />
                    <SPLIT distance="700" swimtime="00:09:20.68" />
                    <SPLIT distance="750" swimtime="00:10:02.16" />
                    <SPLIT distance="800" swimtime="00:10:43.31" />
                    <SPLIT distance="850" swimtime="00:11:24.18" />
                    <SPLIT distance="900" swimtime="00:12:06.41" />
                    <SPLIT distance="950" swimtime="00:12:47.74" />
                    <SPLIT distance="1000" swimtime="00:13:29.03" />
                    <SPLIT distance="1050" swimtime="00:14:11.06" />
                    <SPLIT distance="1100" swimtime="00:14:52.96" />
                    <SPLIT distance="1150" swimtime="00:15:34.56" />
                    <SPLIT distance="1200" swimtime="00:16:17.09" />
                    <SPLIT distance="1250" swimtime="00:16:58.91" />
                    <SPLIT distance="1300" swimtime="00:17:41.94" />
                    <SPLIT distance="1350" swimtime="00:18:22.95" />
                    <SPLIT distance="1400" swimtime="00:19:05.04" />
                    <SPLIT distance="1450" swimtime="00:19:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="2040" heatid="9013" lane="7" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-12-02" firstname="Krzysztof" gender="M" lastname="Drózd" nation="POL" athleteid="6344">
              <RESULTS>
                <RESULT eventid="1205" points="318" reactiontime="+64" swimtime="00:00:32.55" resultid="6345" heatid="8959" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1307" points="320" reactiontime="+64" swimtime="00:01:14.04" resultid="6346" heatid="9015" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="276" reactiontime="+72" swimtime="00:01:15.16" resultid="6347" heatid="9083" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 18:57)" eventid="1508" reactiontime="+54" status="DSQ" swimtime="00:02:27.99" resultid="6348" heatid="9100" lane="0" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                    <SPLIT distance="150" swimtime="00:01:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="258" reactiontime="+69" swimtime="00:02:46.63" resultid="6349" heatid="9148" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:01:21.18" />
                    <SPLIT distance="150" swimtime="00:02:05.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-19" firstname="Michał" gender="M" lastname="Łączny" nation="POL" athleteid="3369">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="3370" heatid="8909" lane="5" entrytime="00:00:27.85" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3371" heatid="8994" lane="9" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-08-01" firstname="Mieczysław" gender="M" lastname="Putek" nation="POL" athleteid="3127">
              <RESULTS>
                <RESULT eventid="1205" points="12" reactiontime="+103" swimtime="00:01:36.19" resultid="3128" heatid="8954" lane="3" />
                <RESULT eventid="1273" points="25" reactiontime="+131" swimtime="00:02:31.87" resultid="3129" heatid="8986" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-18" firstname="Kazimierz" gender="M" lastname="Sinicki" nation="POL" athleteid="1887">
              <RESULTS>
                <RESULT eventid="1079" points="332" reactiontime="+82" swimtime="00:00:29.24" resultid="1888" heatid="8905" lane="5" entrytime="00:00:29.95" />
                <RESULT eventid="1273" points="295" reactiontime="+88" swimtime="00:01:07.44" resultid="1889" heatid="8991" lane="4" entrytime="00:01:08.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="245" reactiontime="+92" swimtime="00:00:34.83" resultid="1890" heatid="9063" lane="4" entrytime="00:00:35.75" />
                <RESULT eventid="1508" points="246" reactiontime="+97" swimtime="00:02:38.54" resultid="1891" heatid="9099" lane="2" entrytime="00:02:37.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                    <SPLIT distance="150" swimtime="00:01:56.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-07-07" firstname="Ryszard" gender="M" lastname="Tatarczuk" nation="POL" athleteid="3372">
              <RESULTS>
                <RESULT eventid="1508" points="184" reactiontime="+109" swimtime="00:02:54.41" resultid="3373" heatid="9097" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:20.40" />
                    <SPLIT distance="150" swimtime="00:02:06.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="181" reactiontime="+100" swimtime="00:06:15.22" resultid="3374" heatid="9185" lane="3" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:25.41" />
                    <SPLIT distance="150" swimtime="00:02:11.92" />
                    <SPLIT distance="200" swimtime="00:02:59.18" />
                    <SPLIT distance="250" swimtime="00:03:48.14" />
                    <SPLIT distance="300" swimtime="00:04:37.72" />
                    <SPLIT distance="350" swimtime="00:05:28.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-22" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="9193">
              <RESULTS>
                <RESULT eventid="1165" points="144" reactiontime="+114" swimtime="00:26:59.72" resultid="9194" heatid="8940" lane="8" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:01:30.43" />
                    <SPLIT distance="150" swimtime="00:02:22.28" />
                    <SPLIT distance="200" swimtime="00:03:15.54" />
                    <SPLIT distance="250" swimtime="00:04:09.91" />
                    <SPLIT distance="300" swimtime="00:06:00.52" />
                    <SPLIT distance="350" swimtime="00:06:56.25" />
                    <SPLIT distance="400" swimtime="00:07:52.35" />
                    <SPLIT distance="450" swimtime="00:08:47.27" />
                    <SPLIT distance="500" swimtime="00:09:43.43" />
                    <SPLIT distance="550" swimtime="00:10:39.13" />
                    <SPLIT distance="600" swimtime="00:11:33.53" />
                    <SPLIT distance="650" swimtime="00:12:28.98" />
                    <SPLIT distance="700" swimtime="00:13:24.39" />
                    <SPLIT distance="750" swimtime="00:14:20.91" />
                    <SPLIT distance="800" swimtime="00:15:15.47" />
                    <SPLIT distance="850" swimtime="00:16:11.03" />
                    <SPLIT distance="900" swimtime="00:17:05.37" />
                    <SPLIT distance="950" swimtime="00:18:00.35" />
                    <SPLIT distance="1000" swimtime="00:18:55.09" />
                    <SPLIT distance="1050" swimtime="00:19:50.80" />
                    <SPLIT distance="1100" swimtime="00:20:46.14" />
                    <SPLIT distance="1150" swimtime="00:21:41.71" />
                    <SPLIT distance="1200" swimtime="00:22:36.28" />
                    <SPLIT distance="1250" swimtime="00:23:30.20" />
                    <SPLIT distance="1300" swimtime="00:24:24.94" />
                    <SPLIT distance="1350" swimtime="00:25:18.93" />
                    <SPLIT distance="1400" swimtime="00:26:12.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="157" reactiontime="+98" swimtime="00:00:37.49" resultid="9195" heatid="8894" lane="8" late="yes" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="9196" heatid="9094" lane="9" late="yes" />
                <RESULT eventid="1744" points="147" reactiontime="+106" swimtime="00:06:42.08" resultid="9197" heatid="9182" lane="9" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:01:29.25" />
                    <SPLIT distance="150" swimtime="00:02:21.60" />
                    <SPLIT distance="200" swimtime="00:03:14.89" />
                    <SPLIT distance="250" swimtime="00:04:08.41" />
                    <SPLIT distance="300" swimtime="00:05:01.02" />
                    <SPLIT distance="350" swimtime="00:05:53.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-14" firstname="Mateusz" gender="M" lastname="Kwaśniewski" nation="POL" athleteid="6326">
              <RESULTS>
                <RESULT eventid="1273" points="567" reactiontime="+71" swimtime="00:00:54.28" resultid="6327" heatid="9000" lane="1" entrytime="00:00:55.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="553" reactiontime="+68" swimtime="00:00:26.55" resultid="6328" heatid="9072" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1508" points="511" reactiontime="+70" swimtime="00:02:04.29" resultid="6329" heatid="9106" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.84" />
                    <SPLIT distance="100" swimtime="00:00:59.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="494" reactiontime="+72" swimtime="00:01:01.25" resultid="6330" heatid="9136" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="6331" heatid="9192" lane="7" entrytime="00:04:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-10" firstname="Jarosław" gender="M" lastname="Wnęk" nation="POL" athleteid="4156">
              <RESULTS>
                <RESULT eventid="1165" points="387" reactiontime="+94" swimtime="00:19:25.78" resultid="4157" heatid="8946" lane="6" entrytime="00:20:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:12.71" />
                    <SPLIT distance="150" swimtime="00:01:50.97" />
                    <SPLIT distance="200" swimtime="00:02:29.77" />
                    <SPLIT distance="250" swimtime="00:03:08.85" />
                    <SPLIT distance="300" swimtime="00:03:47.94" />
                    <SPLIT distance="350" swimtime="00:04:27.43" />
                    <SPLIT distance="400" swimtime="00:05:06.27" />
                    <SPLIT distance="450" swimtime="00:05:45.81" />
                    <SPLIT distance="500" swimtime="00:06:24.66" />
                    <SPLIT distance="550" swimtime="00:07:04.63" />
                    <SPLIT distance="600" swimtime="00:07:43.07" />
                    <SPLIT distance="650" swimtime="00:08:22.31" />
                    <SPLIT distance="700" swimtime="00:09:01.16" />
                    <SPLIT distance="750" swimtime="00:09:40.73" />
                    <SPLIT distance="800" swimtime="00:10:19.96" />
                    <SPLIT distance="850" swimtime="00:10:59.52" />
                    <SPLIT distance="900" swimtime="00:11:38.76" />
                    <SPLIT distance="950" swimtime="00:12:18.28" />
                    <SPLIT distance="1000" swimtime="00:12:57.75" />
                    <SPLIT distance="1050" swimtime="00:13:36.67" />
                    <SPLIT distance="1100" swimtime="00:14:16.14" />
                    <SPLIT distance="1150" swimtime="00:14:55.95" />
                    <SPLIT distance="1200" swimtime="00:15:34.95" />
                    <SPLIT distance="1250" swimtime="00:16:13.23" />
                    <SPLIT distance="1300" swimtime="00:16:53.46" />
                    <SPLIT distance="1350" swimtime="00:17:31.77" />
                    <SPLIT distance="1400" swimtime="00:18:11.10" />
                    <SPLIT distance="1450" swimtime="00:18:49.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="406" reactiontime="+86" swimtime="00:01:00.69" resultid="4158" heatid="8996" lane="3" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="287" reactiontime="+91" swimtime="00:02:44.56" resultid="4159" heatid="9029" lane="1" entrytime="00:02:45.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:02:01.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="404" reactiontime="+86" swimtime="00:02:14.41" resultid="4160" heatid="9103" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:04.72" />
                    <SPLIT distance="150" swimtime="00:01:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="4161" heatid="9121" lane="7" entrytime="00:05:40.00" />
                <RESULT eventid="1744" points="392" reactiontime="+93" swimtime="00:04:49.77" resultid="4162" heatid="9190" lane="4" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:08.62" />
                    <SPLIT distance="150" swimtime="00:01:45.77" />
                    <SPLIT distance="200" swimtime="00:02:23.56" />
                    <SPLIT distance="250" swimtime="00:03:00.66" />
                    <SPLIT distance="300" swimtime="00:03:37.88" />
                    <SPLIT distance="350" swimtime="00:04:15.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-07" firstname="Krzysztof" gender="M" lastname="Nowak" nation="POL" athleteid="4195" />
            <ATHLETE birthdate="1980-01-13" firstname="Michał" gender="M" lastname="Sroka" nation="POL" athleteid="2394">
              <RESULTS>
                <RESULT eventid="1079" points="258" reactiontime="+92" swimtime="00:00:31.82" resultid="2395" heatid="8900" lane="4" entrytime="00:00:32.69" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="2396" heatid="8923" lane="3" entrytime="00:03:30.00" />
                <RESULT eventid="1273" points="229" reactiontime="+81" swimtime="00:01:13.45" resultid="2397" heatid="8990" lane="1" entrytime="00:01:12.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="193" reactiontime="+97" swimtime="00:01:27.58" resultid="2398" heatid="9011" lane="2" entrytime="00:01:28.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="152" reactiontime="+90" swimtime="00:00:40.77" resultid="2399" heatid="9062" lane="8" entrytime="00:00:41.11" />
                <RESULT eventid="1508" points="181" reactiontime="+96" swimtime="00:02:55.43" resultid="2400" heatid="9096" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:21.38" />
                    <SPLIT distance="150" swimtime="00:02:10.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="119" reactiontime="+97" swimtime="00:01:38.37" resultid="2401" heatid="9130" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="163" reactiontime="+100" swimtime="00:06:28.38" resultid="2402" heatid="9184" lane="2" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:30.59" />
                    <SPLIT distance="150" swimtime="00:02:23.95" />
                    <SPLIT distance="200" swimtime="00:03:14.64" />
                    <SPLIT distance="250" swimtime="00:04:05.51" />
                    <SPLIT distance="300" swimtime="00:04:57.64" />
                    <SPLIT distance="350" swimtime="00:05:49.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-16" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="2043">
              <RESULTS>
                <RESULT eventid="1079" points="392" reactiontime="+81" swimtime="00:00:27.66" resultid="2044" heatid="8909" lane="7" entrytime="00:00:27.95" />
                <RESULT eventid="1113" points="352" reactiontime="+84" swimtime="00:02:35.17" resultid="2045" heatid="8928" lane="3" entrytime="00:02:38.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:58.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="381" reactiontime="+83" swimtime="00:01:01.94" resultid="2046" heatid="8995" lane="4" entrytime="00:01:01.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="358" reactiontime="+84" swimtime="00:01:11.29" resultid="2047" heatid="9017" lane="7" entrytime="00:01:10.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="381" reactiontime="+84" swimtime="00:00:30.07" resultid="2048" heatid="9068" lane="1" entrytime="00:00:30.55" />
                <RESULT eventid="1613" points="343" reactiontime="+86" swimtime="00:01:09.14" resultid="2049" heatid="9134" lane="8" entrytime="00:01:09.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="275" reactiontime="+74" swimtime="00:02:43.16" resultid="2050" heatid="9147" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="150" swimtime="00:02:01.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-06-06" firstname="Jolanta" gender="F" lastname="Lipińska" nation="POL" athleteid="1817">
              <RESULTS>
                <RESULT eventid="1096" points="27" reactiontime="+119" swimtime="00:06:42.67" resultid="1818" heatid="8916" lane="6" entrytime="00:06:26.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.94" />
                    <SPLIT distance="100" swimtime="00:03:29.25" />
                    <SPLIT distance="150" swimtime="00:05:16.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="60" reactiontime="+134" swimtime="00:05:42.70" resultid="1819" heatid="8967" lane="0" entrytime="00:05:51.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.26" />
                    <SPLIT distance="100" swimtime="00:02:49.15" />
                    <SPLIT distance="150" swimtime="00:04:19.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="28" reactiontime="+118" swimtime="00:03:05.09" resultid="1820" heatid="9001" lane="3" entrytime="00:02:57.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="51" reactiontime="+113" swimtime="00:02:48.06" resultid="1821" heatid="9037" lane="6" entrytime="00:02:50.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="30" reactiontime="+83" swimtime="00:02:56.78" resultid="1822" heatid="9074" lane="3" entrytime="00:02:53.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="31" reactiontime="+75" swimtime="00:06:18.21" resultid="1823" heatid="9138" lane="6" entrytime="00:05:58.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.85" />
                    <SPLIT distance="100" swimtime="00:03:00.58" />
                    <SPLIT distance="150" swimtime="00:04:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="36" reactiontime="+108" swimtime="00:11:43.81" resultid="1824" heatid="9177" lane="3" entrytime="00:11:36.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.15" />
                    <SPLIT distance="100" swimtime="00:02:49.17" />
                    <SPLIT distance="150" swimtime="00:04:18.92" />
                    <SPLIT distance="200" swimtime="00:05:48.11" />
                    <SPLIT distance="250" swimtime="00:07:17.57" />
                    <SPLIT distance="300" swimtime="00:08:48.20" />
                    <SPLIT distance="350" swimtime="00:10:18.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-08-10" firstname="Robert" gender="M" lastname="Sowa" nation="POL" athleteid="4214">
              <RESULTS>
                <RESULT eventid="1113" points="438" reactiontime="+92" swimtime="00:02:24.34" resultid="4215" heatid="8929" lane="0" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                    <SPLIT distance="150" swimtime="00:01:49.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="395" reactiontime="+67" swimtime="00:00:30.26" resultid="4216" heatid="8962" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1307" points="446" reactiontime="+84" swimtime="00:01:06.26" resultid="4217" heatid="9018" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="448" reactiontime="+62" swimtime="00:01:03.93" resultid="4218" heatid="9086" lane="8" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="4219" heatid="9102" lane="6" entrytime="00:02:18.00" />
                <RESULT eventid="1647" points="432" reactiontime="+66" swimtime="00:02:20.26" resultid="4220" heatid="9148" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:44.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="411" reactiontime="+97" swimtime="00:04:45.29" resultid="4221" heatid="9191" lane="0" entrytime="00:04:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="100" swimtime="00:01:09.10" />
                    <SPLIT distance="150" swimtime="00:01:46.36" />
                    <SPLIT distance="200" swimtime="00:02:23.72" />
                    <SPLIT distance="250" swimtime="00:03:00.67" />
                    <SPLIT distance="300" swimtime="00:03:36.76" />
                    <SPLIT distance="350" swimtime="00:04:12.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-09-08" firstname="Igor" gender="M" lastname="Zalewski" nation="POL" athleteid="1800">
              <RESULTS>
                <RESULT eventid="1113" points="407" reactiontime="+72" swimtime="00:02:27.93" resultid="1801" heatid="8929" lane="3" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:07.82" />
                    <SPLIT distance="150" swimtime="00:01:53.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="386" reactiontime="+81" swimtime="00:19:27.54" resultid="1802" heatid="8947" lane="0" entrytime="00:20:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                    <SPLIT distance="150" swimtime="00:01:50.14" />
                    <SPLIT distance="200" swimtime="00:02:28.81" />
                    <SPLIT distance="250" swimtime="00:03:07.90" />
                    <SPLIT distance="300" swimtime="00:03:47.05" />
                    <SPLIT distance="350" swimtime="00:04:26.15" />
                    <SPLIT distance="400" swimtime="00:05:05.46" />
                    <SPLIT distance="450" swimtime="00:05:45.02" />
                    <SPLIT distance="500" swimtime="00:06:24.43" />
                    <SPLIT distance="550" swimtime="00:07:03.78" />
                    <SPLIT distance="600" swimtime="00:07:43.00" />
                    <SPLIT distance="650" swimtime="00:08:22.69" />
                    <SPLIT distance="700" swimtime="00:09:02.15" />
                    <SPLIT distance="750" swimtime="00:09:41.55" />
                    <SPLIT distance="800" swimtime="00:10:21.22" />
                    <SPLIT distance="850" swimtime="00:11:00.66" />
                    <SPLIT distance="900" swimtime="00:11:39.48" />
                    <SPLIT distance="950" swimtime="00:12:18.57" />
                    <SPLIT distance="1000" swimtime="00:12:57.82" />
                    <SPLIT distance="1050" swimtime="00:13:37.07" />
                    <SPLIT distance="1100" swimtime="00:14:16.29" />
                    <SPLIT distance="1150" swimtime="00:14:55.63" />
                    <SPLIT distance="1200" swimtime="00:15:34.85" />
                    <SPLIT distance="1250" swimtime="00:16:14.26" />
                    <SPLIT distance="1300" swimtime="00:16:53.57" />
                    <SPLIT distance="1350" swimtime="00:17:32.87" />
                    <SPLIT distance="1400" swimtime="00:18:12.56" />
                    <SPLIT distance="1450" swimtime="00:18:51.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="434" reactiontime="+73" swimtime="00:01:06.89" resultid="1803" heatid="9018" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="366" reactiontime="+78" swimtime="00:02:31.69" resultid="1804" heatid="9029" lane="5" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:52.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="424" reactiontime="+73" swimtime="00:02:12.22" resultid="1805" heatid="9101" lane="5" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                    <SPLIT distance="100" swimtime="00:01:01.77" />
                    <SPLIT distance="150" swimtime="00:01:37.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="406" reactiontime="+75" swimtime="00:05:17.96" resultid="1806" heatid="9121" lane="4" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:10.18" />
                    <SPLIT distance="150" swimtime="00:01:51.39" />
                    <SPLIT distance="200" swimtime="00:02:31.93" />
                    <SPLIT distance="250" swimtime="00:03:18.44" />
                    <SPLIT distance="300" swimtime="00:04:05.11" />
                    <SPLIT distance="350" swimtime="00:04:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="438" reactiontime="+77" swimtime="00:01:03.78" resultid="1807" heatid="9134" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="386" reactiontime="+79" swimtime="00:04:51.44" resultid="1808" heatid="9190" lane="0" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:08.69" />
                    <SPLIT distance="150" swimtime="00:01:45.61" />
                    <SPLIT distance="200" swimtime="00:02:22.92" />
                    <SPLIT distance="250" swimtime="00:03:00.77" />
                    <SPLIT distance="300" swimtime="00:03:38.64" />
                    <SPLIT distance="350" swimtime="00:04:16.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-06-26" firstname="Kazimierz" gender="M" lastname="Ślizowski" nation="POL" athleteid="3130">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="3131" heatid="8954" lane="9" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3132" heatid="8985" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-03-06" firstname="Andrzej" gender="M" lastname="Pawlak" nation="POL" athleteid="1904">
              <RESULTS>
                <RESULT eventid="1079" points="193" reactiontime="+120" swimtime="00:00:35.00" resultid="1905" heatid="8900" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1113" points="160" reactiontime="+111" swimtime="00:03:21.87" resultid="1906" heatid="8924" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                    <SPLIT distance="100" swimtime="00:01:36.59" />
                    <SPLIT distance="150" swimtime="00:02:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="174" reactiontime="+76" swimtime="00:00:39.79" resultid="1907" heatid="8957" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1307" points="192" reactiontime="+112" swimtime="00:01:27.81" resultid="1908" heatid="9012" lane="0" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="1909" heatid="9163" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="1910" heatid="9185" lane="8" entrytime="00:06:22.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-12-14" firstname="Jakub" gender="M" lastname="Gorycki" nation="POL" athleteid="5076">
              <RESULTS>
                <RESULT eventid="1113" points="292" reactiontime="+82" swimtime="00:02:45.17" resultid="5077" heatid="8928" lane="6" entrytime="00:02:39.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:15.51" />
                    <SPLIT distance="150" swimtime="00:02:05.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="5078" heatid="8947" lane="2" entrytime="00:19:45.00" />
                <RESULT eventid="1273" points="357" reactiontime="+85" swimtime="00:01:03.31" resultid="5079" heatid="8996" lane="0" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="5080" heatid="9017" lane="2" entrytime="00:01:10.12" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="5081" heatid="9068" lane="5" entrytime="00:00:30.10" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="5082" heatid="9102" lane="0" entrytime="00:02:20.16" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="5083" heatid="9134" lane="1" entrytime="00:01:09.15" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="5084" heatid="9189" lane="4" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-04-13" firstname="Jadwiga" gender="F" lastname="Kowalik" nation="POL" athleteid="5085">
              <RESULTS>
                <RESULT eventid="1062" points="14" swimtime="00:01:36.30" resultid="5086" heatid="8886" lane="8" entrytime="00:00:59.00" />
                <RESULT eventid="1187" points="15" reactiontime="+99" swimtime="00:01:42.65" resultid="5087" heatid="8948" lane="4" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-09-19" firstname="Zygmunt" gender="M" lastname="Lewandowski" nation="POL" athleteid="7224">
              <RESULTS>
                <RESULT eventid="1165" points="107" reactiontime="+111" swimtime="00:29:46.39" resultid="7225" heatid="8941" lane="1" entrytime="00:33:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                    <SPLIT distance="100" swimtime="00:01:46.19" />
                    <SPLIT distance="150" swimtime="00:02:43.15" />
                    <SPLIT distance="200" swimtime="00:03:41.25" />
                    <SPLIT distance="250" swimtime="00:04:39.43" />
                    <SPLIT distance="300" swimtime="00:05:36.88" />
                    <SPLIT distance="350" swimtime="00:06:35.53" />
                    <SPLIT distance="400" swimtime="00:07:34.60" />
                    <SPLIT distance="450" swimtime="00:08:33.93" />
                    <SPLIT distance="500" swimtime="00:09:33.61" />
                    <SPLIT distance="550" swimtime="00:10:33.34" />
                    <SPLIT distance="600" swimtime="00:11:33.51" />
                    <SPLIT distance="650" swimtime="00:12:33.97" />
                    <SPLIT distance="700" swimtime="00:13:33.97" />
                    <SPLIT distance="750" swimtime="00:14:34.32" />
                    <SPLIT distance="800" swimtime="00:15:34.58" />
                    <SPLIT distance="850" swimtime="00:16:35.72" />
                    <SPLIT distance="900" swimtime="00:17:36.29" />
                    <SPLIT distance="950" swimtime="00:18:39.04" />
                    <SPLIT distance="1000" swimtime="00:19:40.39" />
                    <SPLIT distance="1050" swimtime="00:20:42.39" />
                    <SPLIT distance="1100" swimtime="00:21:43.91" />
                    <SPLIT distance="1150" swimtime="00:22:44.45" />
                    <SPLIT distance="1200" swimtime="00:23:44.66" />
                    <SPLIT distance="1250" swimtime="00:24:46.40" />
                    <SPLIT distance="1300" swimtime="00:25:48.43" />
                    <SPLIT distance="1350" swimtime="00:26:49.96" />
                    <SPLIT distance="1400" swimtime="00:27:50.25" />
                    <SPLIT distance="1450" swimtime="00:28:50.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="114" reactiontime="+72" swimtime="00:01:32.49" resultid="7226" heatid="8986" lane="4" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="108" reactiontime="+119" swimtime="00:03:28.65" resultid="7227" heatid="9095" lane="7" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                    <SPLIT distance="100" swimtime="00:01:39.55" />
                    <SPLIT distance="150" swimtime="00:02:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="7228" heatid="9182" lane="4" entrytime="00:08:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-06-11" firstname="Marek" gender="M" lastname="Łukaszewicz" nation="POL" athleteid="1911">
              <RESULTS>
                <RESULT eventid="1079" points="231" reactiontime="+84" swimtime="00:00:33.00" resultid="1912" heatid="8899" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1165" points="176" reactiontime="+88" swimtime="00:25:16.50" resultid="1913" heatid="8941" lane="4" entrytime="00:30:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.55" />
                    <SPLIT distance="100" swimtime="00:01:30.20" />
                    <SPLIT distance="150" swimtime="00:02:18.37" />
                    <SPLIT distance="200" swimtime="00:03:07.03" />
                    <SPLIT distance="250" swimtime="00:03:57.67" />
                    <SPLIT distance="300" swimtime="00:04:47.49" />
                    <SPLIT distance="350" swimtime="00:05:39.28" />
                    <SPLIT distance="400" swimtime="00:06:30.70" />
                    <SPLIT distance="450" swimtime="00:07:23.45" />
                    <SPLIT distance="500" swimtime="00:08:14.96" />
                    <SPLIT distance="550" swimtime="00:09:07.03" />
                    <SPLIT distance="600" swimtime="00:09:57.48" />
                    <SPLIT distance="650" swimtime="00:10:49.39" />
                    <SPLIT distance="700" swimtime="00:11:40.32" />
                    <SPLIT distance="750" swimtime="00:12:31.89" />
                    <SPLIT distance="800" swimtime="00:13:22.42" />
                    <SPLIT distance="850" swimtime="00:14:14.73" />
                    <SPLIT distance="900" swimtime="00:15:05.22" />
                    <SPLIT distance="950" swimtime="00:15:56.68" />
                    <SPLIT distance="1000" swimtime="00:16:46.67" />
                    <SPLIT distance="1050" swimtime="00:17:38.50" />
                    <SPLIT distance="1100" swimtime="00:18:29.39" />
                    <SPLIT distance="1150" swimtime="00:19:22.09" />
                    <SPLIT distance="1200" swimtime="00:20:12.04" />
                    <SPLIT distance="1250" swimtime="00:21:04.57" />
                    <SPLIT distance="1300" swimtime="00:21:55.22" />
                    <SPLIT distance="1350" swimtime="00:22:46.87" />
                    <SPLIT distance="1400" swimtime="00:23:37.27" />
                    <SPLIT distance="1450" swimtime="00:24:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="152" reactiontime="+76" swimtime="00:00:41.59" resultid="1914" heatid="8956" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1341" points="105" reactiontime="+87" swimtime="00:03:49.91" resultid="1915" heatid="9026" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.16" />
                    <SPLIT distance="100" swimtime="00:01:50.31" />
                    <SPLIT distance="150" swimtime="00:02:49.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="187" reactiontime="+89" swimtime="00:00:38.06" resultid="1916" heatid="9063" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1578" points="149" reactiontime="+86" swimtime="00:07:23.81" resultid="1917" heatid="9118" lane="9" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.42" />
                    <SPLIT distance="100" swimtime="00:01:46.33" />
                    <SPLIT distance="150" swimtime="00:02:45.92" />
                    <SPLIT distance="200" swimtime="00:03:45.59" />
                    <SPLIT distance="250" swimtime="00:04:47.95" />
                    <SPLIT distance="300" swimtime="00:05:50.25" />
                    <SPLIT distance="350" swimtime="00:06:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="142" reactiontime="+88" swimtime="00:01:32.68" resultid="1918" heatid="9131" lane="9" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="184" reactiontime="+92" swimtime="00:06:12.89" resultid="1919" heatid="9185" lane="0" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                    <SPLIT distance="100" swimtime="00:01:24.65" />
                    <SPLIT distance="150" swimtime="00:02:11.90" />
                    <SPLIT distance="200" swimtime="00:02:59.66" />
                    <SPLIT distance="250" swimtime="00:03:48.55" />
                    <SPLIT distance="300" swimtime="00:04:37.44" />
                    <SPLIT distance="350" swimtime="00:05:26.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-06-07" firstname="Wiesław" gender="M" lastname="Bar" nation="POL" athleteid="2051">
              <RESULTS>
                <RESULT eventid="1079" points="383" reactiontime="+91" swimtime="00:00:27.89" resultid="2052" heatid="8909" lane="2" entrytime="00:00:27.95" />
                <RESULT eventid="1165" points="362" reactiontime="+98" swimtime="00:19:52.02" resultid="2053" heatid="8946" lane="7" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:11.75" />
                    <SPLIT distance="150" swimtime="00:01:50.78" />
                    <SPLIT distance="200" swimtime="00:02:29.63" />
                    <SPLIT distance="250" swimtime="00:03:09.50" />
                    <SPLIT distance="300" swimtime="00:03:48.26" />
                    <SPLIT distance="350" swimtime="00:04:27.84" />
                    <SPLIT distance="400" swimtime="00:05:07.62" />
                    <SPLIT distance="450" swimtime="00:06:26.89" />
                    <SPLIT distance="550" swimtime="00:07:06.59" />
                    <SPLIT distance="600" swimtime="00:07:46.80" />
                    <SPLIT distance="650" swimtime="00:08:26.91" />
                    <SPLIT distance="800" swimtime="00:10:27.37" />
                    <SPLIT distance="850" swimtime="00:11:07.54" />
                    <SPLIT distance="900" swimtime="00:11:48.37" />
                    <SPLIT distance="950" swimtime="00:12:28.57" />
                    <SPLIT distance="1050" swimtime="00:13:49.12" />
                    <SPLIT distance="1100" swimtime="00:14:29.87" />
                    <SPLIT distance="1150" swimtime="00:15:10.68" />
                    <SPLIT distance="1200" swimtime="00:15:51.38" />
                    <SPLIT distance="1250" swimtime="00:16:31.78" />
                    <SPLIT distance="1300" swimtime="00:17:12.48" />
                    <SPLIT distance="1400" swimtime="00:18:34.37" />
                    <SPLIT distance="1450" swimtime="00:19:14.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="387" reactiontime="+92" swimtime="00:01:01.66" resultid="2054" heatid="8994" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="360" reactiontime="+88" swimtime="00:01:11.16" resultid="2055" heatid="9016" lane="7" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="295" reactiontime="+77" swimtime="00:01:13.48" resultid="2056" heatid="9085" lane="9" entrytime="00:01:10.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="383" reactiontime="+94" swimtime="00:02:16.80" resultid="2057" heatid="9103" lane="0" entrytime="00:02:17.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:07.06" />
                    <SPLIT distance="150" swimtime="00:01:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="381" reactiontime="+96" swimtime="00:04:52.55" resultid="2058" heatid="9190" lane="5" entrytime="00:04:53.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:09.35" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                    <SPLIT distance="200" swimtime="00:02:24.38" />
                    <SPLIT distance="250" swimtime="00:03:02.13" />
                    <SPLIT distance="300" swimtime="00:03:39.15" />
                    <SPLIT distance="350" swimtime="00:04:16.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7088" name="Niezrzeszone Biała Podlaska">
          <ATHLETES>
            <ATHLETE birthdate="1981-11-29" firstname="Iga" gender="F" lastname="Olszanowska" nation="POL" athleteid="6185">
              <RESULTS>
                <RESULT eventid="1096" points="380" reactiontime="+86" swimtime="00:02:48.15" resultid="6186" heatid="8918" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:16.11" />
                    <SPLIT distance="150" swimtime="00:02:05.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="358" reactiontime="+100" swimtime="00:11:14.92" resultid="6187" heatid="8938" lane="6" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                    <SPLIT distance="100" swimtime="00:01:19.66" />
                    <SPLIT distance="150" swimtime="00:02:02.78" />
                    <SPLIT distance="200" swimtime="00:02:46.00" />
                    <SPLIT distance="250" swimtime="00:03:28.87" />
                    <SPLIT distance="300" swimtime="00:04:11.72" />
                    <SPLIT distance="350" swimtime="00:04:54.80" />
                    <SPLIT distance="400" swimtime="00:05:37.47" />
                    <SPLIT distance="450" swimtime="00:06:20.25" />
                    <SPLIT distance="500" swimtime="00:07:02.87" />
                    <SPLIT distance="550" swimtime="00:07:45.25" />
                    <SPLIT distance="600" swimtime="00:08:27.46" />
                    <SPLIT distance="650" swimtime="00:09:09.74" />
                    <SPLIT distance="700" swimtime="00:09:51.76" />
                    <SPLIT distance="750" swimtime="00:10:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="412" reactiontime="+84" swimtime="00:01:16.17" resultid="6188" heatid="9006" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="296" reactiontime="+110" swimtime="00:02:59.38" resultid="6189" heatid="9024" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:21.82" />
                    <SPLIT distance="150" swimtime="00:02:09.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="475" reactiontime="+86" swimtime="00:00:31.24" resultid="6190" heatid="9059" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1555" points="373" reactiontime="+93" swimtime="00:06:00.71" resultid="6191" heatid="9115" lane="8" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:20.12" />
                    <SPLIT distance="150" swimtime="00:02:07.88" />
                    <SPLIT distance="200" swimtime="00:02:54.54" />
                    <SPLIT distance="250" swimtime="00:03:44.65" />
                    <SPLIT distance="300" swimtime="00:04:36.65" />
                    <SPLIT distance="350" swimtime="00:05:20.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="436" reactiontime="+97" swimtime="00:01:11.99" resultid="6192" heatid="9127" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-12-27" firstname="Renata" gender="F" lastname="Kasprowicz" nation="POL" athleteid="6193">
              <RESULTS>
                <RESULT eventid="1062" points="419" reactiontime="+71" swimtime="00:00:31.04" resultid="6194" heatid="8891" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1147" points="202" reactiontime="+87" swimtime="00:13:35.85" resultid="6195" heatid="8937" lane="3" entrytime="00:13:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                    <SPLIT distance="100" swimtime="00:01:23.07" />
                    <SPLIT distance="150" swimtime="00:02:10.72" />
                    <SPLIT distance="200" swimtime="00:03:01.32" />
                    <SPLIT distance="250" swimtime="00:03:53.09" />
                    <SPLIT distance="300" swimtime="00:04:45.05" />
                    <SPLIT distance="350" swimtime="00:05:37.75" />
                    <SPLIT distance="400" swimtime="00:06:29.70" />
                    <SPLIT distance="450" swimtime="00:07:22.06" />
                    <SPLIT distance="500" swimtime="00:08:14.57" />
                    <SPLIT distance="550" swimtime="00:09:06.66" />
                    <SPLIT distance="600" swimtime="00:10:01.49" />
                    <SPLIT distance="650" swimtime="00:10:56.10" />
                    <SPLIT distance="700" swimtime="00:11:51.71" />
                    <SPLIT distance="750" swimtime="00:12:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="378" reactiontime="+77" swimtime="00:01:10.53" resultid="6196" heatid="8983" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="360" reactiontime="+88" swimtime="00:01:19.64" resultid="6197" heatid="9004" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="331" reactiontime="+84" swimtime="00:01:30.12" resultid="6198" heatid="9040" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="364" reactiontime="+77" swimtime="00:00:34.13" resultid="6199" heatid="9057" lane="6" entrytime="00:00:35.20" />
                <RESULT eventid="1664" points="363" reactiontime="+73" swimtime="00:00:40.34" resultid="6200" heatid="9156" lane="5" entrytime="00:00:41.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAŁ" nation="POL" region="MAŁ" clubid="3471" name="niezrzeszony kraków">
          <CONTACT email="piotr_urbanczyk@onet.pl" name="URBAŃCZYK PIOTR" phone="608172201" />
          <ATHLETES>
            <ATHLETE birthdate="1984-03-16" firstname="Piotr" gender="M" lastname="Urbańczyk" nation="POL" athleteid="3472">
              <RESULTS>
                <RESULT eventid="1205" points="412" reactiontime="+70" swimtime="00:00:29.84" resultid="3473" heatid="8965" lane="9" entrytime="00:00:28.12" />
                <RESULT eventid="1474" points="499" reactiontime="+71" swimtime="00:01:01.69" resultid="3474" heatid="9087" lane="6" entrytime="00:01:00.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3764" name="One Man Team">
          <CONTACT city="Daszewice" email="gmo@o2.pl" internet="open-water.pl" name="MONCZAK" street="Przy Lesie" zip="61-160" />
          <ATHLETES>
            <ATHLETE birthdate="1973-05-25" firstname="Grzegorz" gender="M" lastname="Monczak" nation="POL" athleteid="3780">
              <RESULTS>
                <RESULT eventid="1113" points="349" reactiontime="+77" swimtime="00:02:35.70" resultid="3781" heatid="8929" lane="2" entrytime="00:02:31.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="150" swimtime="00:02:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="434" reactiontime="+78" swimtime="00:18:42.48" resultid="3782" heatid="8947" lane="5" entrytime="00:18:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:11.61" />
                    <SPLIT distance="150" swimtime="00:01:49.48" />
                    <SPLIT distance="200" swimtime="00:02:27.30" />
                    <SPLIT distance="250" swimtime="00:03:05.12" />
                    <SPLIT distance="300" swimtime="00:03:42.64" />
                    <SPLIT distance="350" swimtime="00:04:20.58" />
                    <SPLIT distance="400" swimtime="00:04:58.66" />
                    <SPLIT distance="450" swimtime="00:05:36.10" />
                    <SPLIT distance="500" swimtime="00:06:13.63" />
                    <SPLIT distance="550" swimtime="00:06:51.64" />
                    <SPLIT distance="600" swimtime="00:07:29.19" />
                    <SPLIT distance="650" swimtime="00:08:06.69" />
                    <SPLIT distance="700" swimtime="00:08:44.16" />
                    <SPLIT distance="750" swimtime="00:09:21.82" />
                    <SPLIT distance="800" swimtime="00:09:59.85" />
                    <SPLIT distance="850" swimtime="00:10:37.63" />
                    <SPLIT distance="900" swimtime="00:11:15.46" />
                    <SPLIT distance="950" swimtime="00:11:52.56" />
                    <SPLIT distance="1000" swimtime="00:12:30.07" />
                    <SPLIT distance="1050" swimtime="00:13:07.90" />
                    <SPLIT distance="1100" swimtime="00:13:45.45" />
                    <SPLIT distance="1150" swimtime="00:14:23.17" />
                    <SPLIT distance="1200" swimtime="00:15:00.78" />
                    <SPLIT distance="1250" swimtime="00:15:38.54" />
                    <SPLIT distance="1300" swimtime="00:16:15.72" />
                    <SPLIT distance="1350" swimtime="00:16:52.68" />
                    <SPLIT distance="1400" swimtime="00:17:29.60" />
                    <SPLIT distance="1450" swimtime="00:18:06.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="426" reactiontime="+77" swimtime="00:00:59.71" resultid="3783" heatid="8998" lane="2" entrytime="00:00:58.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="341" reactiontime="+72" swimtime="00:01:12.48" resultid="3784" heatid="9017" lane="9" entrytime="00:01:12.00" entrycourse="SCY">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="3785" heatid="9047" lane="6" entrytime="00:01:30.00" />
                <RESULT eventid="1508" points="437" reactiontime="+76" swimtime="00:02:10.92" resultid="3786" heatid="9104" lane="6" entrytime="00:02:09.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:04.60" />
                    <SPLIT distance="150" swimtime="00:01:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="447" reactiontime="+85" swimtime="00:04:37.41" resultid="3787" heatid="9191" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="150" swimtime="00:01:43.60" />
                    <SPLIT distance="200" swimtime="00:02:19.38" />
                    <SPLIT distance="250" swimtime="00:02:54.72" />
                    <SPLIT distance="300" swimtime="00:03:29.69" />
                    <SPLIT distance="350" swimtime="00:04:04.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORSOPOLE" nation="POL" region="OPO" clubid="3339" name="ORS Opole">
          <CONTACT email="wkania62@gmail.com" name="Kania" />
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Waldemar" gender="M" lastname="Kania" nation="POL" athleteid="3340">
              <RESULTS>
                <RESULT eventid="1165" points="223" reactiontime="+93" swimtime="00:23:21.79" resultid="3341" heatid="8944" lane="9" entrytime="00:22:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:24.61" />
                    <SPLIT distance="150" swimtime="00:02:10.44" />
                    <SPLIT distance="200" swimtime="00:02:56.34" />
                    <SPLIT distance="250" swimtime="00:03:42.84" />
                    <SPLIT distance="300" swimtime="00:04:29.90" />
                    <SPLIT distance="350" swimtime="00:05:16.93" />
                    <SPLIT distance="400" swimtime="00:06:04.35" />
                    <SPLIT distance="450" swimtime="00:06:50.95" />
                    <SPLIT distance="500" swimtime="00:07:37.60" />
                    <SPLIT distance="550" swimtime="00:08:24.42" />
                    <SPLIT distance="600" swimtime="00:09:10.66" />
                    <SPLIT distance="650" swimtime="00:09:57.09" />
                    <SPLIT distance="700" swimtime="00:10:44.20" />
                    <SPLIT distance="750" swimtime="00:11:31.50" />
                    <SPLIT distance="800" swimtime="00:12:18.59" />
                    <SPLIT distance="850" swimtime="00:13:05.34" />
                    <SPLIT distance="900" swimtime="00:13:52.37" />
                    <SPLIT distance="950" swimtime="00:14:40.01" />
                    <SPLIT distance="1000" swimtime="00:15:26.86" />
                    <SPLIT distance="1050" swimtime="00:16:13.97" />
                    <SPLIT distance="1100" swimtime="00:17:01.30" />
                    <SPLIT distance="1150" swimtime="00:17:49.06" />
                    <SPLIT distance="1200" swimtime="00:18:36.84" />
                    <SPLIT distance="1250" swimtime="00:19:24.01" />
                    <SPLIT distance="1300" swimtime="00:20:11.37" />
                    <SPLIT distance="1350" swimtime="00:20:59.07" />
                    <SPLIT distance="1400" swimtime="00:21:45.35" />
                    <SPLIT distance="1450" swimtime="00:22:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="238" reactiontime="+101" swimtime="00:02:40.21" resultid="3342" heatid="9098" lane="5" entrytime="00:02:44.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:16.73" />
                    <SPLIT distance="150" swimtime="00:01:59.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="3343" heatid="9186" lane="4" entrytime="00:05:44.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="3344">
              <RESULTS>
                <RESULT eventid="1096" points="392" reactiontime="+78" swimtime="00:02:46.39" resultid="3345" heatid="8920" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:16.79" />
                    <SPLIT distance="150" swimtime="00:02:07.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="3346" heatid="9024" lane="7" entrytime="00:03:01.00" />
                <RESULT eventid="1555" status="DNS" swimtime="00:00:00.00" resultid="3347" heatid="9115" lane="1" entrytime="00:06:10.00" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="3348" heatid="9126" lane="5" entrytime="00:01:18.00" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="3349" heatid="9141" lane="0" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Grzegorz" gender="M" lastname="Stanek" nation="POL" athleteid="3350">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="3351" heatid="8930" lane="0" entrytime="00:02:27.80" />
                <RESULT eventid="1307" points="455" reactiontime="+79" swimtime="00:01:05.86" resultid="3352" heatid="9019" lane="6" entrytime="00:01:06.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="3353" heatid="9105" lane="0" entrytime="00:02:08.90" />
                <RESULT eventid="1744" points="462" reactiontime="+82" swimtime="00:04:34.37" resultid="3354" heatid="9192" lane="9" entrytime="00:04:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:07.23" />
                    <SPLIT distance="150" swimtime="00:01:41.99" />
                    <SPLIT distance="200" swimtime="00:02:17.12" />
                    <SPLIT distance="250" swimtime="00:02:51.73" />
                    <SPLIT distance="300" swimtime="00:03:26.34" />
                    <SPLIT distance="350" swimtime="00:04:00.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Wojciech" gender="M" lastname="Stanek" nation="POL" athleteid="3355">
              <RESULTS>
                <RESULT eventid="1113" points="273" reactiontime="+65" swimtime="00:02:48.98" resultid="3356" heatid="8927" lane="9" entrytime="00:02:49.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:21.32" />
                    <SPLIT distance="150" swimtime="00:02:08.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="284" reactiontime="+84" swimtime="00:01:17.00" resultid="3357" heatid="9014" lane="7" entrytime="00:01:17.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="290" reactiontime="+94" swimtime="00:02:29.99" resultid="3358" heatid="9101" lane="6" entrytime="00:02:22.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:50.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="3359" heatid="9188" lane="5" entrytime="00:05:12.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="9267" name="PK Havirov">
          <ATHLETES>
            <ATHLETE birthdate="1972-08-29" firstname="Libor" gender="M" lastname="Hracki" nation="CZE" athleteid="1892">
              <RESULTS>
                <RESULT eventid="1079" points="308" reactiontime="+82" swimtime="00:00:29.97" resultid="1893" heatid="8906" lane="0" entrytime="00:00:29.50" />
                <RESULT eventid="1165" points="277" reactiontime="+84" swimtime="00:21:42.75" resultid="1894" heatid="8944" lane="2" entrytime="00:22:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:14.65" />
                    <SPLIT distance="150" swimtime="00:01:55.77" />
                    <SPLIT distance="200" swimtime="00:02:37.76" />
                    <SPLIT distance="250" swimtime="00:03:20.39" />
                    <SPLIT distance="300" swimtime="00:04:03.00" />
                    <SPLIT distance="350" swimtime="00:04:46.04" />
                    <SPLIT distance="400" swimtime="00:05:29.94" />
                    <SPLIT distance="450" swimtime="00:06:13.78" />
                    <SPLIT distance="500" swimtime="00:06:57.74" />
                    <SPLIT distance="550" swimtime="00:07:42.50" />
                    <SPLIT distance="600" swimtime="00:08:26.36" />
                    <SPLIT distance="650" swimtime="00:09:10.99" />
                    <SPLIT distance="700" swimtime="00:09:54.89" />
                    <SPLIT distance="750" swimtime="00:10:38.83" />
                    <SPLIT distance="800" swimtime="00:11:22.92" />
                    <SPLIT distance="850" swimtime="00:12:07.11" />
                    <SPLIT distance="900" swimtime="00:12:51.01" />
                    <SPLIT distance="950" swimtime="00:13:35.34" />
                    <SPLIT distance="1000" swimtime="00:14:19.35" />
                    <SPLIT distance="1050" swimtime="00:15:03.64" />
                    <SPLIT distance="1100" swimtime="00:15:47.36" />
                    <SPLIT distance="1150" swimtime="00:16:31.97" />
                    <SPLIT distance="1200" swimtime="00:17:16.09" />
                    <SPLIT distance="1250" swimtime="00:18:00.19" />
                    <SPLIT distance="1300" swimtime="00:18:44.54" />
                    <SPLIT distance="1350" swimtime="00:19:29.37" />
                    <SPLIT distance="1400" swimtime="00:20:14.04" />
                    <SPLIT distance="1450" swimtime="00:20:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="294" reactiontime="+84" swimtime="00:03:01.09" resultid="1895" heatid="8976" lane="6" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:12.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="301" reactiontime="+79" swimtime="00:01:07.05" resultid="1896" heatid="8992" lane="0" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="298" reactiontime="+81" swimtime="00:01:23.17" resultid="1897" heatid="9050" lane="0" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="294" reactiontime="+79" swimtime="00:02:29.31" resultid="1898" heatid="9100" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="150" swimtime="00:01:50.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="3381" name="Pregel">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1963-01-01" firstname="Grigorii" gender="M" lastname="Lopin" nation="RUS" athleteid="3382">
              <RESULTS>
                <RESULT eventid="1165" reactiontime="+99" status="DNF" swimtime="00:00:00.00" resultid="3383" heatid="8943" lane="2" entrytime="00:24:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:26.64" />
                    <SPLIT distance="150" swimtime="00:02:15.01" />
                    <SPLIT distance="200" swimtime="00:03:05.14" />
                    <SPLIT distance="250" swimtime="00:03:57.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="205" reactiontime="+88" swimtime="00:03:24.29" resultid="3384" heatid="8974" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.71" />
                    <SPLIT distance="100" swimtime="00:01:36.59" />
                    <SPLIT distance="150" swimtime="00:02:30.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="248" reactiontime="+88" swimtime="00:01:28.51" resultid="3385" heatid="9048" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="3386" heatid="9119" lane="1" entrytime="00:06:40.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="3387" heatid="9132" lane="9" entrytime="00:01:25.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="3388" heatid="9186" lane="5" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Aleksandr" gender="M" lastname="Smirnov" nation="RUS" athleteid="3396">
              <RESULTS>
                <RESULT eventid="1273" points="402" reactiontime="+82" swimtime="00:01:00.87" resultid="3397" heatid="8997" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="414" reactiontime="+83" swimtime="00:02:13.25" resultid="3398" heatid="9104" lane="8" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                    <SPLIT distance="150" swimtime="00:01:39.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="417" reactiontime="+85" swimtime="00:04:44.05" resultid="3399" heatid="9191" lane="6" entrytime="00:04:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                    <SPLIT distance="150" swimtime="00:01:45.02" />
                    <SPLIT distance="200" swimtime="00:02:21.36" />
                    <SPLIT distance="250" swimtime="00:02:57.71" />
                    <SPLIT distance="300" swimtime="00:03:33.95" />
                    <SPLIT distance="350" swimtime="00:04:09.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Vadim" gender="M" lastname="Ezkov" nation="RUS" athleteid="3389">
              <RESULTS>
                <RESULT eventid="1079" points="291" reactiontime="+81" swimtime="00:00:30.57" resultid="3390" heatid="8904" lane="0" entrytime="00:00:30.50" />
                <RESULT eventid="1113" points="275" reactiontime="+78" swimtime="00:02:48.51" resultid="3391" heatid="8926" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:02:07.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="287" reactiontime="+75" swimtime="00:03:02.46" resultid="3392" heatid="8976" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:24.55" />
                    <SPLIT distance="150" swimtime="00:02:12.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="321" reactiontime="+76" swimtime="00:01:21.16" resultid="3393" heatid="9051" lane="9" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="361" reactiontime="+72" swimtime="00:00:35.44" resultid="3394" heatid="9169" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="3395" heatid="9188" lane="0" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="5088" name="PSK Žilina">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1964-01-01" firstname="Roman" gender="M" lastname="Hrmel" nation="SVK" athleteid="5089">
              <RESULTS>
                <RESULT eventid="1205" points="260" reactiontime="+74" swimtime="00:00:34.80" resultid="5090" heatid="8960" lane="9" entrytime="00:00:34.91" />
                <RESULT eventid="1273" points="327" reactiontime="+79" swimtime="00:01:05.17" resultid="5091" heatid="8993" lane="9" entrytime="00:01:06.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="250" reactiontime="+73" swimtime="00:01:17.68" resultid="5092" heatid="9083" lane="8" entrytime="00:01:18.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Lukas" gender="M" lastname="Smiesko" nation="SVK" athleteid="5102">
              <RESULTS>
                <RESULT eventid="1079" points="568" reactiontime="+73" swimtime="00:00:24.46" resultid="5103" heatid="8915" lane="0" entrytime="00:00:24.12" />
                <RESULT eventid="1113" points="501" reactiontime="+80" swimtime="00:02:17.96" resultid="5104" heatid="8931" lane="0" entrytime="00:02:18.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                    <SPLIT distance="100" swimtime="00:01:04.33" />
                    <SPLIT distance="150" swimtime="00:01:44.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="555" reactiontime="+78" swimtime="00:01:01.64" resultid="5105" heatid="9021" lane="0" entrytime="00:01:01.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="533" reactiontime="+73" swimtime="00:01:08.58" resultid="5106" heatid="9053" lane="7" entrytime="00:01:09.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="519" reactiontime="+68" swimtime="00:00:27.12" resultid="5107" heatid="9073" lane="9" entrytime="00:00:26.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Rastislav" gender="M" lastname="Pavlik" nation="SVK" athleteid="5096">
              <RESULTS>
                <RESULT eventid="1079" points="446" reactiontime="+88" swimtime="00:00:26.50" resultid="5097" heatid="8911" lane="2" entrytime="00:00:26.62" />
                <RESULT eventid="1205" points="397" reactiontime="+73" swimtime="00:00:30.22" resultid="5098" heatid="8963" lane="7" entrytime="00:00:30.65" />
                <RESULT eventid="1307" points="471" reactiontime="+83" swimtime="00:01:05.07" resultid="5099" heatid="9019" lane="5" entrytime="00:01:06.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="441" reactiontime="+94" swimtime="00:01:13.01" resultid="5100" heatid="9052" lane="6" entrytime="00:01:14.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="390" reactiontime="+80" swimtime="00:01:06.93" resultid="5101" heatid="9086" lane="0" entrytime="00:01:07.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Juraj" gender="M" lastname="Jaros" nation="SVK" athleteid="5093">
              <RESULTS>
                <RESULT eventid="1239" points="222" reactiontime="+86" swimtime="00:03:18.83" resultid="5094" heatid="8974" lane="7" entrytime="00:03:21.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                    <SPLIT distance="100" swimtime="00:01:34.67" />
                    <SPLIT distance="150" swimtime="00:02:26.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="250" reactiontime="+82" swimtime="00:01:28.16" resultid="5095" heatid="9048" lane="3" entrytime="00:01:28.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Denisa" gender="F" lastname="Zabkova" nation="SVK" athleteid="5108">
              <RESULTS>
                <RESULT eventid="1256" points="220" reactiontime="+100" swimtime="00:01:24.40" resultid="5109" heatid="8980" lane="7" entrytime="00:01:30.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="147" reactiontime="+75" swimtime="00:01:44.21" resultid="5110" heatid="9075" lane="3" entrytime="00:01:46.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02705" nation="POL" region="SLA" clubid="3664" name="Pływak Tomaszów Maz">
          <CONTACT name="Bucholz" phone="606135860" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-26" firstname="Tomasz" gender="M" lastname="Bucholz" nation="POL" athleteid="3665">
              <RESULTS>
                <RESULT eventid="1165" points="359" reactiontime="+114" swimtime="00:19:56.05" resultid="3666" heatid="8946" lane="0" entrytime="00:21:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:01:52.55" />
                    <SPLIT distance="200" swimtime="00:02:32.52" />
                    <SPLIT distance="250" swimtime="00:03:12.16" />
                    <SPLIT distance="300" swimtime="00:03:50.17" />
                    <SPLIT distance="350" swimtime="00:04:30.14" />
                    <SPLIT distance="400" swimtime="00:05:10.21" />
                    <SPLIT distance="450" swimtime="00:05:50.22" />
                    <SPLIT distance="500" swimtime="00:06:30.09" />
                    <SPLIT distance="550" swimtime="00:07:08.92" />
                    <SPLIT distance="600" swimtime="00:07:49.24" />
                    <SPLIT distance="650" swimtime="00:08:29.38" />
                    <SPLIT distance="700" swimtime="00:09:09.69" />
                    <SPLIT distance="750" swimtime="00:09:50.09" />
                    <SPLIT distance="800" swimtime="00:10:29.69" />
                    <SPLIT distance="850" swimtime="00:11:09.70" />
                    <SPLIT distance="900" swimtime="00:11:50.32" />
                    <SPLIT distance="950" swimtime="00:12:30.77" />
                    <SPLIT distance="1000" swimtime="00:13:11.62" />
                    <SPLIT distance="1050" swimtime="00:13:52.23" />
                    <SPLIT distance="1100" swimtime="00:14:32.99" />
                    <SPLIT distance="1150" swimtime="00:15:12.81" />
                    <SPLIT distance="1200" swimtime="00:15:53.80" />
                    <SPLIT distance="1250" swimtime="00:16:33.93" />
                    <SPLIT distance="1300" swimtime="00:17:14.06" />
                    <SPLIT distance="1350" swimtime="00:17:55.03" />
                    <SPLIT distance="1400" swimtime="00:18:36.42" />
                    <SPLIT distance="1450" swimtime="00:19:17.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-13" firstname="Damian" gender="M" lastname="Hostyński" nation="POL" athleteid="3667" />
            <ATHLETE birthdate="1973-08-30" firstname="Jacek" gender="M" lastname="Kobylczak" nation="POL" athleteid="3668" />
            <ATHLETE birthdate="1972-05-02" firstname="Mateusz" gender="M" lastname="Matusiewicz" nation="POL" athleteid="3669" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="295" reactiontime="+109" swimtime="00:02:04.03" resultid="3670" heatid="9110" lane="0" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                    <SPLIT distance="100" swimtime="00:01:03.48" />
                    <SPLIT distance="150" swimtime="00:01:34.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3667" number="1" reactiontime="+109" />
                    <RELAYPOSITION athleteid="3669" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="3668" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3665" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="259" reactiontime="+88" swimtime="00:02:21.94" resultid="3671" heatid="9032" lane="3" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:16.60" />
                    <SPLIT distance="150" swimtime="00:01:50.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3668" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3667" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3665" number="3" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3669" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="5538" name="Redeco Wrocław">
          <CONTACT city="Wrocław" name="Wolny Dariusz" phone="603630870" state="DOL" street="Rogowska 52a" zip="54-440" />
          <ATHLETES>
            <ATHLETE birthdate="1970-02-10" firstname="Artur" gender="M" lastname="Malina" nation="POL" athleteid="5545">
              <RESULTS>
                <RESULT eventid="1079" points="183" reactiontime="+119" swimtime="00:00:35.68" resultid="5546" heatid="8899" lane="1" entrytime="00:00:35.80" />
                <RESULT eventid="1239" points="170" reactiontime="+117" swimtime="00:03:37.41" resultid="5547" heatid="8973" lane="7" entrytime="00:03:38.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.60" />
                    <SPLIT distance="100" swimtime="00:01:45.64" />
                    <SPLIT distance="150" swimtime="00:02:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="149" reactiontime="+116" swimtime="00:01:24.73" resultid="5548" heatid="8988" lane="7" entrytime="00:01:23.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="189" reactiontime="+111" swimtime="00:01:36.74" resultid="5549" heatid="9046" lane="9" entrytime="00:01:38.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="128" reactiontime="+117" swimtime="00:03:16.73" resultid="5550" heatid="9096" lane="6" entrytime="00:03:18.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="100" swimtime="00:01:30.59" />
                    <SPLIT distance="150" swimtime="00:02:22.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="207" reactiontime="+109" swimtime="00:00:42.65" resultid="5551" heatid="9162" lane="3" entrytime="00:00:44.09" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-03" firstname="Łukasz" gender="M" lastname="Hałada" nation="POL" athleteid="5584">
              <RESULTS>
                <RESULT eventid="1079" points="390" reactiontime="+82" swimtime="00:00:27.72" resultid="5585" heatid="8910" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1205" points="327" reactiontime="+65" swimtime="00:00:32.22" resultid="5586" heatid="8962" lane="3" entrytime="00:00:31.11" />
                <RESULT eventid="1273" points="399" reactiontime="+75" swimtime="00:01:01.02" resultid="5587" heatid="8996" lane="1" entrytime="00:01:01.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="332" reactiontime="+66" swimtime="00:01:10.61" resultid="5588" heatid="9084" lane="4" entrytime="00:01:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="294" reactiontime="+75" swimtime="00:02:39.50" resultid="5589" heatid="9148" lane="0" entrytime="00:02:40.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:01:58.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-13" firstname="Kazimiera" gender="F" lastname="Syguła" nation="POL" athleteid="5567">
              <RESULTS>
                <RESULT eventid="1096" points="112" reactiontime="+115" swimtime="00:04:12.50" resultid="5568" heatid="8917" lane="9" entrytime="00:04:08.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.75" />
                    <SPLIT distance="100" swimtime="00:01:58.00" />
                    <SPLIT distance="150" swimtime="00:03:11.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="117" reactiontime="+105" swimtime="00:01:55.82" resultid="5569" heatid="9002" lane="9" entrytime="00:01:57.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="108" reactiontime="+102" swimtime="00:01:55.41" resultid="5570" heatid="9075" lane="1" entrytime="00:01:55.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="120" reactiontime="+104" swimtime="00:04:01.52" resultid="5571" heatid="9139" lane="1" entrytime="00:04:02.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.92" />
                    <SPLIT distance="100" swimtime="00:01:58.30" />
                    <SPLIT distance="150" swimtime="00:03:00.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-12-13" firstname="Agata" gender="F" lastname="Grochowska" nation="POL" athleteid="5590">
              <RESULTS>
                <RESULT eventid="1062" points="231" reactiontime="+93" swimtime="00:00:37.86" resultid="5591" heatid="8887" lane="3" entrytime="00:00:40.95" />
                <RESULT eventid="1096" points="175" reactiontime="+99" swimtime="00:03:37.86" resultid="5592" heatid="8917" lane="7" entrytime="00:03:45.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.36" />
                    <SPLIT distance="100" swimtime="00:01:42.79" />
                    <SPLIT distance="150" swimtime="00:02:44.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="213" reactiontime="+78" swimtime="00:00:42.95" resultid="5593" heatid="8949" lane="5" entrytime="00:00:47.25" />
                <RESULT eventid="1290" points="211" reactiontime="+96" swimtime="00:01:35.11" resultid="5594" heatid="9003" lane="8" entrytime="00:01:39.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="158" reactiontime="+75" swimtime="00:00:45.09" resultid="5595" heatid="9055" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="1457" points="185" reactiontime="+68" swimtime="00:01:36.41" resultid="5596" heatid="9075" lane="5" entrytime="00:01:42.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-14" firstname="Anna" gender="F" lastname="Jaśkiewicz" nation="POL" athleteid="5559">
              <RESULTS>
                <RESULT eventid="1096" points="244" reactiontime="+99" swimtime="00:03:15.01" resultid="5560" heatid="8918" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:34.79" />
                    <SPLIT distance="150" swimtime="00:02:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="213" reactiontime="+96" swimtime="00:13:21.54" resultid="5561" heatid="8937" lane="4" entrytime="00:13:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:26.49" />
                    <SPLIT distance="150" swimtime="00:02:16.13" />
                    <SPLIT distance="200" swimtime="00:03:07.20" />
                    <SPLIT distance="250" swimtime="00:03:57.97" />
                    <SPLIT distance="300" swimtime="00:04:49.29" />
                    <SPLIT distance="350" swimtime="00:05:40.28" />
                    <SPLIT distance="400" swimtime="00:06:31.53" />
                    <SPLIT distance="450" swimtime="00:07:23.02" />
                    <SPLIT distance="500" swimtime="00:08:14.40" />
                    <SPLIT distance="550" swimtime="00:09:05.24" />
                    <SPLIT distance="600" swimtime="00:09:56.87" />
                    <SPLIT distance="650" swimtime="00:10:48.88" />
                    <SPLIT distance="700" swimtime="00:11:40.93" />
                    <SPLIT distance="750" swimtime="00:12:32.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="297" reactiontime="+104" swimtime="00:03:21.66" resultid="5562" heatid="8970" lane="0" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:36.67" />
                    <SPLIT distance="150" swimtime="00:02:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="294" reactiontime="+98" swimtime="00:01:33.69" resultid="5563" heatid="9040" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="260" reactiontime="+86" swimtime="00:02:53.46" resultid="5564" heatid="9091" lane="9" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:01:22.56" />
                    <SPLIT distance="150" swimtime="00:02:09.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="306" reactiontime="+93" swimtime="00:00:42.70" resultid="5565" heatid="9156" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1721" points="226" reactiontime="+98" swimtime="00:06:24.81" resultid="5566" heatid="9179" lane="7" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.62" />
                    <SPLIT distance="200" swimtime="00:03:09.34" />
                    <SPLIT distance="250" swimtime="00:04:00.02" />
                    <SPLIT distance="300" swimtime="00:04:50.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-09-09" firstname="Michał" gender="M" lastname="Kula" nation="POL" athleteid="5539">
              <RESULTS>
                <RESULT eventid="1079" points="532" reactiontime="+88" swimtime="00:00:24.99" resultid="5540" heatid="8911" lane="9" entrytime="00:00:26.80" />
                <RESULT eventid="1205" points="485" reactiontime="+65" swimtime="00:00:28.27" resultid="5541" heatid="8962" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1273" points="548" reactiontime="+86" swimtime="00:00:54.91" resultid="5542" heatid="8997" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="458" reactiontime="+86" swimtime="00:00:28.27" resultid="5543" heatid="9070" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1474" points="526" reactiontime="+61" swimtime="00:01:00.59" resultid="5544" heatid="9085" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-11-30" firstname="Ryszard" gender="M" lastname="Sowiński" nation="POL" athleteid="6931">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="6932" heatid="8896" lane="0" entrytime="00:00:49.00" />
                <RESULT eventid="1165" points="74" swimtime="00:33:39.28" resultid="6933" heatid="8941" lane="2" entrytime="00:32:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.63" />
                    <SPLIT distance="150" swimtime="00:03:11.66" />
                    <SPLIT distance="200" swimtime="00:04:15.60" />
                    <SPLIT distance="250" swimtime="00:05:22.61" />
                    <SPLIT distance="300" swimtime="00:07:35.57" />
                    <SPLIT distance="350" swimtime="00:08:42.91" />
                    <SPLIT distance="400" swimtime="00:09:52.57" />
                    <SPLIT distance="450" swimtime="00:11:03.01" />
                    <SPLIT distance="500" swimtime="00:12:12.23" />
                    <SPLIT distance="550" swimtime="00:13:23.00" />
                    <SPLIT distance="600" swimtime="00:14:33.02" />
                    <SPLIT distance="650" swimtime="00:15:40.23" />
                    <SPLIT distance="700" swimtime="00:16:49.64" />
                    <SPLIT distance="750" swimtime="00:17:58.00" />
                    <SPLIT distance="800" swimtime="00:19:03.85" />
                    <SPLIT distance="850" swimtime="00:20:13.55" />
                    <SPLIT distance="900" swimtime="00:21:21.73" />
                    <SPLIT distance="950" swimtime="00:22:30.64" />
                    <SPLIT distance="1000" swimtime="00:23:38.41" />
                    <SPLIT distance="1050" swimtime="00:24:45.23" />
                    <SPLIT distance="1100" swimtime="00:25:51.65" />
                    <SPLIT distance="1150" swimtime="00:26:52.88" />
                    <SPLIT distance="1200" swimtime="00:28:01.16" />
                    <SPLIT distance="1250" swimtime="00:29:05.43" />
                    <SPLIT distance="1300" swimtime="00:30:10.33" />
                    <SPLIT distance="1350" swimtime="00:31:16.62" />
                    <SPLIT distance="1400" swimtime="00:32:23.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-12-31" firstname="Agata" gender="F" lastname="Szydło" nation="POL" athleteid="5572">
              <RESULTS>
                <RESULT eventid="1147" points="174" reactiontime="+104" swimtime="00:14:18.29" resultid="5573" heatid="8936" lane="4" entrytime="00:15:55.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.80" />
                    <SPLIT distance="100" swimtime="00:01:38.96" />
                    <SPLIT distance="150" swimtime="00:02:31.74" />
                    <SPLIT distance="200" swimtime="00:03:25.34" />
                    <SPLIT distance="250" swimtime="00:04:18.79" />
                    <SPLIT distance="300" swimtime="00:05:12.98" />
                    <SPLIT distance="350" swimtime="00:06:06.87" />
                    <SPLIT distance="400" swimtime="00:07:01.35" />
                    <SPLIT distance="450" swimtime="00:07:54.98" />
                    <SPLIT distance="500" swimtime="00:08:49.48" />
                    <SPLIT distance="550" swimtime="00:09:43.77" />
                    <SPLIT distance="600" swimtime="00:10:45.36" />
                    <SPLIT distance="650" swimtime="00:11:39.57" />
                    <SPLIT distance="700" swimtime="00:12:33.36" />
                    <SPLIT distance="750" swimtime="00:13:27.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="206" reactiontime="+111" swimtime="00:03:47.85" resultid="5574" heatid="8968" lane="3" entrytime="00:03:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.80" />
                    <SPLIT distance="100" swimtime="00:01:50.92" />
                    <SPLIT distance="150" swimtime="00:02:49.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="169" reactiontime="+107" swimtime="00:01:42.42" resultid="5575" heatid="9003" lane="2" entrytime="00:01:38.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="184" reactiontime="+113" swimtime="00:01:49.51" resultid="5576" heatid="9038" lane="6" entrytime="00:01:50.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="179" reactiontime="+104" swimtime="00:03:16.50" resultid="5577" heatid="9089" lane="3" entrytime="00:03:26.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.62" />
                    <SPLIT distance="100" swimtime="00:01:36.63" />
                    <SPLIT distance="150" swimtime="00:02:27.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="179" reactiontime="+99" swimtime="00:00:51.04" resultid="5578" heatid="9153" lane="1" entrytime="00:00:53.81" />
                <RESULT eventid="1721" points="188" reactiontime="+99" swimtime="00:06:49.23" resultid="5579" heatid="9178" lane="4" entrytime="00:06:45.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                    <SPLIT distance="100" swimtime="00:01:36.67" />
                    <SPLIT distance="150" swimtime="00:02:28.47" />
                    <SPLIT distance="200" swimtime="00:03:20.86" />
                    <SPLIT distance="250" swimtime="00:04:13.66" />
                    <SPLIT distance="300" swimtime="00:05:06.15" />
                    <SPLIT distance="350" swimtime="00:05:58.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-01" firstname="Wojciech" gender="M" lastname="Dobrowolski" nation="POL" athleteid="5580">
              <RESULTS>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="5581" heatid="8994" lane="1" entrytime="00:01:04.00" />
                <RESULT eventid="1440" points="310" reactiontime="+86" swimtime="00:00:32.19" resultid="5582" heatid="9067" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1613" points="223" reactiontime="+86" swimtime="00:01:19.84" resultid="5583" heatid="9132" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-13" firstname="Małgorzata" gender="F" lastname="Bołtuć" nation="POL" athleteid="5552">
              <RESULTS>
                <RESULT eventid="1096" points="194" reactiontime="+113" swimtime="00:03:30.44" resultid="5553" heatid="8917" lane="5" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:43.13" />
                    <SPLIT distance="150" swimtime="00:02:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="192" reactiontime="+113" swimtime="00:13:49.58" resultid="5554" heatid="8937" lane="8" entrytime="00:14:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                    <SPLIT distance="100" swimtime="00:01:37.43" />
                    <SPLIT distance="150" swimtime="00:02:28.57" />
                    <SPLIT distance="200" swimtime="00:03:19.35" />
                    <SPLIT distance="250" swimtime="00:04:11.70" />
                    <SPLIT distance="300" swimtime="00:05:04.36" />
                    <SPLIT distance="350" swimtime="00:05:59.05" />
                    <SPLIT distance="400" swimtime="00:06:50.93" />
                    <SPLIT distance="450" swimtime="00:07:44.72" />
                    <SPLIT distance="500" swimtime="00:08:36.41" />
                    <SPLIT distance="550" swimtime="00:09:29.24" />
                    <SPLIT distance="600" swimtime="00:10:23.23" />
                    <SPLIT distance="650" swimtime="00:11:16.12" />
                    <SPLIT distance="700" swimtime="00:12:08.55" />
                    <SPLIT distance="750" swimtime="00:13:00.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="193" reactiontime="+112" swimtime="00:03:52.58" resultid="5555" heatid="8968" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.24" />
                    <SPLIT distance="100" swimtime="00:01:54.99" />
                    <SPLIT distance="150" swimtime="00:02:54.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="181" reactiontime="+114" swimtime="00:01:40.06" resultid="5556" heatid="9003" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="150" reactiontime="+111" swimtime="00:00:45.83" resultid="5557" heatid="9055" lane="7" entrytime="00:00:48.00" />
                <RESULT eventid="1721" points="179" reactiontime="+110" swimtime="00:06:55.37" resultid="5558" heatid="9179" lane="9" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.23" />
                    <SPLIT distance="100" swimtime="00:01:37.61" />
                    <SPLIT distance="150" swimtime="00:02:29.91" />
                    <SPLIT distance="200" swimtime="00:03:23.10" />
                    <SPLIT distance="250" swimtime="00:04:16.06" />
                    <SPLIT distance="300" swimtime="00:05:10.83" />
                    <SPLIT distance="350" swimtime="00:06:04.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="5597" heatid="9107" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5552" number="1" />
                    <RELAYPOSITION athleteid="5590" number="2" />
                    <RELAYPOSITION athleteid="5559" number="3" />
                    <RELAYPOSITION athleteid="5572" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1358" points="188" reactiontime="+109" swimtime="00:03:01.56" resultid="5598" heatid="9031" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.66" />
                    <SPLIT distance="100" swimtime="00:01:42.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5552" number="1" reactiontime="+109" />
                    <RELAYPOSITION athleteid="5559" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="5567" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5572" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="239" reactiontime="+94" swimtime="00:02:13.09" resultid="5599" heatid="8934" lane="1" entrytime="00:02:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                    <SPLIT distance="100" swimtime="00:01:02.61" />
                    <SPLIT distance="150" swimtime="00:01:40.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5584" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="5545" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="5590" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="5559" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT comment="S4 - Przedwczesna zmiana sztafetowa (stopy pływaka utraciły kontakt z platformą startową słupka zanim poprzedzający go pływak dotkną ściany) (Time: 11:34), Na 3 zmianie" eventid="1698" reactiontime="+67" status="DSQ" swimtime="00:02:31.10" resultid="5600" heatid="9173" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:24.76" />
                    <SPLIT distance="150" swimtime="00:01:58.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5584" number="1" reactiontime="+67" status="DSQ" />
                    <RELAYPOSITION athleteid="5552" number="2" reactiontime="+56" status="DSQ" />
                    <RELAYPOSITION athleteid="5580" number="3" reactiontime="+35" status="DSQ" />
                    <RELAYPOSITION athleteid="5559" number="4" reactiontime="-32" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="RMKS" nation="POL" region="SLA" clubid="3428" name="Rmks Rybnik">
          <CONTACT city="Rybnik" email="aniaduda0511@tlen.pl" name="Duda Anna" phone="792666159" state="SLA" street="orzepowicka 22a/37" zip="44-217" />
          <ATHLETES>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="3439">
              <RESULTS>
                <RESULT eventid="1062" points="534" reactiontime="+83" swimtime="00:00:28.63" resultid="3440" heatid="8893" lane="8" entrytime="00:00:28.80" />
                <RESULT eventid="1256" points="494" reactiontime="+86" swimtime="00:01:04.52" resultid="3441" heatid="8984" lane="1" entrytime="00:01:04.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="494" reactiontime="+89" swimtime="00:00:30.83" resultid="3442" heatid="9059" lane="1" entrytime="00:00:30.80" />
                <RESULT eventid="1491" points="420" reactiontime="+91" swimtime="00:02:27.88" resultid="3443" heatid="9093" lane="8" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:51.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="404" reactiontime="+88" swimtime="00:01:13.87" resultid="3444" heatid="9127" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="394" reactiontime="+91" swimtime="00:00:39.26" resultid="3445" heatid="9158" lane="0" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-11-07" firstname="Iwona" gender="F" lastname="Cymerman" nation="POL" athleteid="3435">
              <RESULTS>
                <RESULT eventid="1290" points="473" reactiontime="+88" swimtime="00:01:12.76" resultid="3436" heatid="9006" lane="3" entrytime="00:01:16.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="414" reactiontime="+87" swimtime="00:00:32.69" resultid="3437" heatid="9058" lane="2" entrytime="00:00:33.80" />
                <RESULT eventid="1664" points="433" reactiontime="+85" swimtime="00:00:38.06" resultid="3438" heatid="9158" lane="8" entrytime="00:00:38.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-03" firstname="Agnieszka" gender="F" lastname="Bieniak" nation="POL" athleteid="3429">
              <RESULTS>
                <RESULT eventid="1187" points="419" reactiontime="+72" swimtime="00:00:34.28" resultid="3430" heatid="8952" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1290" points="440" reactiontime="+88" swimtime="00:01:14.54" resultid="3431" heatid="9006" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="427" reactiontime="+86" swimtime="00:00:32.36" resultid="3432" heatid="9058" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1457" points="429" reactiontime="+106" swimtime="00:01:12.95" resultid="3433" heatid="9078" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="454" reactiontime="+89" swimtime="00:00:37.46" resultid="3434" heatid="9158" lane="1" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SLO" clubid="4222" name="RUDAR Trbovlje">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1963-07-18" firstname="Boris" gender="M" lastname="Novak" nation="SLO" athleteid="4223">
              <RESULTS>
                <RESULT eventid="1205" points="347" reactiontime="+64" swimtime="00:00:31.60" resultid="4224" heatid="8962" lane="7" entrytime="00:00:31.97" />
                <RESULT eventid="1307" points="385" reactiontime="+81" swimtime="00:01:09.58" resultid="4225" heatid="9018" lane="2" entrytime="00:01:09.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="348" reactiontime="+65" swimtime="00:01:09.54" resultid="4226" heatid="9085" lane="6" entrytime="00:01:08.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="315" reactiontime="+63" swimtime="00:02:35.93" resultid="4227" heatid="9149" lane="9" entrytime="00:02:34.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:01:56.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1954" name="Rydułtowska Akademia Aktywnego Seniora 60+" shortname="Rydułtowska Akademia Aktywnego">
          <CONTACT email="otelom.080966@intreria.pl" name="OTLIK Marian" phone="692112775" />
          <ATHLETES>
            <ATHLETE birthdate="1966-09-08" firstname="Marian" gender="M" lastname="Otlik" nation="POL" athleteid="2006">
              <RESULTS>
                <RESULT eventid="1079" points="306" reactiontime="+71" swimtime="00:00:30.05" resultid="2007" heatid="8905" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1113" points="207" reactiontime="+77" swimtime="00:03:05.30" resultid="2008" heatid="8924" lane="6" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="100" swimtime="00:01:26.54" />
                    <SPLIT distance="150" swimtime="00:02:22.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="262" reactiontime="+64" swimtime="00:01:10.17" resultid="2009" heatid="8992" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="235" reactiontime="+79" swimtime="00:01:22.01" resultid="2010" heatid="9012" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="244" reactiontime="+74" swimtime="00:00:34.86" resultid="2011" heatid="9065" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1508" points="222" reactiontime="+74" swimtime="00:02:43.87" resultid="2012" heatid="9099" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:02:02.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="176" reactiontime="+76" swimtime="00:01:26.35" resultid="2013" heatid="9131" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="198" reactiontime="+71" swimtime="00:00:43.28" resultid="2014" heatid="9164" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-07" firstname="Leon" gender="M" lastname="Irczyk" nation="POL" athleteid="1973">
              <RESULTS>
                <RESULT eventid="1113" points="86" reactiontime="+119" swimtime="00:04:07.45" resultid="1974" heatid="8922" lane="2" entrytime="00:03:54.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.54" />
                    <SPLIT distance="100" swimtime="00:02:12.14" />
                    <SPLIT distance="150" swimtime="00:03:10.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="108" reactiontime="+124" swimtime="00:29:42.59" resultid="1975" heatid="8942" lane="9" entrytime="00:29:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                    <SPLIT distance="100" swimtime="00:01:49.73" />
                    <SPLIT distance="150" swimtime="00:02:48.71" />
                    <SPLIT distance="200" swimtime="00:03:47.98" />
                    <SPLIT distance="250" swimtime="00:04:47.03" />
                    <SPLIT distance="300" swimtime="00:05:46.60" />
                    <SPLIT distance="350" swimtime="00:06:45.14" />
                    <SPLIT distance="400" swimtime="00:07:45.47" />
                    <SPLIT distance="450" swimtime="00:08:45.71" />
                    <SPLIT distance="500" swimtime="00:09:46.00" />
                    <SPLIT distance="550" swimtime="00:10:45.91" />
                    <SPLIT distance="600" swimtime="00:11:45.68" />
                    <SPLIT distance="650" swimtime="00:12:46.60" />
                    <SPLIT distance="700" swimtime="00:13:46.27" />
                    <SPLIT distance="750" swimtime="00:14:45.92" />
                    <SPLIT distance="800" swimtime="00:15:45.68" />
                    <SPLIT distance="850" swimtime="00:16:46.43" />
                    <SPLIT distance="900" swimtime="00:17:46.35" />
                    <SPLIT distance="950" swimtime="00:18:46.62" />
                    <SPLIT distance="1000" swimtime="00:19:46.72" />
                    <SPLIT distance="1050" swimtime="00:20:47.11" />
                    <SPLIT distance="1100" swimtime="00:21:47.89" />
                    <SPLIT distance="1150" swimtime="00:22:48.46" />
                    <SPLIT distance="1200" swimtime="00:23:48.64" />
                    <SPLIT distance="1250" swimtime="00:24:48.38" />
                    <SPLIT distance="1300" swimtime="00:25:48.92" />
                    <SPLIT distance="1350" swimtime="00:26:48.14" />
                    <SPLIT distance="1400" swimtime="00:27:48.32" />
                    <SPLIT distance="1450" swimtime="00:28:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="146" reactiontime="+115" swimtime="00:03:48.76" resultid="1976" heatid="8973" lane="9" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.14" />
                    <SPLIT distance="100" swimtime="00:01:52.66" />
                    <SPLIT distance="150" swimtime="00:02:51.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="83" reactiontime="+128" swimtime="00:01:42.76" resultid="1977" heatid="8985" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="137" reactiontime="+115" swimtime="00:01:47.83" resultid="1978" heatid="9045" lane="3" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="1979" heatid="9117" lane="8" entrytime="00:08:30.00" />
                <RESULT eventid="1681" points="132" reactiontime="+110" swimtime="00:00:49.51" resultid="1980" heatid="9161" lane="3" entrytime="00:00:49.00" />
                <RESULT eventid="1744" points="101" reactiontime="+136" swimtime="00:07:35.57" resultid="1981" heatid="9183" lane="1" entrytime="00:07:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.33" />
                    <SPLIT distance="100" swimtime="00:01:49.40" />
                    <SPLIT distance="150" swimtime="00:02:49.22" />
                    <SPLIT distance="200" swimtime="00:03:48.88" />
                    <SPLIT distance="250" swimtime="00:04:47.89" />
                    <SPLIT distance="300" swimtime="00:05:45.18" />
                    <SPLIT distance="350" swimtime="00:06:42.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="1964">
              <RESULTS>
                <RESULT eventid="1113" points="161" reactiontime="+92" swimtime="00:03:21.21" resultid="1965" heatid="8924" lane="2" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                    <SPLIT distance="100" swimtime="00:01:34.40" />
                    <SPLIT distance="150" swimtime="00:02:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="193" reactiontime="+89" swimtime="00:24:29.64" resultid="1966" heatid="8943" lane="7" entrytime="00:24:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="100" swimtime="00:01:29.54" />
                    <SPLIT distance="150" swimtime="00:02:17.97" />
                    <SPLIT distance="200" swimtime="00:03:07.22" />
                    <SPLIT distance="250" swimtime="00:03:56.48" />
                    <SPLIT distance="300" swimtime="00:04:46.08" />
                    <SPLIT distance="350" swimtime="00:05:35.55" />
                    <SPLIT distance="400" swimtime="00:06:24.67" />
                    <SPLIT distance="450" swimtime="00:07:14.38" />
                    <SPLIT distance="500" swimtime="00:08:03.39" />
                    <SPLIT distance="550" swimtime="00:08:52.83" />
                    <SPLIT distance="600" swimtime="00:09:42.32" />
                    <SPLIT distance="650" swimtime="00:10:31.91" />
                    <SPLIT distance="700" swimtime="00:11:21.15" />
                    <SPLIT distance="750" swimtime="00:12:11.01" />
                    <SPLIT distance="800" swimtime="00:13:00.01" />
                    <SPLIT distance="850" swimtime="00:13:49.57" />
                    <SPLIT distance="900" swimtime="00:14:39.25" />
                    <SPLIT distance="950" swimtime="00:15:28.81" />
                    <SPLIT distance="1000" swimtime="00:16:18.34" />
                    <SPLIT distance="1050" swimtime="00:17:08.08" />
                    <SPLIT distance="1100" swimtime="00:17:57.93" />
                    <SPLIT distance="1150" swimtime="00:18:47.70" />
                    <SPLIT distance="1200" swimtime="00:19:37.75" />
                    <SPLIT distance="1250" swimtime="00:20:27.19" />
                    <SPLIT distance="1300" swimtime="00:21:17.18" />
                    <SPLIT distance="1350" swimtime="00:22:06.54" />
                    <SPLIT distance="1400" swimtime="00:22:55.92" />
                    <SPLIT distance="1450" swimtime="00:23:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="158" reactiontime="+74" swimtime="00:00:41.10" resultid="1967" heatid="8957" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1341" points="117" reactiontime="+103" swimtime="00:03:41.59" resultid="1968" heatid="9027" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.20" />
                    <SPLIT distance="100" swimtime="00:01:42.41" />
                    <SPLIT distance="150" swimtime="00:02:43.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="161" reactiontime="+79" swimtime="00:01:29.79" resultid="1969" heatid="9081" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="168" reactiontime="+92" swimtime="00:07:06.79" resultid="1970" heatid="9118" lane="8" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                    <SPLIT distance="100" swimtime="00:01:41.53" />
                    <SPLIT distance="200" swimtime="00:03:32.38" />
                    <SPLIT distance="250" swimtime="00:04:35.29" />
                    <SPLIT distance="300" swimtime="00:05:35.80" />
                    <SPLIT distance="350" swimtime="00:06:22.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="162" reactiontime="+90" swimtime="00:01:28.80" resultid="1971" heatid="9131" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="144" reactiontime="+91" swimtime="00:03:22.13" resultid="1972" heatid="9146" lane="8" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                    <SPLIT distance="100" swimtime="00:01:37.23" />
                    <SPLIT distance="150" swimtime="00:02:30.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-02-02" firstname="Maria" gender="F" lastname="Lippa" nation="POL" athleteid="1997">
              <RESULTS>
                <RESULT eventid="1062" points="31" reactiontime="+131" swimtime="00:01:13.69" resultid="1998" heatid="8885" lane="4" />
                <RESULT eventid="1147" reactiontime="+136" status="OTL" swimtime="00:00:00.00" resultid="1999" heatid="8936" lane="6" entrytime="00:19:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.86" />
                    <SPLIT distance="100" swimtime="00:02:37.24" />
                    <SPLIT distance="150" swimtime="00:04:03.21" />
                    <SPLIT distance="200" swimtime="00:05:29.47" />
                    <SPLIT distance="250" swimtime="00:06:54.00" />
                    <SPLIT distance="300" swimtime="00:08:19.09" />
                    <SPLIT distance="350" swimtime="00:09:44.87" />
                    <SPLIT distance="400" swimtime="00:11:10.04" />
                    <SPLIT distance="450" swimtime="00:12:35.10" />
                    <SPLIT distance="500" swimtime="00:13:58.74" />
                    <SPLIT distance="550" swimtime="00:15:23.76" />
                    <SPLIT distance="600" swimtime="00:16:49.33" />
                    <SPLIT distance="650" swimtime="00:18:13.35" />
                    <SPLIT distance="700" swimtime="00:19:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="25" reactiontime="+139" swimtime="00:01:26.83" resultid="2000" heatid="8948" lane="2" />
                <RESULT eventid="1222" points="40" reactiontime="+153" swimtime="00:06:33.12" resultid="2001" heatid="8966" lane="4" entrytime="00:06:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.94" />
                    <SPLIT distance="100" swimtime="00:03:12.35" />
                    <SPLIT distance="150" swimtime="00:04:54.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="23" reactiontime="+73" swimtime="00:03:11.65" resultid="2002" heatid="9074" lane="2" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="38" reactiontime="+129" swimtime="00:05:29.50" resultid="2003" heatid="9088" lane="4" entrytime="00:05:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.16" />
                    <SPLIT distance="100" swimtime="00:02:40.17" />
                    <SPLIT distance="150" swimtime="00:04:05.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="29" reactiontime="+192" swimtime="00:06:25.62" resultid="2004" heatid="9138" lane="2" entrytime="00:06:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.69" />
                    <SPLIT distance="100" swimtime="00:03:08.56" />
                    <SPLIT distance="150" swimtime="00:04:48.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="47" reactiontime="+160" swimtime="00:10:49.30" resultid="2005" heatid="9177" lane="5" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.25" />
                    <SPLIT distance="100" swimtime="00:02:30.62" />
                    <SPLIT distance="150" swimtime="00:03:52.08" />
                    <SPLIT distance="200" swimtime="00:05:16.40" />
                    <SPLIT distance="250" swimtime="00:06:38.25" />
                    <SPLIT distance="300" swimtime="00:08:00.61" />
                    <SPLIT distance="350" swimtime="00:09:24.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-21" firstname="Michał" gender="M" lastname="Kądzioła" nation="POL" athleteid="2015">
              <RESULTS>
                <RESULT eventid="1205" points="297" reactiontime="+63" swimtime="00:00:33.28" resultid="2016" heatid="8961" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1307" points="317" reactiontime="+89" swimtime="00:01:14.26" resultid="2017" heatid="9015" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="323" reactiontime="+88" swimtime="00:00:31.77" resultid="2018" heatid="9064" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1474" points="280" reactiontime="+71" swimtime="00:01:14.77" resultid="2019" heatid="9082" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="2020" heatid="9146" lane="0" entrytime="00:03:20.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="2021" heatid="9165" lane="8" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="1955">
              <RESULTS>
                <RESULT eventid="1079" points="84" reactiontime="+103" swimtime="00:00:46.09" resultid="1956" heatid="8896" lane="8" entrytime="00:00:45.25" />
                <RESULT eventid="1113" points="76" reactiontime="+102" swimtime="00:04:18.73" resultid="1957" heatid="8922" lane="9" entrytime="00:04:20.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.88" />
                    <SPLIT distance="100" swimtime="00:02:06.14" />
                    <SPLIT distance="150" swimtime="00:03:18.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="58" reactiontime="+69" swimtime="00:00:57.08" resultid="1958" heatid="8955" lane="3" entrytime="00:00:56.24" />
                <RESULT comment="Rekord Polski" eventid="1341" points="55" reactiontime="+91" swimtime="00:04:43.93" resultid="1959" heatid="9025" lane="3" entrytime="00:04:50.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.27" />
                    <SPLIT distance="100" swimtime="00:02:14.70" />
                    <SPLIT distance="150" swimtime="00:03:29.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="55" reactiontime="+100" swimtime="00:00:57.16" resultid="1960" heatid="9060" lane="2" entrytime="00:00:55.24" />
                <RESULT eventid="1578" points="71" reactiontime="+100" swimtime="00:09:26.37" resultid="1961" heatid="9116" lane="4" entrytime="00:09:40.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.48" />
                    <SPLIT distance="100" swimtime="00:02:16.19" />
                    <SPLIT distance="150" swimtime="00:03:30.03" />
                    <SPLIT distance="200" swimtime="00:04:43.99" />
                    <SPLIT distance="250" swimtime="00:05:59.31" />
                    <SPLIT distance="300" swimtime="00:07:14.91" />
                    <SPLIT distance="350" swimtime="00:08:21.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="50" reactiontime="+97" swimtime="00:02:11.37" resultid="1962" heatid="9129" lane="1" entrytime="00:02:06.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="100" reactiontime="+94" swimtime="00:00:54.26" resultid="1963" heatid="9160" lane="5" entrytime="00:00:55.09" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-12-07" firstname="Miron" gender="M" lastname="Starosta" nation="POL" athleteid="1989">
              <RESULTS>
                <RESULT eventid="1079" points="38" reactiontime="+104" swimtime="00:01:00.03" resultid="1990" heatid="8895" lane="4" entrytime="00:00:51.00" />
                <RESULT eventid="1239" points="72" reactiontime="+115" swimtime="00:04:49.38" resultid="1991" heatid="8971" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.54" />
                    <SPLIT distance="100" swimtime="00:02:23.77" />
                    <SPLIT distance="150" swimtime="00:03:37.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="63" reactiontime="+106" swimtime="00:01:52.55" resultid="1992" heatid="8985" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="65" reactiontime="+151" swimtime="00:02:18.25" resultid="1993" heatid="9043" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="52" reactiontime="+106" swimtime="00:04:25.50" resultid="1994" heatid="9095" lane="9" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.27" />
                    <SPLIT distance="100" swimtime="00:02:07.75" />
                    <SPLIT distance="150" swimtime="00:03:17.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="52" reactiontime="+123" swimtime="00:04:43.05" resultid="1995" heatid="9143" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.35" />
                    <SPLIT distance="100" swimtime="00:02:16.80" />
                    <SPLIT distance="150" swimtime="00:03:30.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="81" reactiontime="+105" swimtime="00:00:58.17" resultid="1996" heatid="9159" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-26" firstname="Władysław" gender="M" lastname="Szurek" nation="POL" athleteid="1982">
              <RESULTS>
                <RESULT eventid="1079" points="21" reactiontime="+108" swimtime="00:01:12.58" resultid="1983" heatid="8895" lane="8" entrytime="00:01:06.00" />
                <RESULT eventid="1205" points="13" reactiontime="+109" swimtime="00:01:33.98" resultid="1984" heatid="8954" lane="4" entrytime="00:01:23.00" />
                <RESULT eventid="1273" points="24" reactiontime="+115" swimtime="00:02:35.75" resultid="1985" heatid="8986" lane="8" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="16" reactiontime="+85" swimtime="00:03:12.70" resultid="1986" heatid="9079" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="18" reactiontime="+105" swimtime="00:06:14.94" resultid="1987" heatid="9094" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.24" />
                    <SPLIT distance="150" swimtime="00:04:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="16" reactiontime="+81" swimtime="00:06:55.65" resultid="1988" heatid="9142" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.98" />
                    <SPLIT distance="100" swimtime="00:03:18.90" />
                    <SPLIT distance="150" swimtime="00:05:07.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="2022" heatid="9109" lane="9">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1964" number="1" />
                    <RELAYPOSITION athleteid="1973" number="2" />
                    <RELAYPOSITION athleteid="2015" number="3" />
                    <RELAYPOSITION athleteid="2006" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="2023" heatid="9032" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1964" number="1" />
                    <RELAYPOSITION athleteid="1973" number="2" />
                    <RELAYPOSITION athleteid="2015" number="3" />
                    <RELAYPOSITION athleteid="2006" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SERLOD" nation="POL" region="LOD" clubid="3141" name="Sergiusz Olejniczak Team Łódź">
          <CONTACT city="Łódź" email="jblasiak@biol.uni.lodz.pl" name="Błasiak" phone="696033013" state="ŁÓDZK" street="Podchorążych 35A m 20" zip="94-234" />
          <ATHLETES>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" athleteid="3142">
              <RESULTS>
                <RESULT eventid="1079" points="326" reactiontime="+103" swimtime="00:00:29.41" resultid="3143" heatid="8897" lane="8" entrytime="00:00:40.18" />
                <RESULT eventid="1113" points="84" reactiontime="+110" swimtime="00:04:09.76" resultid="3144" heatid="8922" lane="0" entrytime="00:04:10.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.86" />
                    <SPLIT distance="100" swimtime="00:02:01.18" />
                    <SPLIT distance="150" swimtime="00:03:18.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="122" reactiontime="+100" swimtime="00:01:30.44" resultid="3145" heatid="8987" lane="2" entrytime="00:01:32.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="89" reactiontime="+103" swimtime="00:01:53.18" resultid="3146" heatid="9009" lane="2" entrytime="00:01:54.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="86" reactiontime="+84" swimtime="00:00:49.37" resultid="3147" heatid="9060" lane="3" entrytime="00:00:52.73" />
                <RESULT eventid="1508" points="90" reactiontime="+110" swimtime="00:03:41.01" resultid="3148" heatid="9095" lane="4" entrytime="00:03:30.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.08" />
                    <SPLIT distance="100" swimtime="00:01:48.23" />
                    <SPLIT distance="150" swimtime="00:02:49.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="57" reactiontime="+107" swimtime="00:04:35.18" resultid="3149" heatid="9144" lane="7" entrytime="00:04:27.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:03:28.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="89" reactiontime="+115" swimtime="00:07:54.43" resultid="3150" heatid="9183" lane="0" entrytime="00:07:45.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.75" />
                    <SPLIT distance="100" swimtime="00:01:53.74" />
                    <SPLIT distance="200" swimtime="00:03:55.96" />
                    <SPLIT distance="250" swimtime="00:04:57.44" />
                    <SPLIT distance="300" swimtime="00:05:58.49" />
                    <SPLIT distance="350" swimtime="00:07:00.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3183" name="SIKRET Gliwice">
          <CONTACT city="Gliwice" email="joannaeco@teln.pl" name="Zagała" phone="601427257" state="ŚLĄSK" street="Jagielońska 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1960-04-28" firstname="Marek" gender="M" lastname="Paściak" nation="POL" athleteid="3217">
              <RESULTS>
                <RESULT eventid="1079" points="144" reactiontime="+103" swimtime="00:00:38.61" resultid="3218" heatid="8897" lane="5" entrytime="00:00:39.50" />
                <RESULT eventid="1205" points="90" reactiontime="+110" swimtime="00:00:49.54" resultid="3219" heatid="8956" lane="2" entrytime="00:00:49.50" />
                <RESULT eventid="1273" points="129" reactiontime="+135" swimtime="00:01:28.72" resultid="3220" heatid="8988" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="103" reactiontime="+124" swimtime="00:01:44.37" resultid="3221" heatid="9080" lane="6" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="3222" heatid="9096" lane="8" entrytime="00:03:24.00" />
                <RESULT eventid="1744" points="123" reactiontime="+135" swimtime="00:07:06.12" resultid="3223" heatid="9183" lane="5" entrytime="00:07:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                    <SPLIT distance="100" swimtime="00:01:38.80" />
                    <SPLIT distance="150" swimtime="00:02:32.52" />
                    <SPLIT distance="200" swimtime="00:03:27.58" />
                    <SPLIT distance="250" swimtime="00:04:22.42" />
                    <SPLIT distance="300" swimtime="00:05:16.78" />
                    <SPLIT distance="350" swimtime="00:06:12.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-15" firstname="Mieczysław" gender="M" lastname="Mydłowski" nation="POL" athleteid="3230">
              <RESULTS>
                <RESULT eventid="1079" points="289" reactiontime="+98" swimtime="00:00:30.62" resultid="3231" heatid="8903" lane="6" entrytime="00:00:30.80" />
                <RESULT eventid="1205" points="189" reactiontime="+76" swimtime="00:00:38.66" resultid="3232" heatid="8959" lane="9" entrytime="00:00:38.00" />
                <RESULT eventid="1307" points="272" reactiontime="+95" swimtime="00:01:18.12" resultid="3233" heatid="9015" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K2 - Brak wynurzenia głowy po rozpoczęciu ruchu ramion do wewnątrz z jego najszerszego położenia w drugim cyklu ruchu ramion po starcie lub nawrocie (Time: 16:44)" eventid="1406" reactiontime="+91" status="DSQ" swimtime="00:01:29.05" resultid="3234" heatid="9051" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="187" reactiontime="+76" swimtime="00:01:25.49" resultid="3235" heatid="9082" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-10-21" firstname="Krystian" gender="M" lastname="Kapias" nation="POL" athleteid="3236">
              <RESULTS>
                <RESULT eventid="1079" points="180" reactiontime="+88" swimtime="00:00:35.83" resultid="3237" heatid="8900" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1273" points="145" reactiontime="+89" swimtime="00:01:25.51" resultid="3238" heatid="8989" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-14" firstname="Dawid" gender="M" lastname="Zimkowski" nation="POL" athleteid="3208">
              <RESULTS>
                <RESULT eventid="1079" points="313" reactiontime="+86" swimtime="00:00:29.81" resultid="3209" heatid="8904" lane="1" entrytime="00:00:30.26" />
                <RESULT eventid="1205" points="257" reactiontime="+78" swimtime="00:00:34.91" resultid="3210" heatid="8960" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1440" points="293" reactiontime="+82" swimtime="00:00:32.82" resultid="3211" heatid="9066" lane="6" entrytime="00:00:32.50" />
                <RESULT eventid="1474" points="223" reactiontime="+81" swimtime="00:01:20.64" resultid="3212" heatid="9082" lane="0" entrytime="00:01:26.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="225" reactiontime="+100" swimtime="00:05:48.90" resultid="3213" heatid="9185" lane="2" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:19.64" />
                    <SPLIT distance="150" swimtime="00:02:04.94" />
                    <SPLIT distance="200" swimtime="00:02:50.29" />
                    <SPLIT distance="250" swimtime="00:03:35.12" />
                    <SPLIT distance="300" swimtime="00:04:20.17" />
                    <SPLIT distance="350" swimtime="00:05:05.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-11" firstname="Agnieszka" gender="F" lastname="Drejka" nation="POL" athleteid="3201">
              <RESULTS>
                <RESULT eventid="1062" points="194" reactiontime="+95" swimtime="00:00:40.11" resultid="3202" heatid="8887" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1222" points="181" reactiontime="+107" swimtime="00:03:57.84" resultid="3203" heatid="8968" lane="8" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.98" />
                    <SPLIT distance="100" swimtime="00:01:50.29" />
                    <SPLIT distance="150" swimtime="00:02:54.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="160" reactiontime="+102" swimtime="00:01:33.79" resultid="3204" heatid="8980" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="181" reactiontime="+95" swimtime="00:01:50.11" resultid="3205" heatid="9039" lane="8" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="149" reactiontime="+103" swimtime="00:03:28.50" resultid="3206" heatid="9089" lane="4" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.34" />
                    <SPLIT distance="100" swimtime="00:01:37.11" />
                    <SPLIT distance="150" swimtime="00:02:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="185" reactiontime="+101" swimtime="00:00:50.52" resultid="3207" heatid="9154" lane="0" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-10-06" firstname="Arkadiusz" gender="M" lastname="Bednarek" nation="POL" athleteid="3224">
              <RESULTS>
                <RESULT eventid="1079" points="191" reactiontime="+80" swimtime="00:00:35.15" resultid="3225" heatid="8899" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1273" points="201" reactiontime="+80" swimtime="00:01:16.63" resultid="3226" heatid="8988" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="178" reactiontime="+91" swimtime="00:00:38.69" resultid="3227" heatid="9065" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1508" points="151" reactiontime="+89" swimtime="00:03:06.22" resultid="3228" heatid="9097" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:26.59" />
                    <SPLIT distance="150" swimtime="00:02:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="142" reactiontime="+89" swimtime="00:06:46.41" resultid="3229" heatid="9184" lane="4" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:01:29.75" />
                    <SPLIT distance="150" swimtime="00:02:20.86" />
                    <SPLIT distance="200" swimtime="00:03:13.10" />
                    <SPLIT distance="250" swimtime="00:04:06.36" />
                    <SPLIT distance="300" swimtime="00:04:59.12" />
                    <SPLIT distance="350" swimtime="00:05:53.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="3192">
              <RESULTS>
                <RESULT eventid="1062" points="238" reactiontime="+76" swimtime="00:00:37.48" resultid="3193" heatid="8888" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="3194" heatid="8937" lane="9" entrytime="00:15:30.00" />
                <RESULT eventid="1256" points="220" reactiontime="+78" swimtime="00:01:24.41" resultid="3195" heatid="8979" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="189" reactiontime="+82" swimtime="00:01:38.68" resultid="3196" heatid="9002" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="168" reactiontime="+82" swimtime="00:01:39.69" resultid="3197" heatid="9075" lane="0" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="189" reactiontime="+83" swimtime="00:03:12.91" resultid="3198" heatid="9089" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.44" />
                    <SPLIT distance="100" swimtime="00:01:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="200" reactiontime="+77" swimtime="00:00:49.19" resultid="3199" heatid="9152" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1721" points="178" reactiontime="+83" swimtime="00:06:56.26" resultid="3200" heatid="9178" lane="8" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                    <SPLIT distance="100" swimtime="00:01:37.28" />
                    <SPLIT distance="350" swimtime="00:06:08.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-03-14" firstname="Tomasz" gender="M" lastname="Bartosik" nation="POL" athleteid="3214">
              <RESULTS>
                <RESULT eventid="1079" points="394" reactiontime="+81" swimtime="00:00:27.63" resultid="3215" heatid="8909" lane="1" entrytime="00:00:27.98" />
                <RESULT eventid="1273" points="375" reactiontime="+77" swimtime="00:01:02.31" resultid="3216" heatid="8995" lane="9" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="3184">
              <RESULTS>
                <RESULT eventid="1062" points="209" reactiontime="+95" swimtime="00:00:39.14" resultid="3185" heatid="8887" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1222" points="197" reactiontime="+86" swimtime="00:03:51.25" resultid="3186" heatid="8967" lane="5" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.88" />
                    <SPLIT distance="100" swimtime="00:01:52.58" />
                    <SPLIT distance="150" swimtime="00:02:54.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="91" reactiontime="+101" swimtime="00:04:25.00" resultid="3187" heatid="9023" lane="1" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.68" />
                    <SPLIT distance="100" swimtime="00:02:05.48" />
                    <SPLIT distance="150" swimtime="00:03:15.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="204" reactiontime="+85" swimtime="00:01:45.93" resultid="3188" heatid="9038" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="139" reactiontime="+85" swimtime="00:08:21.05" resultid="3189" heatid="9113" lane="5" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.81" />
                    <SPLIT distance="100" swimtime="00:02:02.11" />
                    <SPLIT distance="150" swimtime="00:03:16.40" />
                    <SPLIT distance="200" swimtime="00:04:26.99" />
                    <SPLIT distance="250" swimtime="00:05:28.03" />
                    <SPLIT distance="300" swimtime="00:06:28.36" />
                    <SPLIT distance="350" swimtime="00:07:27.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="101" reactiontime="+90" swimtime="00:01:56.92" resultid="3190" heatid="9124" lane="7" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="233" reactiontime="+85" swimtime="00:00:46.74" resultid="3191" heatid="9154" lane="1" entrytime="00:00:48.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-29" firstname="Szymon" gender="M" lastname="Chrzanowski" nation="POL" athleteid="3252">
              <RESULTS>
                <RESULT eventid="1079" points="292" reactiontime="+70" swimtime="00:00:30.53" resultid="3253" heatid="8906" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1205" points="199" reactiontime="+55" swimtime="00:00:38.00" resultid="3254" heatid="8960" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1406" points="283" reactiontime="+75" swimtime="00:01:24.66" resultid="3255" heatid="9052" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="209" reactiontime="+69" swimtime="00:00:36.73" resultid="3256" heatid="9066" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1681" points="305" reactiontime="+71" swimtime="00:00:37.48" resultid="3257" heatid="9169" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="3258" heatid="9190" lane="9" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="308" reactiontime="+97" swimtime="00:02:02.19" resultid="3239" heatid="9110" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:05.96" />
                    <SPLIT distance="150" swimtime="00:01:34.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3230" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="3236" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="3208" number="3" reactiontime="+5" />
                    <RELAYPOSITION athleteid="3214" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="258" reactiontime="+79" swimtime="00:02:22.12" resultid="3240" heatid="9033" lane="0" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:54.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3208" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="3230" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="3224" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3214" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="229" reactiontime="+84" swimtime="00:02:14.92" resultid="3241" heatid="8934" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:17.23" />
                    <SPLIT distance="150" swimtime="00:01:47.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3184" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3192" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3230" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3214" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="187" reactiontime="+78" swimtime="00:02:38.02" resultid="3242" heatid="9174" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.19" />
                    <SPLIT distance="100" swimtime="00:01:33.54" />
                    <SPLIT distance="150" swimtime="00:02:10.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3192" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3184" number="2" reactiontime="+74" />
                    <RELAYPOSITION athleteid="3230" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3214" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="2238" name="SK Spolchemie Usti nad Labem">
          <CONTACT email="benova.dana@seznam.cz" name="SK Spolchemie Usti nad Labem" />
          <ATHLETES>
            <ATHLETE birthdate="1956-07-10" firstname="Vaclav" gender="M" lastname="Valtr" nation="CZE" athleteid="2248" />
            <ATHLETE birthdate="1956-01-26" firstname="Dana" gender="F" lastname="Benova" nation="CZE" athleteid="2239">
              <RESULTS>
                <RESULT eventid="1096" points="87" reactiontime="+87" swimtime="00:04:34.21" resultid="2240" heatid="8916" lane="2" entrytime="00:09:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.15" />
                    <SPLIT distance="100" swimtime="00:02:17.27" />
                    <SPLIT distance="150" swimtime="00:03:28.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="93" reactiontime="+102" swimtime="00:17:37.30" resultid="2241" heatid="8936" lane="3" entrytime="00:17:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.93" />
                    <SPLIT distance="100" swimtime="00:02:01.69" />
                    <SPLIT distance="150" swimtime="00:03:07.71" />
                    <SPLIT distance="200" swimtime="00:04:13.75" />
                    <SPLIT distance="250" swimtime="00:05:19.46" />
                    <SPLIT distance="300" swimtime="00:06:26.55" />
                    <SPLIT distance="350" swimtime="00:07:33.78" />
                    <SPLIT distance="400" swimtime="00:08:41.40" />
                    <SPLIT distance="450" swimtime="00:09:49.49" />
                    <SPLIT distance="500" swimtime="00:10:57.89" />
                    <SPLIT distance="550" swimtime="00:12:05.34" />
                    <SPLIT distance="600" swimtime="00:13:12.93" />
                    <SPLIT distance="650" swimtime="00:14:20.54" />
                    <SPLIT distance="700" swimtime="00:15:26.59" />
                    <SPLIT distance="750" swimtime="00:16:33.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="99" reactiontime="+93" swimtime="00:04:50.70" resultid="2242" heatid="8967" lane="7" entrytime="00:04:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.58" />
                    <SPLIT distance="100" swimtime="00:02:20.47" />
                    <SPLIT distance="150" swimtime="00:03:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="30" reactiontime="+98" swimtime="00:06:21.12" resultid="2243" heatid="9023" lane="0" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.21" />
                    <SPLIT distance="100" swimtime="00:03:01.85" />
                    <SPLIT distance="150" swimtime="00:04:44.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="83" reactiontime="+96" swimtime="00:04:13.78" resultid="2244" heatid="9089" lane="0" entrytime="00:04:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.30" />
                    <SPLIT distance="100" swimtime="00:02:02.29" />
                    <SPLIT distance="150" swimtime="00:03:10.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="82" reactiontime="+92" swimtime="00:09:57.37" resultid="2245" heatid="9113" lane="7" entrytime="00:09:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.46" />
                    <SPLIT distance="100" swimtime="00:04:08.98" />
                    <SPLIT distance="150" swimtime="00:05:17.74" />
                    <SPLIT distance="200" swimtime="00:06:32.32" />
                    <SPLIT distance="250" swimtime="00:07:44.88" />
                    <SPLIT distance="350" swimtime="00:08:53.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="84" reactiontime="+82" swimtime="00:04:32.18" resultid="2246" heatid="9138" lane="4" entrytime="00:04:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.92" />
                    <SPLIT distance="100" swimtime="00:02:13.04" />
                    <SPLIT distance="150" swimtime="00:03:24.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="88" swimtime="00:08:46.62" resultid="2247" heatid="9178" lane="9" entrytime="00:08:49.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.26" />
                    <SPLIT distance="100" swimtime="00:02:03.11" />
                    <SPLIT distance="150" swimtime="00:03:12.04" />
                    <SPLIT distance="200" swimtime="00:04:19.33" />
                    <SPLIT distance="250" swimtime="00:05:27.04" />
                    <SPLIT distance="300" swimtime="00:06:33.99" />
                    <SPLIT distance="350" swimtime="00:07:41.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4079" name="SMT Szczecin">
          <CONTACT city="Szczecin" email="aga.krzyzostaniak@gmail.com" name="Krzyżostaniak" phone="603772862" street="Szafera 110/1" zip="71-245" />
          <ATHLETES>
            <ATHLETE birthdate="1984-03-20" firstname="Marcin" gender="M" lastname="Łogin" nation="POL" athleteid="7058">
              <RESULTS>
                <RESULT eventid="1079" points="298" reactiontime="+83" swimtime="00:00:30.33" resultid="7059" heatid="8905" lane="9" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="7060" heatid="8976" lane="1" entrytime="00:03:05.00" entrycourse="SCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="7061" heatid="9051" lane="3" entrytime="00:01:18.23" entrycourse="SCM" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="7062" heatid="9169" lane="2" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="Roenig" nation="POL" athleteid="7023">
              <RESULTS>
                <RESULT eventid="1113" points="356" reactiontime="+103" swimtime="00:02:34.56" resultid="7024" heatid="8931" lane="2" entrytime="00:02:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:09.83" />
                    <SPLIT distance="150" swimtime="00:01:54.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="7025" heatid="8977" lane="4" entrytime="00:02:45.00" entrycourse="SCM" />
                <RESULT eventid="1307" points="390" reactiontime="+95" swimtime="00:01:09.28" resultid="7026" heatid="9016" lane="1" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="394" reactiontime="+94" swimtime="00:01:15.80" resultid="7027" heatid="9052" lane="8" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="413" reactiontime="+86" swimtime="00:00:33.89" resultid="7028" heatid="9171" lane="8" entrytime="00:00:34.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-12" firstname="Kamila" gender="F" lastname="Gębka" nation="POL" athleteid="7002">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="7003" heatid="8919" lane="4" entrytime="00:02:55.00" entrycourse="SCM" />
                <RESULT eventid="1222" points="305" reactiontime="+97" swimtime="00:03:19.75" resultid="7004" heatid="8970" lane="7" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                    <SPLIT distance="100" swimtime="00:01:35.63" />
                    <SPLIT distance="150" swimtime="00:02:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="7005" heatid="9024" lane="0" entrytime="00:03:20.00" entrycourse="SCM" />
                <RESULT eventid="1388" points="283" reactiontime="+93" swimtime="00:01:34.88" resultid="7006" heatid="9041" lane="8" entrytime="00:01:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" status="DNS" swimtime="00:00:00.00" resultid="7007" heatid="9115" lane="9" entrytime="00:06:20.00" entrycourse="SCM" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="7008" heatid="9126" lane="8" entrytime="00:01:25.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-14" firstname="Kinga" gender="F" lastname="Maciupa" nation="POL" athleteid="7015">
              <RESULTS>
                <RESULT eventid="1062" points="412" reactiontime="+81" swimtime="00:00:31.21" resultid="7016" heatid="8893" lane="0" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1096" points="424" reactiontime="+76" swimtime="00:02:42.12" resultid="7017" heatid="8920" lane="8" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                    <SPLIT distance="150" swimtime="00:02:02.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="461" reactiontime="+66" swimtime="00:00:33.21" resultid="7018" heatid="8952" lane="6" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1290" points="435" reactiontime="+79" swimtime="00:01:14.81" resultid="7019" heatid="9006" lane="4" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="407" reactiontime="+73" swimtime="00:00:32.89" resultid="7020" heatid="9059" lane="9" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1555" points="454" reactiontime="+82" swimtime="00:05:37.86" resultid="7021" heatid="9115" lane="5" entrytime="00:05:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="150" swimtime="00:01:59.69" />
                    <SPLIT distance="200" swimtime="00:02:42.27" />
                    <SPLIT distance="250" swimtime="00:03:31.06" />
                    <SPLIT distance="300" swimtime="00:04:20.15" />
                    <SPLIT distance="350" swimtime="00:05:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="409" reactiontime="+77" swimtime="00:01:13.51" resultid="7022" heatid="9127" lane="1" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-20" firstname="Agnieszka" gender="F" lastname="Krzyżostaniak" nation="POL" athleteid="7051">
              <RESULTS>
                <RESULT eventid="1062" points="563" reactiontime="+74" swimtime="00:00:28.13" resultid="7052" heatid="8892" lane="5" entrytime="00:00:29.50" entrycourse="SCM" />
                <RESULT eventid="1147" points="537" reactiontime="+79" swimtime="00:09:49.68" resultid="7053" heatid="8939" lane="4" entrytime="00:10:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:07.37" />
                    <SPLIT distance="150" swimtime="00:01:43.48" />
                    <SPLIT distance="200" swimtime="00:02:20.66" />
                    <SPLIT distance="250" swimtime="00:02:57.98" />
                    <SPLIT distance="300" swimtime="00:03:35.34" />
                    <SPLIT distance="350" swimtime="00:04:13.02" />
                    <SPLIT distance="400" swimtime="00:04:50.14" />
                    <SPLIT distance="450" swimtime="00:05:27.40" />
                    <SPLIT distance="500" swimtime="00:06:04.68" />
                    <SPLIT distance="550" swimtime="00:06:42.36" />
                    <SPLIT distance="600" swimtime="00:07:20.13" />
                    <SPLIT distance="650" swimtime="00:07:57.88" />
                    <SPLIT distance="700" swimtime="00:08:36.06" />
                    <SPLIT distance="750" swimtime="00:09:13.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="588" reactiontime="+72" swimtime="00:00:30.63" resultid="7054" heatid="8953" lane="1" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1290" points="548" reactiontime="+83" swimtime="00:01:09.26" resultid="7055" heatid="9007" lane="0" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="506" reactiontime="+79" swimtime="00:05:25.97" resultid="7056" heatid="9115" lane="4" entrytime="00:05:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="150" swimtime="00:01:57.31" />
                    <SPLIT distance="200" swimtime="00:02:37.74" />
                    <SPLIT distance="250" swimtime="00:03:26.20" />
                    <SPLIT distance="300" swimtime="00:04:14.51" />
                    <SPLIT distance="350" swimtime="00:04:51.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="555" reactiontime="+78" swimtime="00:04:45.25" resultid="7057" heatid="9181" lane="3" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="150" swimtime="00:01:42.77" />
                    <SPLIT distance="200" swimtime="00:02:19.62" />
                    <SPLIT distance="250" swimtime="00:02:56.27" />
                    <SPLIT distance="300" swimtime="00:03:33.85" />
                    <SPLIT distance="350" swimtime="00:04:10.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-09" firstname="Helena" gender="F" lastname="Szulc" nation="POL" athleteid="7009">
              <RESULTS>
                <RESULT eventid="1096" points="326" reactiontime="+80" swimtime="00:02:56.93" resultid="7010" heatid="8920" lane="9" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:21.71" />
                    <SPLIT distance="150" swimtime="00:02:14.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="351" reactiontime="+96" swimtime="00:01:20.31" resultid="7011" heatid="9005" lane="1" entrytime="00:01:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="216" reactiontime="+98" swimtime="00:03:19.06" resultid="7012" heatid="9024" lane="8" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                    <SPLIT distance="100" swimtime="00:01:36.64" />
                    <SPLIT distance="150" swimtime="00:02:28.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="319" reactiontime="+93" swimtime="00:06:19.97" resultid="7013" heatid="9115" lane="0" entrytime="00:06:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:32.95" />
                    <SPLIT distance="150" swimtime="00:02:20.08" />
                    <SPLIT distance="200" swimtime="00:03:06.15" />
                    <SPLIT distance="250" swimtime="00:03:59.05" />
                    <SPLIT distance="300" swimtime="00:04:52.68" />
                    <SPLIT distance="350" swimtime="00:05:37.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="7014" heatid="9126" lane="9" entrytime="00:01:26.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-21" firstname="Michał" gender="M" lastname="Krysiak" nation="POL" athleteid="7037">
              <RESULTS>
                <RESULT eventid="1079" points="455" reactiontime="+78" swimtime="00:00:26.34" resultid="7038" heatid="8912" lane="9" entrytime="00:00:26.50" entrycourse="SCM" />
                <RESULT eventid="1113" points="335" reactiontime="+79" swimtime="00:02:37.71" resultid="7039" heatid="8928" lane="9" entrytime="00:02:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:02:03.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="464" reactiontime="+80" swimtime="00:00:58.04" resultid="7040" heatid="8997" lane="4" entrytime="00:01:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="392" reactiontime="+82" swimtime="00:02:28.30" resultid="7041" heatid="9030" lane="1" entrytime="00:02:33.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="100" swimtime="00:01:10.76" />
                    <SPLIT distance="150" swimtime="00:01:50.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="430" reactiontime="+83" swimtime="00:00:28.88" resultid="7042" heatid="9070" lane="1" entrytime="00:00:29.15" entrycourse="SCM" />
                <RESULT eventid="1508" points="345" reactiontime="+83" swimtime="00:02:21.60" resultid="7043" heatid="9102" lane="8" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:01:48.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="451" reactiontime="+82" swimtime="00:01:03.12" resultid="7044" heatid="9135" lane="5" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="332" reactiontime="+81" swimtime="00:05:06.29" resultid="7045" heatid="9189" lane="3" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:15.21" />
                    <SPLIT distance="150" swimtime="00:01:55.48" />
                    <SPLIT distance="200" swimtime="00:02:35.87" />
                    <SPLIT distance="250" swimtime="00:03:16.03" />
                    <SPLIT distance="300" swimtime="00:03:54.95" />
                    <SPLIT distance="350" swimtime="00:04:31.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-07-21" firstname="Wiktoria" gender="F" lastname="Podkowińska" nation="POL" athleteid="7029">
              <RESULTS>
                <RESULT eventid="1062" points="351" reactiontime="+78" swimtime="00:00:32.94" resultid="7030" heatid="8891" lane="7" entrytime="00:00:31.25" entrycourse="SCM" />
                <RESULT eventid="1096" points="319" reactiontime="+74" swimtime="00:02:58.22" resultid="7031" heatid="8919" lane="5" entrytime="00:02:56.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:27.03" />
                    <SPLIT distance="150" swimtime="00:02:18.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="321" reactiontime="+79" swimtime="00:01:22.74" resultid="7032" heatid="9005" lane="2" entrytime="00:01:22.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="275" reactiontime="+79" swimtime="00:00:37.46" resultid="7033" heatid="9057" lane="4" entrytime="00:00:34.87" entrycourse="SCM" />
                <RESULT eventid="1555" points="325" reactiontime="+86" swimtime="00:06:17.64" resultid="7034" heatid="9115" lane="3" entrytime="00:05:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:29.77" />
                    <SPLIT distance="150" swimtime="00:02:21.29" />
                    <SPLIT distance="200" swimtime="00:03:10.46" />
                    <SPLIT distance="250" swimtime="00:04:02.42" />
                    <SPLIT distance="300" swimtime="00:04:55.60" />
                    <SPLIT distance="350" swimtime="00:05:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="257" reactiontime="+83" swimtime="00:01:25.85" resultid="7035" heatid="9126" lane="1" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="286" reactiontime="+83" swimtime="00:00:43.71" resultid="7036" heatid="9157" lane="0" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-12" firstname="Marek" gender="M" lastname="Zienkiewicz" nation="POL" athleteid="7046">
              <RESULTS>
                <RESULT eventid="1079" points="292" reactiontime="+76" swimtime="00:00:30.53" resultid="7047" heatid="8903" lane="3" entrytime="00:00:30.78" entrycourse="SCM" />
                <RESULT eventid="1307" points="212" reactiontime="+73" swimtime="00:01:24.94" resultid="7048" heatid="9012" lane="9" entrytime="00:01:26.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="241" reactiontime="+80" swimtime="00:01:29.24" resultid="7049" heatid="9047" lane="2" entrytime="00:01:30.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="262" reactiontime="+77" swimtime="00:00:39.42" resultid="7050" heatid="9164" lane="3" entrytime="00:00:40.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="7067" heatid="9034" lane="8" entrytime="00:02:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7046" number="1" />
                    <RELAYPOSITION athleteid="7058" number="2" />
                    <RELAYPOSITION athleteid="7037" number="3" />
                    <RELAYPOSITION athleteid="7023" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="7068" heatid="9110" lane="9" entrytime="00:02:12.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7023" number="1" />
                    <RELAYPOSITION athleteid="7046" number="2" />
                    <RELAYPOSITION athleteid="7058" number="3" />
                    <RELAYPOSITION athleteid="7037" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="297" reactiontime="+87" swimtime="00:02:03.78" resultid="7065" heatid="8933" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:03.69" />
                    <SPLIT distance="150" swimtime="00:01:37.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7002" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="7046" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="7009" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="7037" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="251" reactiontime="+73" swimtime="00:02:23.37" resultid="7066" heatid="9175" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                    <SPLIT distance="150" swimtime="00:01:55.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7002" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="7023" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="7009" number="3" />
                    <RELAYPOSITION athleteid="7046" number="4" reactiontime="+96" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="SMT Szczecin 2" number="1">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="7069" heatid="8933" lane="7" entrytime="00:02:25.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7023" number="1" />
                    <RELAYPOSITION athleteid="7015" number="2" />
                    <RELAYPOSITION athleteid="7029" number="3" />
                    <RELAYPOSITION athleteid="7058" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="7070" heatid="9175" lane="4" entrytime="00:02:15.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7051" number="1" />
                    <RELAYPOSITION athleteid="7058" number="2" />
                    <RELAYPOSITION athleteid="7015" number="3" />
                    <RELAYPOSITION athleteid="7037" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4804" name="Start Poznań">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" street="os. Batorego 8/67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1987-06-06" firstname="Joanna" gender="F" lastname="Kostencka" nation="POL" athleteid="4841">
              <RESULTS>
                <RESULT eventid="1096" points="373" reactiontime="+87" swimtime="00:02:49.28" resultid="4842" heatid="8919" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                    <SPLIT distance="100" swimtime="00:01:17.98" />
                    <SPLIT distance="150" swimtime="00:02:09.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="349" reactiontime="+89" swimtime="00:11:20.64" resultid="4843" heatid="8938" lane="4" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:01:18.66" />
                    <SPLIT distance="150" swimtime="00:02:00.35" />
                    <SPLIT distance="200" swimtime="00:02:42.56" />
                    <SPLIT distance="250" swimtime="00:03:24.93" />
                    <SPLIT distance="300" swimtime="00:04:08.06" />
                    <SPLIT distance="350" swimtime="00:04:50.99" />
                    <SPLIT distance="400" swimtime="00:05:34.20" />
                    <SPLIT distance="450" swimtime="00:06:17.68" />
                    <SPLIT distance="500" swimtime="00:07:01.45" />
                    <SPLIT distance="550" swimtime="00:07:45.76" />
                    <SPLIT distance="600" swimtime="00:08:29.43" />
                    <SPLIT distance="650" swimtime="00:09:12.40" />
                    <SPLIT distance="700" swimtime="00:09:55.42" />
                    <SPLIT distance="750" swimtime="00:10:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="353" reactiontime="+77" swimtime="00:00:36.30" resultid="4844" heatid="8952" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1290" points="356" reactiontime="+87" swimtime="00:01:19.99" resultid="4845" heatid="9005" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="365" reactiontime="+77" swimtime="00:01:16.99" resultid="4846" heatid="9078" lane="9" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="388" reactiontime="+81" swimtime="00:02:43.42" resultid="4847" heatid="9141" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:01:19.56" />
                    <SPLIT distance="150" swimtime="00:02:01.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="375" reactiontime="+88" swimtime="00:05:25.18" resultid="4848" heatid="9180" lane="5" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                    <SPLIT distance="100" swimtime="00:01:18.77" />
                    <SPLIT distance="150" swimtime="00:01:59.45" />
                    <SPLIT distance="200" swimtime="00:02:40.62" />
                    <SPLIT distance="250" swimtime="00:03:21.75" />
                    <SPLIT distance="300" swimtime="00:04:03.46" />
                    <SPLIT distance="350" swimtime="00:04:44.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-06-06" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="4818">
              <RESULTS>
                <RESULT eventid="1079" points="446" reactiontime="+71" swimtime="00:00:26.50" resultid="4819" heatid="8912" lane="2" entrytime="00:00:26.40" />
                <RESULT eventid="1113" points="401" reactiontime="+79" swimtime="00:02:28.62" resultid="4820" heatid="8930" lane="8" entrytime="00:02:27.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="100" swimtime="00:01:11.70" />
                    <SPLIT distance="150" swimtime="00:01:55.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="480" reactiontime="+75" swimtime="00:00:57.39" resultid="4821" heatid="8999" lane="6" entrytime="00:00:57.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="418" reactiontime="+76" swimtime="00:01:07.74" resultid="4822" heatid="9019" lane="7" entrytime="00:01:07.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="470" reactiontime="+79" swimtime="00:02:07.75" resultid="4823" heatid="9104" lane="4" entrytime="00:02:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:04.33" />
                    <SPLIT distance="150" swimtime="00:01:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="390" reactiontime="+70" swimtime="00:05:22.22" resultid="4824" heatid="9121" lane="3" entrytime="00:05:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:13.23" />
                    <SPLIT distance="150" swimtime="00:01:55.58" />
                    <SPLIT distance="200" swimtime="00:02:37.67" />
                    <SPLIT distance="250" swimtime="00:03:24.29" />
                    <SPLIT distance="300" swimtime="00:04:12.00" />
                    <SPLIT distance="350" swimtime="00:04:48.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="450" reactiontime="+77" swimtime="00:04:36.78" resultid="4825" heatid="9191" lane="4" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:07.66" />
                    <SPLIT distance="150" swimtime="00:01:43.33" />
                    <SPLIT distance="200" swimtime="00:02:19.25" />
                    <SPLIT distance="250" swimtime="00:02:53.97" />
                    <SPLIT distance="300" swimtime="00:03:28.80" />
                    <SPLIT distance="350" swimtime="00:04:03.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-06" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="4826">
              <RESULTS>
                <RESULT eventid="1079" points="475" reactiontime="+72" swimtime="00:00:25.96" resultid="4827" heatid="8908" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="4828" heatid="8928" lane="2" entrytime="00:02:40.00" />
                <RESULT eventid="1205" points="392" reactiontime="+78" swimtime="00:00:30.36" resultid="4829" heatid="8961" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1307" points="478" reactiontime="+73" swimtime="00:01:04.78" resultid="4830" heatid="9018" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="434" reactiontime="+72" swimtime="00:01:04.63" resultid="4831" heatid="9085" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="4832" heatid="9134" lane="0" entrytime="00:01:10.00" />
                <RESULT eventid="1647" points="421" reactiontime="+70" swimtime="00:02:21.56" resultid="4833" heatid="9148" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                    <SPLIT distance="100" swimtime="00:01:08.50" />
                    <SPLIT distance="150" swimtime="00:01:44.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-06-06" firstname="Anna" gender="F" lastname="Rostkowska-Kaczmarek" nation="POL" athleteid="4849">
              <RESULTS>
                <RESULT eventid="1062" points="294" reactiontime="+94" swimtime="00:00:34.95" resultid="4850" heatid="8889" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1147" points="164" reactiontime="+99" swimtime="00:14:34.42" resultid="4851" heatid="8937" lane="1" entrytime="00:14:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                    <SPLIT distance="100" swimtime="00:01:34.66" />
                    <SPLIT distance="150" swimtime="00:02:28.40" />
                    <SPLIT distance="200" swimtime="00:03:24.51" />
                    <SPLIT distance="250" swimtime="00:04:20.22" />
                    <SPLIT distance="300" swimtime="00:05:17.50" />
                    <SPLIT distance="350" swimtime="00:06:14.24" />
                    <SPLIT distance="400" swimtime="00:07:11.38" />
                    <SPLIT distance="450" swimtime="00:08:07.92" />
                    <SPLIT distance="500" swimtime="00:10:01.15" />
                    <SPLIT distance="550" swimtime="00:10:56.31" />
                    <SPLIT distance="600" swimtime="00:11:51.55" />
                    <SPLIT distance="650" swimtime="00:12:47.06" />
                    <SPLIT distance="750" swimtime="00:13:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="239" reactiontime="+83" swimtime="00:01:22.14" resultid="4852" heatid="8980" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="205" reactiontime="+97" swimtime="00:01:36.15" resultid="4853" heatid="9003" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="173" reactiontime="+100" swimtime="00:00:43.72" resultid="4854" heatid="9056" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1664" points="236" reactiontime="+101" swimtime="00:00:46.55" resultid="4855" heatid="9154" lane="6" entrytime="00:00:47.50" />
                <RESULT eventid="1721" points="169" reactiontime="+100" swimtime="00:07:04.09" resultid="4856" heatid="9179" lane="1" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.48" />
                    <SPLIT distance="150" swimtime="00:02:33.86" />
                    <SPLIT distance="200" swimtime="00:03:28.79" />
                    <SPLIT distance="300" swimtime="00:05:17.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-06" firstname="Mikołaj" gender="M" lastname="Osuch" nation="POL" athleteid="4834">
              <RESULTS>
                <RESULT eventid="1079" points="540" reactiontime="+75" swimtime="00:00:24.87" resultid="4835" heatid="8914" lane="5" entrytime="00:00:24.50" />
                <RESULT eventid="1205" points="502" reactiontime="+62" swimtime="00:00:27.94" resultid="4836" heatid="8964" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1307" points="539" reactiontime="+78" swimtime="00:01:02.22" resultid="4837" heatid="9020" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="549" reactiontime="+57" swimtime="00:00:59.74" resultid="4838" heatid="9087" lane="7" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="500" reactiontime="+65" swimtime="00:02:13.67" resultid="4839" heatid="9150" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                    <SPLIT distance="100" swimtime="00:01:05.19" />
                    <SPLIT distance="150" swimtime="00:01:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="448" reactiontime="+78" swimtime="00:00:32.98" resultid="4840" heatid="9171" lane="3" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-06" firstname="Aneta" gender="F" lastname="Maduzia" nation="POL" athleteid="4811">
              <RESULTS>
                <RESULT eventid="1062" points="357" reactiontime="+93" swimtime="00:00:32.76" resultid="4812" heatid="8889" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1147" points="279" reactiontime="+92" swimtime="00:12:12.73" resultid="4813" heatid="8938" lane="8" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="150" swimtime="00:02:07.15" />
                    <SPLIT distance="200" swimtime="00:02:53.25" />
                    <SPLIT distance="250" swimtime="00:03:39.53" />
                    <SPLIT distance="300" swimtime="00:04:25.79" />
                    <SPLIT distance="450" swimtime="00:08:21.55" />
                    <SPLIT distance="700" swimtime="00:11:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="344" reactiontime="+85" swimtime="00:01:12.74" resultid="4814" heatid="8981" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="269" reactiontime="+89" swimtime="00:01:36.50" resultid="4815" heatid="9039" lane="6" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="325" reactiontime="+94" swimtime="00:02:41.12" resultid="4816" heatid="9091" lane="7" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                    <SPLIT distance="150" swimtime="00:02:01.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="316" reactiontime="+93" swimtime="00:05:44.10" resultid="4817" heatid="9180" lane="8" entrytime="00:06:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                    <SPLIT distance="150" swimtime="00:02:08.42" />
                    <SPLIT distance="200" swimtime="00:02:52.24" />
                    <SPLIT distance="250" swimtime="00:03:35.54" />
                    <SPLIT distance="300" swimtime="00:04:19.79" />
                    <SPLIT distance="350" swimtime="00:05:03.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-06-06" firstname="Krzysztof" gender="M" lastname="Kapałczyński" nation="POL" athleteid="4805">
              <RESULTS>
                <RESULT eventid="1113" points="265" reactiontime="+94" swimtime="00:02:50.57" resultid="4806" heatid="8927" lane="1" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:19.75" />
                    <SPLIT distance="150" swimtime="00:02:11.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="207" reactiontime="+93" swimtime="00:03:03.48" resultid="4807" heatid="9028" lane="4" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:22.87" />
                    <SPLIT distance="150" swimtime="00:02:12.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="307" reactiontime="+88" swimtime="00:01:22.41" resultid="4808" heatid="9050" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="278" reactiontime="+91" swimtime="00:06:00.72" resultid="4809" heatid="9120" lane="6" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="150" swimtime="00:02:05.82" />
                    <SPLIT distance="200" swimtime="00:02:51.58" />
                    <SPLIT distance="250" swimtime="00:03:43.83" />
                    <SPLIT distance="300" swimtime="00:04:35.79" />
                    <SPLIT distance="350" swimtime="00:05:20.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="205" reactiontime="+94" swimtime="00:01:22.06" resultid="4810" heatid="9133" lane="0" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="474" reactiontime="+74" swimtime="00:01:45.93" resultid="4857" heatid="9111" lane="8" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                    <SPLIT distance="100" swimtime="00:00:55.50" />
                    <SPLIT distance="150" swimtime="00:01:21.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4805" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4826" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="4818" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="4834" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="3475" name="Steef Wrocław">
          <CONTACT city="Wrocław" email="ste1@wp.pl" name="Skrzypek Stefan" phone="500388374" street="Edyty Stein 6/1" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="3476">
              <RESULTS>
                <RESULT eventid="1113" points="164" reactiontime="+99" swimtime="00:03:20.18" resultid="3477" heatid="8924" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                    <SPLIT distance="100" swimtime="00:01:37.57" />
                    <SPLIT distance="150" swimtime="00:02:34.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="191" reactiontime="+103" swimtime="00:24:34.24" resultid="3478" heatid="8943" lane="9" entrytime="00:25:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                    <SPLIT distance="100" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:02:14.51" />
                    <SPLIT distance="200" swimtime="00:03:01.61" />
                    <SPLIT distance="250" swimtime="00:03:48.79" />
                    <SPLIT distance="300" swimtime="00:04:37.44" />
                    <SPLIT distance="350" swimtime="00:05:26.31" />
                    <SPLIT distance="400" swimtime="00:06:14.45" />
                    <SPLIT distance="450" swimtime="00:07:03.40" />
                    <SPLIT distance="500" swimtime="00:07:52.18" />
                    <SPLIT distance="550" swimtime="00:08:39.77" />
                    <SPLIT distance="600" swimtime="00:09:26.66" />
                    <SPLIT distance="650" swimtime="00:10:13.60" />
                    <SPLIT distance="700" swimtime="00:11:01.61" />
                    <SPLIT distance="750" swimtime="00:11:49.59" />
                    <SPLIT distance="800" swimtime="00:12:36.76" />
                    <SPLIT distance="850" swimtime="00:13:25.25" />
                    <SPLIT distance="900" swimtime="00:14:14.83" />
                    <SPLIT distance="950" swimtime="00:15:04.48" />
                    <SPLIT distance="1000" swimtime="00:15:54.36" />
                    <SPLIT distance="1050" swimtime="00:16:44.81" />
                    <SPLIT distance="1100" swimtime="00:17:38.08" />
                    <SPLIT distance="1150" swimtime="00:18:31.26" />
                    <SPLIT distance="1200" swimtime="00:19:24.69" />
                    <SPLIT distance="1250" swimtime="00:20:18.20" />
                    <SPLIT distance="1300" swimtime="00:21:12.66" />
                    <SPLIT distance="1350" swimtime="00:22:06.49" />
                    <SPLIT distance="1400" swimtime="00:22:56.81" />
                    <SPLIT distance="1450" swimtime="00:23:47.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="3479" heatid="9010" lane="5" entrytime="00:01:35.00" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="3480" heatid="9027" lane="6" entrytime="00:03:35.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="3481" heatid="9097" lane="9" entrytime="00:03:05.00" />
                <RESULT eventid="1578" points="176" reactiontime="+103" swimtime="00:07:00.12" resultid="3482" heatid="9118" lane="1" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                    <SPLIT distance="100" swimtime="00:01:38.97" />
                    <SPLIT distance="150" swimtime="00:02:35.79" />
                    <SPLIT distance="200" swimtime="00:03:32.04" />
                    <SPLIT distance="250" swimtime="00:04:31.50" />
                    <SPLIT distance="300" swimtime="00:05:27.06" />
                    <SPLIT distance="350" swimtime="00:06:15.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="163" reactiontime="+102" swimtime="00:01:28.66" resultid="3483" heatid="9131" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="215" reactiontime="+104" swimtime="00:05:54.16" resultid="3484" heatid="9185" lane="4" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:09.48" />
                    <SPLIT distance="200" swimtime="00:02:54.79" />
                    <SPLIT distance="250" swimtime="00:03:40.20" />
                    <SPLIT distance="300" swimtime="00:04:25.34" />
                    <SPLIT distance="350" swimtime="00:05:10.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WA" clubid="5894" name="SWIMMERS St. Pływackie">
          <CONTACT city="WARSZAWA" email="INFO@SWIMMERSTEAM.PL" name="GOŁĘBIOWSKI REMIGIUSZ" phone="601333782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1993-12-20" firstname="Arkadiusz" gender="M" lastname="Aptewicz" nation="POL" athleteid="5947">
              <RESULTS>
                <RESULT eventid="1239" points="616" reactiontime="+72" swimtime="00:02:21.55" resultid="5948" heatid="8978" lane="4" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="574" reactiontime="+73" swimtime="00:01:00.95" resultid="5949" heatid="9021" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="638" reactiontime="+70" swimtime="00:01:04.57" resultid="5950" heatid="9053" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="567" reactiontime="+68" swimtime="00:00:30.50" resultid="5951" heatid="9172" lane="3" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-03-03" firstname="Katarzyna" gender="F" lastname="Napora" nation="POL" athleteid="5903">
              <RESULTS>
                <RESULT eventid="1062" points="364" reactiontime="+82" swimtime="00:00:32.54" resultid="5904" heatid="8892" lane="9" entrytime="00:00:30.55" />
                <RESULT eventid="1256" points="326" reactiontime="+86" swimtime="00:01:14.09" resultid="5905" heatid="8983" lane="1" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="221" reactiontime="+82" swimtime="00:00:40.29" resultid="5906" heatid="9056" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1491" points="284" reactiontime="+89" swimtime="00:02:48.38" resultid="5907" heatid="9092" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.47" />
                    <SPLIT distance="150" swimtime="00:02:04.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brożyna" nation="POL" athleteid="5937">
              <RESULTS>
                <RESULT eventid="1205" points="269" reactiontime="+70" swimtime="00:00:34.41" resultid="5938" heatid="8961" lane="0" entrytime="00:00:33.40" />
                <RESULT eventid="1474" points="300" reactiontime="+71" swimtime="00:01:13.06" resultid="5939" heatid="9084" lane="3" entrytime="00:01:11.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="298" reactiontime="+80" swimtime="00:02:38.71" resultid="5940" heatid="9147" lane="5" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="100" swimtime="00:01:17.00" />
                    <SPLIT distance="150" swimtime="00:01:58.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-07-07" firstname="Remigiusz" gender="M" lastname="Gołębiowski" nation="POL" athleteid="5913">
              <RESULTS>
                <RESULT eventid="1079" points="451" reactiontime="+93" swimtime="00:00:26.40" resultid="5914" heatid="8912" lane="0" entrytime="00:00:26.50" />
                <RESULT eventid="1273" points="490" reactiontime="+87" swimtime="00:00:56.97" resultid="5915" heatid="8998" lane="3" entrytime="00:00:58.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="504" reactiontime="+85" swimtime="00:00:27.39" resultid="5916" heatid="9072" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1508" points="486" reactiontime="+83" swimtime="00:02:06.37" resultid="5917" heatid="9105" lane="3" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                    <SPLIT distance="100" swimtime="00:01:01.67" />
                    <SPLIT distance="150" swimtime="00:01:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="489" reactiontime="+84" swimtime="00:01:01.48" resultid="5918" heatid="9136" lane="3" entrytime="00:01:00.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-12-11" firstname="Mikołaj" gender="M" lastname="Tusiński" nation="POL" athleteid="5895">
              <RESULTS>
                <RESULT eventid="1079" points="437" reactiontime="+89" swimtime="00:00:26.68" resultid="5896" heatid="8911" lane="1" entrytime="00:00:26.70" />
                <RESULT eventid="1113" points="399" reactiontime="+86" swimtime="00:02:28.90" resultid="5897" heatid="8926" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="100" swimtime="00:01:10.89" />
                    <SPLIT distance="150" swimtime="00:01:54.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="463" reactiontime="+89" swimtime="00:00:58.06" resultid="5898" heatid="8999" lane="1" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="395" reactiontime="+89" swimtime="00:00:29.69" resultid="5899" heatid="9069" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1508" points="443" reactiontime="+84" swimtime="00:02:10.33" resultid="5900" heatid="9101" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:04.04" />
                    <SPLIT distance="150" swimtime="00:01:36.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="353" reactiontime="+86" swimtime="00:01:08.48" resultid="5901" heatid="9134" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="393" reactiontime="+88" swimtime="00:04:49.63" resultid="5902" heatid="9189" lane="0" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:47.08" />
                    <SPLIT distance="200" swimtime="00:02:24.69" />
                    <SPLIT distance="250" swimtime="00:03:01.24" />
                    <SPLIT distance="300" swimtime="00:03:37.01" />
                    <SPLIT distance="350" swimtime="00:04:13.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-12" firstname="Jan" gender="M" lastname="Rekowski" nation="POL" athleteid="5941">
              <RESULTS>
                <RESULT eventid="1079" points="480" reactiontime="+78" swimtime="00:00:25.87" resultid="5942" heatid="8914" lane="7" entrytime="00:00:25.80" />
                <RESULT eventid="1273" points="473" reactiontime="+75" swimtime="00:00:57.67" resultid="5943" heatid="8999" lane="9" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="357" reactiontime="+86" swimtime="00:01:11.38" resultid="5944" heatid="9019" lane="0" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="410" reactiontime="+78" swimtime="00:00:29.33" resultid="5945" heatid="9070" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1681" points="373" reactiontime="+76" swimtime="00:00:35.06" resultid="5946" heatid="9169" lane="5" entrytime="00:00:35.68" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-27" firstname="Remigiusz" gender="M" lastname="Miklewski" nation="POL" athleteid="5924">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="5925" heatid="8908" lane="9" entrytime="00:00:28.30" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="5926" heatid="8992" lane="5" entrytime="00:01:06.99" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="5927" heatid="9064" lane="9" entrytime="00:00:35.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-01" firstname="Katarzyna" gender="F" lastname="Koba" nation="POL" athleteid="5908">
              <RESULTS>
                <RESULT eventid="1062" points="433" reactiontime="+94" swimtime="00:00:30.71" resultid="5909" heatid="8892" lane="0" entrytime="00:00:30.40" />
                <RESULT eventid="1256" points="391" reactiontime="+91" swimtime="00:01:09.72" resultid="5910" heatid="8983" lane="2" entrytime="00:01:08.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="357" reactiontime="+90" swimtime="00:02:36.03" resultid="5911" heatid="9092" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:56.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="230" reactiontime="+96" swimtime="00:01:29.04" resultid="5912" heatid="9126" lane="2" entrytime="00:01:24.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-04" firstname="Norbert" gender="M" lastname="Tchorzewski" nation="POL" athleteid="5928">
              <RESULTS>
                <RESULT eventid="1113" points="218" reactiontime="+98" swimtime="00:03:02.00" resultid="5929" heatid="8925" lane="5" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                    <SPLIT distance="150" swimtime="00:02:18.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="236" reactiontime="+137" swimtime="00:22:54.35" resultid="5930" heatid="8943" lane="4" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="150" swimtime="00:02:08.26" />
                    <SPLIT distance="200" swimtime="00:02:54.32" />
                    <SPLIT distance="250" swimtime="00:03:39.90" />
                    <SPLIT distance="300" swimtime="00:04:26.17" />
                    <SPLIT distance="350" swimtime="00:05:11.22" />
                    <SPLIT distance="400" swimtime="00:05:56.92" />
                    <SPLIT distance="450" swimtime="00:06:42.38" />
                    <SPLIT distance="500" swimtime="00:07:27.80" />
                    <SPLIT distance="550" swimtime="00:08:13.46" />
                    <SPLIT distance="600" swimtime="00:08:59.58" />
                    <SPLIT distance="650" swimtime="00:09:45.44" />
                    <SPLIT distance="700" swimtime="00:10:31.41" />
                    <SPLIT distance="750" swimtime="00:11:16.60" />
                    <SPLIT distance="800" swimtime="00:12:03.81" />
                    <SPLIT distance="850" swimtime="00:12:49.44" />
                    <SPLIT distance="900" swimtime="00:13:35.25" />
                    <SPLIT distance="950" swimtime="00:14:21.98" />
                    <SPLIT distance="1000" swimtime="00:15:09.95" />
                    <SPLIT distance="1050" swimtime="00:15:55.71" />
                    <SPLIT distance="1100" swimtime="00:16:42.43" />
                    <SPLIT distance="1150" swimtime="00:17:30.05" />
                    <SPLIT distance="1200" swimtime="00:18:15.79" />
                    <SPLIT distance="1250" swimtime="00:19:01.65" />
                    <SPLIT distance="1300" swimtime="00:19:49.20" />
                    <SPLIT distance="1350" swimtime="00:20:35.92" />
                    <SPLIT distance="1400" swimtime="00:21:22.33" />
                    <SPLIT distance="1450" swimtime="00:22:09.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="277" reactiontime="+102" swimtime="00:01:08.92" resultid="5931" heatid="8993" lane="6" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="172" reactiontime="+114" swimtime="00:03:15.18" resultid="5932" heatid="9028" lane="2" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:28.47" />
                    <SPLIT distance="150" swimtime="00:02:19.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="271" reactiontime="+106" swimtime="00:02:33.50" resultid="5933" heatid="9099" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                    <SPLIT distance="150" swimtime="00:01:54.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="183" reactiontime="+113" swimtime="00:06:54.10" resultid="5934" heatid="9119" lane="0" entrytime="00:06:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:01:33.55" />
                    <SPLIT distance="150" swimtime="00:02:29.32" />
                    <SPLIT distance="200" swimtime="00:03:26.12" />
                    <SPLIT distance="250" swimtime="00:04:26.03" />
                    <SPLIT distance="300" swimtime="00:05:25.01" />
                    <SPLIT distance="350" swimtime="00:06:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="225" reactiontime="+107" swimtime="00:01:19.59" resultid="5935" heatid="9133" lane="9" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="250" reactiontime="+108" swimtime="00:05:36.88" resultid="5936" heatid="9187" lane="8" entrytime="00:05:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:17.11" />
                    <SPLIT distance="150" swimtime="00:02:00.09" />
                    <SPLIT distance="200" swimtime="00:02:44.30" />
                    <SPLIT distance="250" swimtime="00:03:27.66" />
                    <SPLIT distance="300" swimtime="00:04:12.90" />
                    <SPLIT distance="350" swimtime="00:04:58.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-03" firstname="Bolesław" gender="M" lastname="Porolniczak" nation="POL" athleteid="5919">
              <RESULTS>
                <RESULT eventid="1079" points="422" reactiontime="+84" swimtime="00:00:27.01" resultid="5920" heatid="8910" lane="5" entrytime="00:00:26.90" />
                <RESULT eventid="1273" points="400" reactiontime="+91" swimtime="00:01:00.95" resultid="5921" heatid="8997" lane="1" entrytime="00:01:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="362" reactiontime="+88" swimtime="00:01:11.07" resultid="5922" heatid="9017" lane="8" entrytime="00:01:11.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="365" reactiontime="+88" swimtime="00:00:30.48" resultid="5923" heatid="9069" lane="4" entrytime="00:00:29.70" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="404" reactiontime="+75" swimtime="00:02:02.40" resultid="5954" heatid="9035" lane="9" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:08.83" />
                    <SPLIT distance="150" swimtime="00:01:36.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5937" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="5941" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="5913" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="5895" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="499" reactiontime="+88" swimtime="00:01:44.07" resultid="5955" heatid="9111" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.00" />
                    <SPLIT distance="100" swimtime="00:00:53.31" />
                    <SPLIT distance="150" swimtime="00:01:18.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5919" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="5895" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="5913" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="5941" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="370" reactiontime="+85" swimtime="00:01:54.98" resultid="5952" heatid="8935" lane="1" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:00:58.34" />
                    <SPLIT distance="150" swimtime="00:01:28.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5903" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="5895" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="5908" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="5941" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="274" reactiontime="+80" swimtime="00:02:19.34" resultid="5953" heatid="9176" lane="9" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:01:13.06" />
                    <SPLIT distance="150" swimtime="00:01:46.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5903" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5941" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="5908" number="3" reactiontime="+85" />
                    <RELAYPOSITION athleteid="5928" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="U.B.O.T." nation="POL" region="OPO" clubid="2434" name="T.P &quot;U.B.O.T&quot; Masters Kędzierzyn-Koźle" shortname="T.P &quot;U.B.O.T&quot; Masters Kędzierz">
          <CONTACT city="Kędzierzyn-Koźle" email="marekkopij@wp.pl" name="Kopij Marek" phone="503-002-225" state="OPOLS" street="ul. Kościelna 17" zip="47-220" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-14" firstname="Sławomir" gender="M" lastname="Strzelczyk" nation="POL" athleteid="2459">
              <RESULTS>
                <RESULT eventid="1113" points="265" reactiontime="+94" swimtime="00:02:50.56" resultid="2460" heatid="8924" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:20.32" />
                    <SPLIT distance="150" swimtime="00:02:09.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="264" reactiontime="+87" swimtime="00:03:07.69" resultid="2461" heatid="8975" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                    <SPLIT distance="100" swimtime="00:01:30.67" />
                    <SPLIT distance="150" swimtime="00:02:19.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="286" reactiontime="+94" swimtime="00:01:16.85" resultid="2462" heatid="9012" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="220" reactiontime="+80" swimtime="00:02:55.60" resultid="2463" heatid="9146" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:26.48" />
                    <SPLIT distance="150" swimtime="00:02:12.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2464" heatid="9186" lane="1" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-05-14" firstname="Ewa" gender="F" lastname="Rojewska" nation="POL" athleteid="2442">
              <RESULTS>
                <RESULT eventid="1096" points="180" reactiontime="+74" swimtime="00:03:35.81" resultid="2443" heatid="8918" lane="9" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="100" swimtime="00:01:40.85" />
                    <SPLIT distance="150" swimtime="00:02:43.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="201" reactiontime="+94" swimtime="00:03:49.43" resultid="2444" heatid="8969" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.70" />
                    <SPLIT distance="100" swimtime="00:01:49.27" />
                    <SPLIT distance="150" swimtime="00:02:49.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="230" reactiontime="+77" swimtime="00:01:32.52" resultid="2445" heatid="9003" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="2446" heatid="9038" lane="3" entrytime="00:01:50.00" />
                <RESULT eventid="1423" points="218" reactiontime="+84" swimtime="00:00:40.45" resultid="2447" heatid="9056" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1595" points="144" reactiontime="+83" swimtime="00:01:44.17" resultid="2448" heatid="9125" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="218" reactiontime="+85" swimtime="00:00:47.79" resultid="2449" heatid="9153" lane="5" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-11" firstname="Aleksandra" gender="F" lastname="Dul" nation="POL" athleteid="2465">
              <RESULTS>
                <RESULT eventid="1187" points="410" reactiontime="+79" swimtime="00:00:34.54" resultid="2466" heatid="8951" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1290" points="358" reactiontime="+87" swimtime="00:01:19.79" resultid="2467" heatid="9004" lane="2" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="353" reactiontime="+90" swimtime="00:00:34.49" resultid="2468" heatid="9056" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1457" points="392" reactiontime="+83" swimtime="00:01:15.16" resultid="2469" heatid="9077" lane="8" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-08-18" firstname="Dorota" gender="F" lastname="Jaskulska" nation="POL" athleteid="2450">
              <RESULTS>
                <RESULT eventid="1062" points="251" reactiontime="+95" swimtime="00:00:36.82" resultid="2451" heatid="8889" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1096" points="188" reactiontime="+99" swimtime="00:03:32.54" resultid="2452" heatid="8917" lane="3" entrytime="00:03:35.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.56" />
                    <SPLIT distance="100" swimtime="00:01:41.67" />
                    <SPLIT distance="150" swimtime="00:02:45.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="230" reactiontime="+62" swimtime="00:00:41.86" resultid="2453" heatid="8950" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1290" points="217" reactiontime="+95" swimtime="00:01:34.33" resultid="2454" heatid="9003" lane="7" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="201" reactiontime="+62" swimtime="00:01:33.92" resultid="2455" heatid="9076" lane="9" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="215" reactiontime="+105" swimtime="00:03:04.73" resultid="2456" heatid="9090" lane="6" entrytime="00:03:12.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:27.01" />
                    <SPLIT distance="150" swimtime="00:02:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="197" reactiontime="+70" swimtime="00:03:24.79" resultid="2457" heatid="9139" lane="2" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                    <SPLIT distance="100" swimtime="00:01:39.82" />
                    <SPLIT distance="150" swimtime="00:02:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="221" reactiontime="+107" swimtime="00:06:27.73" resultid="2458" heatid="9179" lane="0" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                    <SPLIT distance="100" swimtime="00:01:26.12" />
                    <SPLIT distance="150" swimtime="00:02:14.71" />
                    <SPLIT distance="300" swimtime="00:04:45.59" />
                    <SPLIT distance="350" swimtime="00:05:37.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7089" name="T.P. Masters Opole">
          <CONTACT name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1967-01-01" firstname="Oskar" gender="M" lastname="Orski" nation="POL" athleteid="7116">
              <RESULTS>
                <RESULT eventid="1273" points="293" reactiontime="+103" swimtime="00:01:07.60" resultid="7117" heatid="8991" lane="6" entrytime="00:01:09.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Jerzy" gender="M" lastname="Minkiewicz" nation="POL" athleteid="7111">
              <RESULTS>
                <RESULT eventid="1079" points="257" reactiontime="+96" swimtime="00:00:31.83" resultid="7112" heatid="8903" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1273" points="253" reactiontime="+93" swimtime="00:01:10.98" resultid="7113" heatid="8991" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="201" reactiontime="+100" swimtime="00:01:26.37" resultid="7114" heatid="9012" lane="2" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="227" reactiontime="+98" swimtime="00:00:35.70" resultid="7115" heatid="9065" lane="0" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Grzegorz" gender="M" lastname="Radomski" nation="POL" athleteid="7090">
              <RESULTS>
                <RESULT eventid="1113" points="559" reactiontime="+76" swimtime="00:02:13.04" resultid="7091" heatid="8931" lane="8" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                    <SPLIT distance="100" swimtime="00:01:01.99" />
                    <SPLIT distance="150" swimtime="00:01:40.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="526" reactiontime="+74" swimtime="00:02:03.03" resultid="7092" heatid="9106" lane="9" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="100" swimtime="00:00:58.88" />
                    <SPLIT distance="150" swimtime="00:01:31.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="531" reactiontime="+75" swimtime="00:04:50.65" resultid="7093" heatid="9122" lane="5" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="150" swimtime="00:01:43.93" />
                    <SPLIT distance="200" swimtime="00:02:20.44" />
                    <SPLIT distance="250" swimtime="00:03:00.14" />
                    <SPLIT distance="300" swimtime="00:03:41.34" />
                    <SPLIT distance="350" swimtime="00:04:16.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="491" reactiontime="+64" swimtime="00:02:14.43" resultid="7094" heatid="9150" lane="7" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:05.17" />
                    <SPLIT distance="150" swimtime="00:01:39.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="532" reactiontime="+80" swimtime="00:04:21.94" resultid="7095" heatid="9192" lane="6" entrytime="00:04:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                    <SPLIT distance="100" swimtime="00:01:00.51" />
                    <SPLIT distance="150" swimtime="00:01:33.20" />
                    <SPLIT distance="200" swimtime="00:02:06.52" />
                    <SPLIT distance="250" swimtime="00:02:40.16" />
                    <SPLIT distance="300" swimtime="00:03:13.97" />
                    <SPLIT distance="350" swimtime="00:03:48.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="7104">
              <RESULTS>
                <RESULT eventid="1079" points="396" reactiontime="+87" swimtime="00:00:27.58" resultid="7105" heatid="8909" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1205" points="353" reactiontime="+67" swimtime="00:00:31.44" resultid="7106" heatid="8962" lane="2" entrytime="00:00:31.80" />
                <RESULT eventid="1273" points="393" reactiontime="+85" swimtime="00:01:01.32" resultid="7107" heatid="8996" lane="8" entrytime="00:01:01.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="390" reactiontime="+87" swimtime="00:00:29.82" resultid="7108" heatid="9061" lane="0" entrytime="00:00:47.50" />
                <RESULT eventid="1474" points="379" reactiontime="+65" swimtime="00:01:07.57" resultid="7109" heatid="9086" lane="9" entrytime="00:01:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="380" reactiontime="+67" swimtime="00:02:26.41" resultid="7110" heatid="9149" lane="2" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:11.49" />
                    <SPLIT distance="150" swimtime="00:01:49.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Witkowski" nation="POL" athleteid="7096">
              <RESULTS>
                <RESULT eventid="1079" points="142" reactiontime="+124" swimtime="00:00:38.77" resultid="7097" heatid="8898" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="7098" heatid="8921" lane="6" entrytime="00:04:55.00" />
                <RESULT eventid="1205" points="74" reactiontime="+98" swimtime="00:00:52.78" resultid="7099" heatid="8956" lane="1" entrytime="00:00:52.00" />
                <RESULT eventid="1273" points="99" reactiontime="+124" swimtime="00:01:37.08" resultid="7100" heatid="8987" lane="7" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="61" reactiontime="+95" swimtime="00:02:03.98" resultid="7101" heatid="9080" lane="7" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="7102" heatid="9144" lane="6" entrytime="00:04:25.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="7103" heatid="9161" lane="0" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Zbigniew" gender="M" lastname="Krasnodębski" nation="POL" athleteid="7118">
              <RESULTS>
                <RESULT eventid="1681" points="221" reactiontime="+85" swimtime="00:00:41.76" resultid="7119" heatid="9164" lane="8" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="242" reactiontime="+91" swimtime="00:02:12.40" resultid="7120" heatid="9110" lane="2" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="150" swimtime="00:01:42.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7104" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="7096" number="2" reactiontime="+92" />
                    <RELAYPOSITION athleteid="7111" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="7116" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3133" name="T.P. Skalar Słupsk">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-01" firstname="Beata" gender="F" lastname="Zubel" nation="POL" athleteid="3136">
              <RESULTS>
                <RESULT eventid="1147" points="342" reactiontime="+87" swimtime="00:11:24.97" resultid="3137" heatid="8939" lane="9" entrytime="00:11:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:19.04" />
                    <SPLIT distance="150" swimtime="00:02:00.98" />
                    <SPLIT distance="200" swimtime="00:02:43.58" />
                    <SPLIT distance="250" swimtime="00:03:26.71" />
                    <SPLIT distance="300" swimtime="00:04:10.18" />
                    <SPLIT distance="350" swimtime="00:04:53.47" />
                    <SPLIT distance="400" swimtime="00:05:36.67" />
                    <SPLIT distance="450" swimtime="00:06:20.20" />
                    <SPLIT distance="500" swimtime="00:07:03.80" />
                    <SPLIT distance="550" swimtime="00:07:48.08" />
                    <SPLIT distance="600" swimtime="00:08:32.38" />
                    <SPLIT distance="650" swimtime="00:09:17.16" />
                    <SPLIT distance="700" swimtime="00:10:01.22" />
                    <SPLIT distance="750" swimtime="00:10:44.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="335" reactiontime="+105" swimtime="00:02:39.35" resultid="3138" heatid="9092" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:01:57.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="352" reactiontime="+91" swimtime="00:05:31.99" resultid="3139" heatid="9180" lane="3" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:19.03" />
                    <SPLIT distance="150" swimtime="00:02:00.76" />
                    <SPLIT distance="200" swimtime="00:02:42.68" />
                    <SPLIT distance="250" swimtime="00:03:24.88" />
                    <SPLIT distance="300" swimtime="00:04:07.75" />
                    <SPLIT distance="350" swimtime="00:04:50.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5997" name="Tkkf Koszalin Masters">
          <CONTACT email="jakubkielar3@gmail.com" name="Jakub Kielar" />
          <ATHLETES>
            <ATHLETE birthdate="1960-01-01" firstname="Dorota" gender="F" lastname="Gudaniec" nation="POL" athleteid="6021">
              <RESULTS>
                <RESULT eventid="1147" points="232" reactiontime="+106" swimtime="00:12:59.19" resultid="6022" heatid="8938" lane="9" entrytime="00:13:15.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                    <SPLIT distance="150" swimtime="00:02:18.66" />
                    <SPLIT distance="200" swimtime="00:03:08.21" />
                    <SPLIT distance="250" swimtime="00:03:57.93" />
                    <SPLIT distance="300" swimtime="00:04:48.02" />
                    <SPLIT distance="350" swimtime="00:05:38.20" />
                    <SPLIT distance="400" swimtime="00:06:27.73" />
                    <SPLIT distance="450" swimtime="00:07:17.58" />
                    <SPLIT distance="500" swimtime="00:08:07.29" />
                    <SPLIT distance="550" swimtime="00:08:56.86" />
                    <SPLIT distance="600" swimtime="00:09:46.17" />
                    <SPLIT distance="650" swimtime="00:10:35.20" />
                    <SPLIT distance="700" swimtime="00:11:23.75" />
                    <SPLIT distance="750" swimtime="00:12:12.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="206" reactiontime="+110" swimtime="00:03:47.67" resultid="6023" heatid="8968" lane="5" entrytime="00:03:47.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.77" />
                    <SPLIT distance="100" swimtime="00:01:48.01" />
                    <SPLIT distance="150" swimtime="00:02:48.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="198" reactiontime="+95" swimtime="00:01:37.12" resultid="6024" heatid="9004" lane="9" entrytime="00:01:33.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="6025" heatid="9039" lane="2" entrytime="00:01:43.50" entrycourse="SCM" />
                <RESULT eventid="1555" points="207" reactiontime="+103" swimtime="00:07:19.28" resultid="6026" heatid="9114" lane="0" entrytime="00:07:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                    <SPLIT distance="100" swimtime="00:01:45.81" />
                    <SPLIT distance="150" swimtime="00:02:41.49" />
                    <SPLIT distance="200" swimtime="00:03:36.33" />
                    <SPLIT distance="250" swimtime="00:04:36.01" />
                    <SPLIT distance="300" swimtime="00:05:36.82" />
                    <SPLIT distance="350" swimtime="00:06:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="229" reactiontime="+103" swimtime="00:06:23.27" resultid="6027" heatid="9179" lane="8" entrytime="00:06:30.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                    <SPLIT distance="100" swimtime="00:01:29.53" />
                    <SPLIT distance="150" swimtime="00:02:17.80" />
                    <SPLIT distance="200" swimtime="00:03:07.39" />
                    <SPLIT distance="250" swimtime="00:03:57.00" />
                    <SPLIT distance="300" swimtime="00:04:46.69" />
                    <SPLIT distance="350" swimtime="00:05:35.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Aleksandra" gender="F" lastname="Kamińska" nation="POL" athleteid="6028">
              <RESULTS>
                <RESULT eventid="1062" points="117" reactiontime="+139" swimtime="00:00:47.50" resultid="6029" heatid="8887" lane="0" entrytime="00:00:43.00" entrycourse="SCM" />
                <RESULT eventid="1256" points="138" reactiontime="+112" swimtime="00:01:38.49" resultid="6030" heatid="8979" lane="5" entrytime="00:01:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="114" reactiontime="+125" swimtime="00:02:08.39" resultid="6031" heatid="9038" lane="8" entrytime="00:01:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="119" reactiontime="+132" swimtime="00:00:58.54" resultid="6032" heatid="9153" lane="0" entrytime="00:00:55.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Krzysztof" gender="M" lastname="Stefański" nation="POL" athleteid="5998">
              <RESULTS>
                <RESULT eventid="1079" points="368" reactiontime="+78" swimtime="00:00:28.25" resultid="5999" heatid="8907" lane="2" entrytime="00:00:28.90" entrycourse="SCM" />
                <RESULT eventid="1273" points="350" reactiontime="+72" swimtime="00:01:03.74" resultid="6000" heatid="8993" lane="3" entrytime="00:01:05.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="260" reactiontime="+83" swimtime="00:02:35.62" resultid="6001" heatid="9098" lane="2" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K15 - Brak dotknięcia ściany obydwoma rozłączonymi dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 20:40)" eventid="1578" reactiontime="+84" status="DSQ" swimtime="00:07:00.32" resultid="6002" heatid="9118" lane="4" entrytime="00:06:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:33.12" />
                    <SPLIT distance="150" swimtime="00:02:27.25" />
                    <SPLIT distance="200" swimtime="00:03:22.18" />
                    <SPLIT distance="250" swimtime="00:04:27.81" />
                    <SPLIT distance="300" swimtime="00:05:31.18" />
                    <SPLIT distance="350" swimtime="00:06:18.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="6003" heatid="9164" lane="1" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Jarosław" gender="M" lastname="Winiarczyk" nation="POL" athleteid="6004">
              <RESULTS>
                <RESULT eventid="1165" points="292" reactiontime="+89" swimtime="00:21:20.08" resultid="6005" heatid="8945" lane="8" entrytime="00:21:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:12.87" />
                    <SPLIT distance="150" swimtime="00:01:52.42" />
                    <SPLIT distance="200" swimtime="00:02:33.15" />
                    <SPLIT distance="250" swimtime="00:03:14.55" />
                    <SPLIT distance="300" swimtime="00:03:56.72" />
                    <SPLIT distance="350" swimtime="00:04:39.23" />
                    <SPLIT distance="400" swimtime="00:05:22.60" />
                    <SPLIT distance="450" swimtime="00:06:06.12" />
                    <SPLIT distance="500" swimtime="00:06:50.10" />
                    <SPLIT distance="550" swimtime="00:07:33.96" />
                    <SPLIT distance="600" swimtime="00:08:18.06" />
                    <SPLIT distance="650" swimtime="00:09:01.48" />
                    <SPLIT distance="700" swimtime="00:09:45.25" />
                    <SPLIT distance="750" swimtime="00:10:29.11" />
                    <SPLIT distance="800" swimtime="00:11:13.18" />
                    <SPLIT distance="850" swimtime="00:11:57.57" />
                    <SPLIT distance="900" swimtime="00:12:41.79" />
                    <SPLIT distance="950" swimtime="00:13:25.57" />
                    <SPLIT distance="1000" swimtime="00:14:09.83" />
                    <SPLIT distance="1050" swimtime="00:14:54.63" />
                    <SPLIT distance="1100" swimtime="00:15:39.03" />
                    <SPLIT distance="1150" swimtime="00:16:23.00" />
                    <SPLIT distance="1200" swimtime="00:17:06.21" />
                    <SPLIT distance="1250" swimtime="00:17:49.63" />
                    <SPLIT distance="1300" swimtime="00:18:32.92" />
                    <SPLIT distance="1350" swimtime="00:19:14.92" />
                    <SPLIT distance="1400" swimtime="00:19:57.72" />
                    <SPLIT distance="1450" swimtime="00:20:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="351" reactiontime="+83" swimtime="00:01:03.65" resultid="6006" heatid="8994" lane="6" entrytime="00:01:03.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="316" reactiontime="+69" swimtime="00:02:25.83" resultid="6007" heatid="9103" lane="9" entrytime="00:02:17.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                    <SPLIT distance="100" swimtime="00:01:08.54" />
                    <SPLIT distance="150" swimtime="00:01:48.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="314" reactiontime="+84" swimtime="00:05:11.98" resultid="6008" heatid="9188" lane="3" entrytime="00:05:13.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="150" swimtime="00:01:49.63" />
                    <SPLIT distance="200" swimtime="00:02:30.06" />
                    <SPLIT distance="250" swimtime="00:03:11.28" />
                    <SPLIT distance="300" swimtime="00:03:52.96" />
                    <SPLIT distance="350" swimtime="00:04:34.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Stankiewicz - Majkowska" gender="F" lastname="Joanna" nation="POL" athleteid="6009">
              <RESULTS>
                <RESULT eventid="1096" points="182" reactiontime="+91" swimtime="00:03:34.97" resultid="6010" heatid="8917" lane="4" entrytime="00:03:33.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                    <SPLIT distance="100" swimtime="00:01:41.50" />
                    <SPLIT distance="150" swimtime="00:02:41.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="6011" heatid="8949" lane="4" entrytime="00:00:46.91" entrycourse="SCM" />
                <RESULT eventid="1290" points="198" reactiontime="+83" swimtime="00:01:37.12" resultid="6012" heatid="9003" lane="4" entrytime="00:01:34.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="6013" heatid="9039" lane="1" entrytime="00:01:46.72" entrycourse="SCM" />
                <RESULT eventid="1555" points="193" reactiontime="+81" swimtime="00:07:29.07" resultid="6014" heatid="9114" lane="9" entrytime="00:07:51.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                    <SPLIT distance="100" swimtime="00:01:47.16" />
                    <SPLIT distance="150" swimtime="00:02:45.89" />
                    <SPLIT distance="200" swimtime="00:03:44.04" />
                    <SPLIT distance="250" swimtime="00:04:43.65" />
                    <SPLIT distance="300" swimtime="00:05:43.96" />
                    <SPLIT distance="350" swimtime="00:06:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="218" reactiontime="+84" swimtime="00:00:47.79" resultid="6015" heatid="9154" lane="3" entrytime="00:00:47.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Joanna" gender="F" lastname="Wojciechowska" nation="POL" athleteid="6016">
              <RESULTS>
                <RESULT eventid="1062" points="243" reactiontime="+81" swimtime="00:00:37.22" resultid="6017" heatid="8889" lane="9" entrytime="00:00:37.05" entrycourse="SCM" />
                <RESULT eventid="1187" points="163" reactiontime="+77" swimtime="00:00:46.95" resultid="6018" heatid="8950" lane="9" entrytime="00:00:46.70" entrycourse="SCM" />
                <RESULT eventid="1256" points="207" reactiontime="+88" swimtime="00:01:26.23" resultid="6019" heatid="8980" lane="5" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="194" reactiontime="+87" swimtime="00:00:49.67" resultid="6020" heatid="9154" lane="7" entrytime="00:00:48.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="6035" heatid="9108" lane="0" entrytime="00:03:25.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6021" number="1" />
                    <RELAYPOSITION athleteid="6028" number="2" />
                    <RELAYPOSITION athleteid="6009" number="3" />
                    <RELAYPOSITION athleteid="6016" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="247" reactiontime="+73" swimtime="00:02:11.50" resultid="6033" heatid="8933" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="100" swimtime="00:01:07.58" />
                    <SPLIT distance="150" swimtime="00:01:43.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6009" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="6016" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="6004" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="5998" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="206" reactiontime="+77" swimtime="00:02:33.21" resultid="6034" heatid="9174" lane="2" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.34" />
                    <SPLIT distance="100" swimtime="00:01:32.73" />
                    <SPLIT distance="150" swimtime="00:02:05.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6009" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="6021" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="5998" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="6004" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02602" nation="POL" region="KUJ" clubid="2476" name="Toruń Multisport Team">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1978-01-23" firstname="Marcin" gender="M" lastname="Mykowski" nation="POL" athleteid="2501">
              <RESULTS>
                <RESULT eventid="1273" points="486" reactiontime="+77" swimtime="00:00:57.13" resultid="2502" heatid="8997" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="422" reactiontime="+66" swimtime="00:01:05.23" resultid="2503" heatid="9085" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="369" reactiontime="+93" swimtime="00:02:18.53" resultid="2504" heatid="9103" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="150" swimtime="00:01:45.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="379" reactiontime="+70" swimtime="00:02:26.60" resultid="2505" heatid="9149" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                    <SPLIT distance="150" swimtime="00:01:49.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="2506">
              <RESULTS>
                <RESULT eventid="1096" points="308" reactiontime="+80" swimtime="00:03:00.42" resultid="2507" heatid="8918" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:24.48" />
                    <SPLIT distance="150" swimtime="00:02:17.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="276" reactiontime="+80" swimtime="00:12:16.19" resultid="2508" heatid="8938" lane="7" entrytime="00:12:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:08.40" />
                    <SPLIT distance="200" swimtime="00:02:54.54" />
                    <SPLIT distance="250" swimtime="00:03:40.85" />
                    <SPLIT distance="300" swimtime="00:04:27.06" />
                    <SPLIT distance="350" swimtime="00:05:13.20" />
                    <SPLIT distance="400" swimtime="00:06:00.46" />
                    <SPLIT distance="450" swimtime="00:06:46.87" />
                    <SPLIT distance="500" swimtime="00:07:33.15" />
                    <SPLIT distance="550" swimtime="00:08:20.10" />
                    <SPLIT distance="600" swimtime="00:09:07.07" />
                    <SPLIT distance="650" swimtime="00:09:54.53" />
                    <SPLIT distance="700" swimtime="00:10:42.62" />
                    <SPLIT distance="750" swimtime="00:11:30.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="288" reactiontime="+80" swimtime="00:03:23.70" resultid="2509" heatid="8969" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                    <SPLIT distance="100" swimtime="00:01:34.68" />
                    <SPLIT distance="150" swimtime="00:02:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="2510" heatid="9023" lane="3" entrytime="00:03:50.00" />
                <RESULT eventid="1388" points="288" reactiontime="+75" swimtime="00:01:34.42" resultid="2511" heatid="9040" lane="8" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="296" reactiontime="+84" swimtime="00:06:29.52" resultid="2512" heatid="9114" lane="1" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:31.89" />
                    <SPLIT distance="150" swimtime="00:02:19.95" />
                    <SPLIT distance="200" swimtime="00:03:06.27" />
                    <SPLIT distance="250" swimtime="00:03:59.96" />
                    <SPLIT distance="300" swimtime="00:04:55.65" />
                    <SPLIT distance="350" swimtime="00:05:43.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="219" reactiontime="+82" swimtime="00:01:30.58" resultid="2513" heatid="9124" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="289" reactiontime="+78" swimtime="00:05:54.52" resultid="2514" heatid="9180" lane="9" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:22.57" />
                    <SPLIT distance="150" swimtime="00:02:06.97" />
                    <SPLIT distance="200" swimtime="00:02:51.77" />
                    <SPLIT distance="250" swimtime="00:03:37.33" />
                    <SPLIT distance="300" swimtime="00:04:23.39" />
                    <SPLIT distance="350" swimtime="00:05:09.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="2477">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="2478" heatid="8896" lane="3" entrytime="00:00:42.45" />
                <RESULT eventid="1205" points="71" reactiontime="+80" swimtime="00:00:53.58" resultid="2479" heatid="8956" lane="8" entrytime="00:00:53.10" />
                <RESULT eventid="1239" points="86" reactiontime="+104" swimtime="00:04:32.42" resultid="2480" heatid="8972" lane="8" entrytime="00:04:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.68" />
                    <SPLIT distance="100" swimtime="00:02:05.08" />
                    <SPLIT distance="150" swimtime="00:03:19.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="102" reactiontime="+108" swimtime="00:01:58.80" resultid="2481" heatid="9044" lane="6" entrytime="00:01:59.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="2482" heatid="9079" lane="4" entrytime="00:02:11.24" />
                <RESULT eventid="1681" points="116" reactiontime="+97" swimtime="00:00:51.75" resultid="2483" heatid="9161" lane="2" entrytime="00:00:49.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="2493">
              <RESULTS>
                <RESULT eventid="1079" points="110" reactiontime="+101" swimtime="00:00:42.24" resultid="2494" heatid="8896" lane="5" entrytime="00:00:41.25" />
                <RESULT eventid="1205" points="45" reactiontime="+95" swimtime="00:01:02.41" resultid="2495" heatid="8955" lane="2" entrytime="00:00:59.24" />
                <RESULT eventid="1273" points="81" reactiontime="+102" swimtime="00:01:43.67" resultid="2496" heatid="8987" lane="9" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="39" reactiontime="+102" swimtime="00:05:12.03" resultid="2497" heatid="9143" lane="5" entrytime="00:05:18.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.35" />
                    <SPLIT distance="100" swimtime="00:02:30.85" />
                    <SPLIT distance="150" swimtime="00:03:53.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="43" reactiontime="+69" swimtime="00:02:19.03" resultid="3041" heatid="9079" lane="5" entrytime="00:02:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="Szufarski" nation="POL" athleteid="2523">
              <RESULTS>
                <RESULT eventid="1113" reactiontime="+103" status="DNF" swimtime="00:00:00.00" resultid="2524" heatid="8923" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="134" reactiontime="+102" swimtime="00:01:38.76" resultid="2525" heatid="9010" lane="2" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="125" reactiontime="+102" swimtime="00:00:43.55" resultid="2526" heatid="9061" lane="5" entrytime="00:00:42.50" />
                <RESULT eventid="1578" points="94" reactiontime="+112" swimtime="00:08:37.16" resultid="2527" heatid="9117" lane="2" entrytime="00:08:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.03" />
                    <SPLIT distance="100" swimtime="00:03:00.93" />
                    <SPLIT distance="150" swimtime="00:04:04.55" />
                    <SPLIT distance="200" swimtime="00:05:10.33" />
                    <SPLIT distance="250" swimtime="00:06:18.55" />
                    <SPLIT distance="300" swimtime="00:07:18.11" />
                    <SPLIT distance="350" swimtime="00:08:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="87" reactiontime="+113" swimtime="00:01:48.92" resultid="2528" heatid="9130" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="139" reactiontime="+103" swimtime="00:00:48.73" resultid="2529" heatid="9162" lane="9" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-14" firstname="Marta" gender="F" lastname="Lord" nation="POL" athleteid="2530">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1062" points="569" reactiontime="+76" swimtime="00:00:28.03" resultid="2531" heatid="8892" lane="4" entrytime="00:00:29.50" />
                <RESULT comment="Rekord Polski" eventid="1187" points="445" reactiontime="+77" swimtime="00:00:33.61" resultid="2532" heatid="8953" lane="9" entrytime="00:00:33.90" />
                <RESULT comment="Rekord Polski" eventid="1290" points="480" reactiontime="+76" swimtime="00:01:12.39" resultid="2533" heatid="9007" lane="8" entrytime="00:01:13.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="448" reactiontime="+81" swimtime="00:01:21.45" resultid="2534" heatid="9042" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1457" points="450" reactiontime="+81" swimtime="00:01:11.81" resultid="2535" heatid="9078" lane="8" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1630" points="447" reactiontime="+88" swimtime="00:02:35.85" resultid="2536" heatid="9141" lane="6" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:01:56.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="443" reactiontime="+82" swimtime="00:00:37.77" resultid="2537" heatid="9158" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="Osóbka" nation="POL" athleteid="2498">
              <RESULTS>
                <RESULT eventid="1079" points="34" reactiontime="+122" swimtime="00:01:02.27" resultid="2499" heatid="8895" lane="3" entrytime="00:00:59.58" />
                <RESULT eventid="1681" points="27" reactiontime="+126" swimtime="00:01:23.26" resultid="2500" heatid="9160" lane="0" entrytime="00:01:19.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="2538">
              <RESULTS>
                <RESULT eventid="1079" points="312" reactiontime="+82" swimtime="00:00:29.85" resultid="2539" heatid="8898" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1113" points="240" reactiontime="+94" swimtime="00:02:56.21" resultid="2540" heatid="8925" lane="0" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:01:24.04" />
                    <SPLIT distance="150" swimtime="00:02:16.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="303" reactiontime="+85" swimtime="00:01:06.84" resultid="2541" heatid="8991" lane="9" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="218" reactiontime="+99" swimtime="00:03:00.36" resultid="2542" heatid="9028" lane="8" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="150" swimtime="00:02:11.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="275" reactiontime="+87" swimtime="00:02:32.79" resultid="2543" heatid="9097" lane="4" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                    <SPLIT distance="150" swimtime="00:01:53.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="233" reactiontime="+106" swimtime="00:06:22.46" resultid="2544" heatid="9119" lane="2" entrytime="00:06:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:21.86" />
                    <SPLIT distance="150" swimtime="00:02:16.48" />
                    <SPLIT distance="200" swimtime="00:03:09.07" />
                    <SPLIT distance="250" swimtime="00:04:01.96" />
                    <SPLIT distance="300" swimtime="00:04:56.65" />
                    <SPLIT distance="350" swimtime="00:05:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="274" reactiontime="+92" swimtime="00:01:14.51" resultid="2545" heatid="9132" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2546" heatid="9186" lane="3" entrytime="00:05:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="2515">
              <RESULTS>
                <RESULT eventid="1096" points="430" reactiontime="+84" swimtime="00:02:41.40" resultid="2516" heatid="8920" lane="6" entrytime="00:02:44.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:15.62" />
                    <SPLIT distance="150" swimtime="00:02:01.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="425" reactiontime="+81" swimtime="00:02:58.97" resultid="2517" heatid="8970" lane="5" entrytime="00:03:05.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:25.87" />
                    <SPLIT distance="150" swimtime="00:02:12.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="443" reactiontime="+79" swimtime="00:01:14.33" resultid="2518" heatid="9007" lane="9" entrytime="00:01:14.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="411" reactiontime="+87" swimtime="00:01:23.87" resultid="2519" heatid="9042" lane="2" entrytime="00:01:24.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1555" points="394" reactiontime="+92" swimtime="00:05:54.44" resultid="2520" heatid="9115" lane="2" entrytime="00:06:01.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:23.10" />
                    <SPLIT distance="150" swimtime="00:02:08.45" />
                    <SPLIT distance="200" swimtime="00:02:53.64" />
                    <SPLIT distance="250" swimtime="00:03:41.92" />
                    <SPLIT distance="300" swimtime="00:04:30.62" />
                    <SPLIT distance="350" swimtime="00:05:13.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="381" reactiontime="+86" swimtime="00:01:15.31" resultid="2521" heatid="9127" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="416" reactiontime="+80" swimtime="00:00:38.57" resultid="2522" heatid="9157" lane="5" entrytime="00:00:39.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-01" firstname="Adrian" gender="M" lastname="Bilski" nation="POL" athleteid="2547">
              <RESULTS>
                <RESULT eventid="1079" points="187" reactiontime="+130" swimtime="00:00:35.40" resultid="2548" heatid="8898" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1273" points="182" reactiontime="+122" swimtime="00:01:19.23" resultid="2549" heatid="8988" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="155" reactiontime="+110" swimtime="00:03:04.95" resultid="2550" heatid="9094" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                    <SPLIT distance="100" swimtime="00:01:29.78" />
                    <SPLIT distance="150" swimtime="00:02:17.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="142" reactiontime="+112" swimtime="00:06:46.51" resultid="2551" heatid="9183" lane="8" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="2484">
              <RESULTS>
                <RESULT eventid="1113" points="53" reactiontime="+124" swimtime="00:04:51.42" resultid="2485" heatid="8921" lane="3" entrytime="00:04:31.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.73" />
                    <SPLIT distance="100" swimtime="00:02:31.86" />
                    <SPLIT distance="150" swimtime="00:03:56.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2486" heatid="8940" lane="4" entrytime="00:38:24.14" />
                <RESULT eventid="1273" points="63" reactiontime="+125" swimtime="00:01:52.50" resultid="2487" heatid="8987" lane="8" entrytime="00:01:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="2488" heatid="9025" lane="6" entrytime="00:05:10.00" />
                <RESULT eventid="1508" points="60" reactiontime="+134" swimtime="00:04:13.37" resultid="2489" heatid="9095" lane="6" entrytime="00:03:42.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.91" />
                    <SPLIT distance="100" swimtime="00:02:04.77" />
                    <SPLIT distance="150" swimtime="00:03:12.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="2490" heatid="9116" lane="5" entrytime="00:09:48.45" />
                <RESULT eventid="1613" points="34" reactiontime="+124" swimtime="00:02:28.34" resultid="2491" heatid="9129" lane="8" entrytime="00:02:14.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="31" reactiontime="+88" swimtime="00:05:37.72" resultid="2492" heatid="9143" lane="4" entrytime="00:05:15.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.63" />
                    <SPLIT distance="100" swimtime="00:02:46.26" />
                    <SPLIT distance="150" swimtime="00:04:13.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="56" reactiontime="+80" swimtime="00:03:56.11" resultid="2552" heatid="9032" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.72" />
                    <SPLIT distance="100" swimtime="00:02:14.65" />
                    <SPLIT distance="150" swimtime="00:03:16.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2477" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2498" number="2" reactiontime="+84" />
                    <RELAYPOSITION athleteid="2484" number="3" reactiontime="+104" />
                    <RELAYPOSITION athleteid="2493" number="4" reactiontime="+91" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="76" reactiontime="+103" swimtime="00:03:14.59" resultid="2553" heatid="9109" lane="7" entrytime="00:03:21.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="100" swimtime="00:01:44.36" />
                    <SPLIT distance="150" swimtime="00:02:31.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2477" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="2498" number="2" reactiontime="+91" />
                    <RELAYPOSITION athleteid="2484" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2493" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="381" reactiontime="+81" swimtime="00:01:53.85" resultid="2554" heatid="8935" lane="8" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:00:59.38" />
                    <SPLIT distance="150" swimtime="00:01:27.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2538" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2515" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2530" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="2501" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="331" reactiontime="+77" swimtime="00:02:10.82" resultid="2555" heatid="9176" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="150" swimtime="00:01:44.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2530" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2515" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2538" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2501" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="4628" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="4643">
              <RESULTS>
                <RESULT eventid="1079" points="145" reactiontime="+105" swimtime="00:00:38.53" resultid="4644" heatid="8898" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1113" points="117" reactiontime="+106" swimtime="00:03:43.55" resultid="4645" heatid="8923" lane="9" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.88" />
                    <SPLIT distance="100" swimtime="00:01:50.10" />
                    <SPLIT distance="150" swimtime="00:02:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="117" reactiontime="+80" swimtime="00:00:45.32" resultid="4646" heatid="8957" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="1307" points="119" reactiontime="+96" swimtime="00:01:42.79" resultid="4647" heatid="9010" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="106" reactiontime="+97" swimtime="00:01:43.36" resultid="4648" heatid="9081" lane="0" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="104" reactiontime="+85" swimtime="00:03:44.96" resultid="4649" heatid="9145" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.96" />
                    <SPLIT distance="100" swimtime="00:01:48.94" />
                    <SPLIT distance="150" swimtime="00:02:47.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="137" reactiontime="+103" swimtime="00:00:48.93" resultid="4650" heatid="9161" lane="6" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="4671" />
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="4651">
              <RESULTS>
                <RESULT eventid="1079" points="157" reactiontime="+84" swimtime="00:00:37.49" resultid="4652" heatid="8898" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1205" points="145" reactiontime="+86" swimtime="00:00:42.21" resultid="4653" heatid="8957" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1474" points="136" reactiontime="+80" swimtime="00:01:34.95" resultid="4654" heatid="9081" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="106" reactiontime="+92" swimtime="00:03:43.97" resultid="4655" heatid="9145" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.64" />
                    <SPLIT distance="100" swimtime="00:01:51.09" />
                    <SPLIT distance="150" swimtime="00:02:49.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="4656" heatid="9184" lane="0" entrytime="00:07:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" athleteid="4665">
              <RESULTS>
                <RESULT eventid="1113" points="190" reactiontime="+95" swimtime="00:03:10.44" resultid="4666" heatid="8924" lane="3" entrytime="00:03:15.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:30.23" />
                    <SPLIT distance="150" swimtime="00:02:23.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="215" reactiontime="+100" swimtime="00:03:20.93" resultid="4667" heatid="8973" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                    <SPLIT distance="100" swimtime="00:01:34.93" />
                    <SPLIT distance="150" swimtime="00:02:26.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="214" reactiontime="+89" swimtime="00:01:32.87" resultid="4668" heatid="9047" lane="7" entrytime="00:01:30.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="162" reactiontime="+103" swimtime="00:07:11.21" resultid="4669" heatid="9118" lane="7" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                    <SPLIT distance="100" swimtime="00:01:43.72" />
                    <SPLIT distance="150" swimtime="00:02:40.76" />
                    <SPLIT distance="200" swimtime="00:03:37.33" />
                    <SPLIT distance="250" swimtime="00:04:36.00" />
                    <SPLIT distance="300" swimtime="00:05:33.74" />
                    <SPLIT distance="350" swimtime="00:06:23.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="136" reactiontime="+91" swimtime="00:03:25.85" resultid="4670" heatid="9145" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.13" />
                    <SPLIT distance="100" swimtime="00:01:38.76" />
                    <SPLIT distance="150" swimtime="00:02:31.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="4629">
              <RESULTS>
                <RESULT eventid="1062" points="209" reactiontime="+91" swimtime="00:00:39.15" resultid="4630" heatid="8888" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="1187" points="139" reactiontime="+80" swimtime="00:00:49.53" resultid="4631" heatid="8949" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1290" points="149" reactiontime="+97" swimtime="00:01:46.79" resultid="4632" heatid="9002" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="118" reactiontime="+96" swimtime="00:00:49.59" resultid="4633" heatid="9054" lane="5" entrytime="00:00:53.00" />
                <RESULT eventid="1457" points="119" reactiontime="+86" swimtime="00:01:51.82" resultid="4634" heatid="9075" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="153" reactiontime="+97" swimtime="00:00:53.76" resultid="4635" heatid="9153" lane="7" entrytime="00:00:53.00" />
                <RESULT eventid="1721" points="160" reactiontime="+103" swimtime="00:07:11.88" resultid="4636" heatid="9178" lane="7" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                    <SPLIT distance="100" swimtime="00:01:40.98" />
                    <SPLIT distance="150" swimtime="00:02:39.72" />
                    <SPLIT distance="200" swimtime="00:03:34.80" />
                    <SPLIT distance="250" swimtime="00:04:29.96" />
                    <SPLIT distance="300" swimtime="00:05:27.16" />
                    <SPLIT distance="350" swimtime="00:06:20.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Anna" gender="F" lastname="Gano-Kosturkiewicz" nation="POL" athleteid="4637">
              <RESULTS>
                <RESULT eventid="1062" points="157" reactiontime="+111" swimtime="00:00:43.06" resultid="4638" heatid="8887" lane="8" entrytime="00:00:43.00" />
                <RESULT eventid="1187" points="104" reactiontime="+93" swimtime="00:00:54.55" resultid="4639" heatid="8949" lane="1" entrytime="00:00:54.00" />
                <RESULT eventid="1423" points="122" reactiontime="+113" swimtime="00:00:49.04" resultid="4640" heatid="9055" lane="6" entrytime="00:00:47.00" />
                <RESULT eventid="1457" points="88" reactiontime="+82" swimtime="00:02:03.40" resultid="4641" heatid="9075" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="88" reactiontime="+125" swimtime="00:02:02.46" resultid="4642" heatid="9124" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="4657">
              <RESULTS>
                <RESULT eventid="1113" points="202" reactiontime="+99" swimtime="00:03:06.54" resultid="4658" heatid="8925" lane="1" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                    <SPLIT distance="100" swimtime="00:01:31.02" />
                    <SPLIT distance="150" swimtime="00:02:23.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="163" reactiontime="+73" swimtime="00:00:40.66" resultid="4659" heatid="8958" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1307" points="210" reactiontime="+93" swimtime="00:01:25.10" resultid="4660" heatid="9012" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="181" reactiontime="+75" swimtime="00:01:26.46" resultid="4661" heatid="9082" lane="7" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="193" reactiontime="+96" swimtime="00:06:47.21" resultid="4662" heatid="9119" lane="6" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                    <SPLIT distance="100" swimtime="00:01:42.60" />
                    <SPLIT distance="150" swimtime="00:02:32.58" />
                    <SPLIT distance="200" swimtime="00:03:22.13" />
                    <SPLIT distance="250" swimtime="00:04:17.82" />
                    <SPLIT distance="300" swimtime="00:05:13.87" />
                    <SPLIT distance="350" swimtime="00:06:01.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="174" reactiontime="+80" swimtime="00:03:10.01" resultid="4663" heatid="9147" lane="9" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                    <SPLIT distance="100" swimtime="00:01:33.24" />
                    <SPLIT distance="150" swimtime="00:02:22.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="226" reactiontime="+98" swimtime="00:00:41.44" resultid="4664" heatid="9165" lane="0" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="184" reactiontime="+89" swimtime="00:02:39.10" resultid="4677" heatid="9032" lane="4" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:01:23.55" />
                    <SPLIT distance="150" swimtime="00:02:00.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4651" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="4657" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="4665" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="4643" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WIE" clubid="2089" name="UKS CITYZEN Poznań">
          <CONTACT name="roszak" />
          <ATHLETES>
            <ATHLETE birthdate="1977-09-24" firstname="Adam" gender="M" lastname="Kijowski" nation="POL" athleteid="2099">
              <RESULTS>
                <RESULT eventid="1079" points="234" reactiontime="+80" swimtime="00:00:32.86" resultid="2100" heatid="8894" lane="7" />
                <RESULT eventid="1239" points="213" reactiontime="+83" swimtime="00:03:21.47" resultid="2101" heatid="8977" lane="1" entrytime="00:02:50.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:01:28.71" />
                    <SPLIT distance="150" swimtime="00:02:23.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="194" reactiontime="+80" swimtime="00:01:27.41" resultid="2102" heatid="9011" lane="5" entrytime="00:01:27.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="251" reactiontime="+82" swimtime="00:01:28.10" resultid="2103" heatid="9050" lane="6" entrytime="00:01:22.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="230" reactiontime="+81" swimtime="00:00:41.16" resultid="2104" heatid="9166" lane="5" entrytime="00:00:38.48" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-10" firstname="Krzysztof" gender="M" lastname="Grzegorzewicz" nation="POL" athleteid="2152">
              <RESULTS>
                <RESULT eventid="1113" points="345" reactiontime="+80" swimtime="00:02:36.20" resultid="2153" heatid="8930" lane="3" entrytime="00:02:20.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:11.24" />
                    <SPLIT distance="150" swimtime="00:01:58.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="380" reactiontime="+83" swimtime="00:01:09.92" resultid="2154" heatid="9019" lane="3" entrytime="00:01:06.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="399" reactiontime="+88" swimtime="00:00:29.60" resultid="2155" heatid="9071" lane="4" entrytime="00:00:27.63" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="2156" heatid="9136" lane="6" entrytime="00:01:01.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-05" firstname="Kinga" gender="F" lastname="Jaruga" nation="POL" athleteid="2147">
              <RESULTS>
                <RESULT eventid="1147" points="262" reactiontime="+84" swimtime="00:12:28.26" resultid="2148" heatid="8937" lane="5" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:23.03" />
                    <SPLIT distance="150" swimtime="00:02:10.16" />
                    <SPLIT distance="200" swimtime="00:02:57.44" />
                    <SPLIT distance="250" swimtime="00:03:45.12" />
                    <SPLIT distance="300" swimtime="00:04:32.88" />
                    <SPLIT distance="350" swimtime="00:05:20.54" />
                    <SPLIT distance="400" swimtime="00:06:08.60" />
                    <SPLIT distance="450" swimtime="00:06:56.53" />
                    <SPLIT distance="500" swimtime="00:07:44.59" />
                    <SPLIT distance="550" swimtime="00:08:32.41" />
                    <SPLIT distance="600" swimtime="00:09:20.68" />
                    <SPLIT distance="650" swimtime="00:10:08.54" />
                    <SPLIT distance="700" swimtime="00:10:56.73" />
                    <SPLIT distance="750" swimtime="00:11:44.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="264" reactiontime="+81" swimtime="00:01:19.50" resultid="2149" heatid="8981" lane="2" entrytime="00:01:18.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="259" reactiontime="+81" swimtime="00:02:53.67" resultid="2150" heatid="9092" lane="9" entrytime="00:02:41.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                    <SPLIT distance="100" swimtime="00:01:23.54" />
                    <SPLIT distance="150" swimtime="00:02:08.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="254" reactiontime="+83" swimtime="00:06:09.83" resultid="2151" heatid="9179" lane="5" entrytime="00:06:12.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:25.76" />
                    <SPLIT distance="150" swimtime="00:02:13.02" />
                    <SPLIT distance="200" swimtime="00:03:00.52" />
                    <SPLIT distance="250" swimtime="00:03:47.47" />
                    <SPLIT distance="300" swimtime="00:04:35.41" />
                    <SPLIT distance="350" swimtime="00:05:23.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-11-16" firstname="Karolina" gender="F" lastname="Głuszkowska" nation="POL" athleteid="2124">
              <RESULTS>
                <RESULT eventid="1187" points="406" reactiontime="+67" swimtime="00:00:34.64" resultid="2125" heatid="8953" lane="3" entrytime="00:00:32.48" />
                <RESULT eventid="1423" points="396" reactiontime="+68" swimtime="00:00:33.18" resultid="2126" heatid="9058" lane="3" entrytime="00:00:32.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-18" firstname="Marcin" gender="M" lastname="Jabłoński" nation="POL" athleteid="2090">
              <RESULTS>
                <RESULT eventid="1079" points="609" reactiontime="+64" swimtime="00:00:23.89" resultid="2091" heatid="8915" lane="5" entrytime="00:00:23.20" />
                <RESULT eventid="1113" points="550" reactiontime="+67" swimtime="00:02:13.79" resultid="2092" heatid="8931" lane="4" entrytime="00:02:09.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                    <SPLIT distance="100" swimtime="00:01:02.87" />
                    <SPLIT distance="150" swimtime="00:01:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="517" reactiontime="+62" swimtime="00:00:27.67" resultid="2093" heatid="8965" lane="2" entrytime="00:00:27.18" />
                <RESULT eventid="1273" points="629" reactiontime="+69" swimtime="00:00:52.43" resultid="2094" heatid="9000" lane="5" entrytime="00:00:51.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="576" reactiontime="+73" swimtime="00:00:26.20" resultid="2095" heatid="9073" lane="3" entrytime="00:00:25.32" />
                <RESULT eventid="1508" points="619" reactiontime="+74" swimtime="00:01:56.57" resultid="2096" heatid="9106" lane="4" entrytime="00:01:53.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                    <SPLIT distance="100" swimtime="00:00:57.44" />
                    <SPLIT distance="150" swimtime="00:01:27.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="611" reactiontime="+70" swimtime="00:00:57.06" resultid="2097" heatid="9137" lane="5" entrytime="00:00:55.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1744" points="581" reactiontime="+70" swimtime="00:04:14.30" resultid="2098" heatid="9192" lane="4" entrytime="00:04:12.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="100" swimtime="00:00:59.71" />
                    <SPLIT distance="150" swimtime="00:01:31.79" />
                    <SPLIT distance="200" swimtime="00:02:04.33" />
                    <SPLIT distance="250" swimtime="00:02:37.16" />
                    <SPLIT distance="300" swimtime="00:03:10.24" />
                    <SPLIT distance="350" swimtime="00:03:42.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-09" firstname="Bartosz" gender="M" lastname="Turla" nation="POL" athleteid="2127">
              <RESULTS>
                <RESULT eventid="1113" points="215" reactiontime="+92" swimtime="00:03:02.93" resultid="2128" heatid="8929" lane="8" entrytime="00:02:32.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:29.83" />
                    <SPLIT distance="150" swimtime="00:02:20.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="255" reactiontime="+101" swimtime="00:22:19.63" resultid="2129" heatid="8945" lane="1" entrytime="00:21:28.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:15.83" />
                    <SPLIT distance="150" swimtime="00:01:57.13" />
                    <SPLIT distance="200" swimtime="00:02:39.49" />
                    <SPLIT distance="250" swimtime="00:03:22.82" />
                    <SPLIT distance="300" swimtime="00:04:05.98" />
                    <SPLIT distance="350" swimtime="00:04:50.23" />
                    <SPLIT distance="400" swimtime="00:05:35.53" />
                    <SPLIT distance="450" swimtime="00:06:20.75" />
                    <SPLIT distance="500" swimtime="00:07:06.78" />
                    <SPLIT distance="550" swimtime="00:07:52.88" />
                    <SPLIT distance="600" swimtime="00:08:38.37" />
                    <SPLIT distance="650" swimtime="00:09:23.83" />
                    <SPLIT distance="700" swimtime="00:10:08.90" />
                    <SPLIT distance="750" swimtime="00:10:53.76" />
                    <SPLIT distance="800" swimtime="00:11:39.12" />
                    <SPLIT distance="850" swimtime="00:12:24.44" />
                    <SPLIT distance="900" swimtime="00:13:10.03" />
                    <SPLIT distance="950" swimtime="00:13:55.74" />
                    <SPLIT distance="1000" swimtime="00:14:41.54" />
                    <SPLIT distance="1050" swimtime="00:15:27.34" />
                    <SPLIT distance="1100" swimtime="00:16:13.60" />
                    <SPLIT distance="1150" swimtime="00:16:59.35" />
                    <SPLIT distance="1200" swimtime="00:17:45.52" />
                    <SPLIT distance="1250" swimtime="00:18:31.28" />
                    <SPLIT distance="1300" swimtime="00:19:16.87" />
                    <SPLIT distance="1350" swimtime="00:20:02.96" />
                    <SPLIT distance="1400" swimtime="00:20:49.56" />
                    <SPLIT distance="1450" swimtime="00:21:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="293" reactiontime="+88" swimtime="00:01:07.61" resultid="2130" heatid="8993" lane="2" entrytime="00:01:05.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="219" reactiontime="+89" swimtime="00:01:23.98" resultid="2131" heatid="9015" lane="5" entrytime="00:01:14.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="234" reactiontime="+94" swimtime="00:01:30.24" resultid="2132" heatid="9047" lane="1" entrytime="00:01:30.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="288" reactiontime="+88" swimtime="00:02:30.36" resultid="2133" heatid="9102" lane="9" entrytime="00:02:20.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                    <SPLIT distance="150" swimtime="00:01:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="217" reactiontime="+94" swimtime="00:00:41.99" resultid="2134" heatid="9166" lane="7" entrytime="00:00:38.76" />
                <RESULT eventid="1744" points="271" reactiontime="+95" swimtime="00:05:27.60" resultid="2135" heatid="9188" lane="7" entrytime="00:05:15.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:11.74" />
                    <SPLIT distance="150" swimtime="00:01:51.17" />
                    <SPLIT distance="200" swimtime="00:02:32.22" />
                    <SPLIT distance="250" swimtime="00:03:15.45" />
                    <SPLIT distance="300" swimtime="00:03:58.84" />
                    <SPLIT distance="350" swimtime="00:04:43.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-06-23" firstname="Ireneusz" gender="M" lastname="Stachecki" nation="POL" athleteid="2157">
              <RESULTS>
                <RESULT eventid="1079" points="218" reactiontime="+94" swimtime="00:00:33.62" resultid="2158" heatid="8900" lane="2" entrytime="00:00:33.15" />
                <RESULT eventid="1165" points="185" reactiontime="+96" swimtime="00:24:49.93" resultid="2159" heatid="8942" lane="3" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:26.16" />
                    <SPLIT distance="150" swimtime="00:02:14.80" />
                    <SPLIT distance="200" swimtime="00:03:03.46" />
                    <SPLIT distance="250" swimtime="00:03:52.72" />
                    <SPLIT distance="300" swimtime="00:04:42.11" />
                    <SPLIT distance="350" swimtime="00:05:32.30" />
                    <SPLIT distance="400" swimtime="00:06:22.34" />
                    <SPLIT distance="450" swimtime="00:07:12.37" />
                    <SPLIT distance="500" swimtime="00:08:02.41" />
                    <SPLIT distance="550" swimtime="00:08:53.16" />
                    <SPLIT distance="600" swimtime="00:09:42.09" />
                    <SPLIT distance="650" swimtime="00:10:31.96" />
                    <SPLIT distance="700" swimtime="00:11:22.17" />
                    <SPLIT distance="750" swimtime="00:12:12.99" />
                    <SPLIT distance="800" swimtime="00:13:03.21" />
                    <SPLIT distance="850" swimtime="00:13:53.49" />
                    <SPLIT distance="900" swimtime="00:14:44.01" />
                    <SPLIT distance="950" swimtime="00:15:34.13" />
                    <SPLIT distance="1000" swimtime="00:16:24.65" />
                    <SPLIT distance="1050" swimtime="00:17:15.51" />
                    <SPLIT distance="1100" swimtime="00:18:06.37" />
                    <SPLIT distance="1150" swimtime="00:18:56.63" />
                    <SPLIT distance="1200" swimtime="00:19:47.76" />
                    <SPLIT distance="1250" swimtime="00:20:37.93" />
                    <SPLIT distance="1300" swimtime="00:21:28.28" />
                    <SPLIT distance="1350" swimtime="00:22:19.26" />
                    <SPLIT distance="1400" swimtime="00:23:10.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="208" reactiontime="+91" swimtime="00:01:15.79" resultid="2160" heatid="8988" lane="4" entrytime="00:01:18.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-11-21" firstname="Tomasz" gender="M" lastname="Stankowski" nation="POL" athleteid="2111">
              <RESULTS>
                <RESULT eventid="1307" points="547" reactiontime="+68" swimtime="00:01:01.93" resultid="2113" heatid="9020" lane="5" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="582" reactiontime="+68" swimtime="00:00:26.10" resultid="2114" heatid="9073" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1613" points="585" reactiontime="+62" swimtime="00:00:57.90" resultid="2115" heatid="9136" lane="4" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="575" reactiontime="+68" swimtime="00:00:30.36" resultid="2116" heatid="9172" lane="2" entrytime="00:00:31.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-11-15" firstname="Aleksander" gender="M" lastname="Sęczkowski" nation="POL" athleteid="2117">
              <RESULTS>
                <RESULT eventid="1079" points="378" reactiontime="+72" swimtime="00:00:28.01" resultid="2118" heatid="8910" lane="0" entrytime="00:00:27.36" />
                <RESULT eventid="1205" points="343" reactiontime="+66" swimtime="00:00:31.73" resultid="2119" heatid="8963" lane="6" entrytime="00:00:30.51" />
                <RESULT eventid="1307" points="401" reactiontime="+68" swimtime="00:01:08.65" resultid="2120" heatid="9018" lane="4" entrytime="00:01:08.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="371" reactiontime="+58" swimtime="00:01:08.07" resultid="2121" heatid="9085" lane="7" entrytime="00:01:09.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="329" reactiontime="+64" swimtime="00:01:10.15" resultid="2122" heatid="9135" lane="4" entrytime="00:01:04.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="394" reactiontime="+62" swimtime="00:00:34.43" resultid="2123" heatid="9170" lane="5" entrytime="00:00:34.29" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-19" firstname="Łukasz" gender="M" lastname="Dziubaty" nation="POL" athleteid="2105">
              <RESULTS>
                <RESULT eventid="1165" points="226" reactiontime="+116" swimtime="00:23:15.59" resultid="2106" heatid="8943" lane="3" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:22.14" />
                    <SPLIT distance="150" swimtime="00:02:06.20" />
                    <SPLIT distance="200" swimtime="00:02:51.58" />
                    <SPLIT distance="250" swimtime="00:03:38.60" />
                    <SPLIT distance="300" swimtime="00:04:24.66" />
                    <SPLIT distance="350" swimtime="00:05:10.50" />
                    <SPLIT distance="400" swimtime="00:05:56.97" />
                    <SPLIT distance="450" swimtime="00:06:43.46" />
                    <SPLIT distance="500" swimtime="00:07:29.88" />
                    <SPLIT distance="550" swimtime="00:08:16.93" />
                    <SPLIT distance="600" swimtime="00:09:04.12" />
                    <SPLIT distance="650" swimtime="00:09:51.29" />
                    <SPLIT distance="700" swimtime="00:10:39.00" />
                    <SPLIT distance="750" swimtime="00:11:26.48" />
                    <SPLIT distance="800" swimtime="00:12:13.92" />
                    <SPLIT distance="850" swimtime="00:13:01.43" />
                    <SPLIT distance="900" swimtime="00:13:48.83" />
                    <SPLIT distance="950" swimtime="00:14:36.53" />
                    <SPLIT distance="1000" swimtime="00:15:23.68" />
                    <SPLIT distance="1050" swimtime="00:16:10.74" />
                    <SPLIT distance="1100" swimtime="00:16:57.97" />
                    <SPLIT distance="1150" swimtime="00:17:45.57" />
                    <SPLIT distance="1200" swimtime="00:18:33.02" />
                    <SPLIT distance="1250" swimtime="00:19:20.56" />
                    <SPLIT distance="1300" swimtime="00:20:07.65" />
                    <SPLIT distance="1350" swimtime="00:20:54.31" />
                    <SPLIT distance="1400" swimtime="00:21:42.87" />
                    <SPLIT distance="1450" swimtime="00:22:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="273" reactiontime="+88" swimtime="00:01:09.26" resultid="2107" heatid="8991" lane="3" entrytime="00:01:09.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="186" reactiontime="+91" swimtime="00:00:38.18" resultid="2108" heatid="9065" lane="6" entrytime="00:00:33.99" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="2109" heatid="9133" lane="8" entrytime="00:01:16.37" />
                <RESULT eventid="1744" points="234" reactiontime="+97" swimtime="00:05:44.04" resultid="2110" heatid="9188" lane="1" entrytime="00:05:15.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                    <SPLIT distance="150" swimtime="00:02:00.16" />
                    <SPLIT distance="200" swimtime="00:02:43.94" />
                    <SPLIT distance="250" swimtime="00:03:28.76" />
                    <SPLIT distance="300" swimtime="00:04:14.46" />
                    <SPLIT distance="350" swimtime="00:04:59.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-02-29" firstname="Adrian" gender="M" lastname="Roszak" nation="POL" athleteid="2136">
              <RESULTS>
                <RESULT eventid="1079" points="578" reactiontime="+76" swimtime="00:00:24.31" resultid="2137" heatid="8915" lane="3" entrytime="00:00:23.50" />
                <RESULT eventid="1273" points="578" reactiontime="+83" swimtime="00:00:53.92" resultid="2138" heatid="9000" lane="2" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="481" reactiontime="+82" swimtime="00:00:27.81" resultid="2139" heatid="9072" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1613" points="528" reactiontime="+85" swimtime="00:00:59.90" resultid="2140" heatid="9136" lane="5" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-03-14" firstname="Tadeusz" gender="M" lastname="Gołembiewski" nation="POL" athleteid="2141">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="2142" heatid="8912" lane="6" entrytime="00:00:26.32" />
                <RESULT eventid="1273" points="531" reactiontime="+87" swimtime="00:00:55.48" resultid="2143" heatid="8999" lane="2" entrytime="00:00:57.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="431" reactiontime="+87" swimtime="00:00:28.86" resultid="2144" heatid="9072" lane="7" entrytime="00:00:27.28" />
                <RESULT eventid="1508" points="495" reactiontime="+83" swimtime="00:02:05.59" resultid="2145" heatid="9105" lane="4" entrytime="00:02:05.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                    <SPLIT distance="100" swimtime="00:01:00.81" />
                    <SPLIT distance="150" swimtime="00:01:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2146" heatid="9192" lane="8" entrytime="00:04:32.76" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="568" reactiontime="+59" swimtime="00:01:49.28" resultid="2163" heatid="9035" lane="5" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                    <SPLIT distance="100" swimtime="00:00:57.91" />
                    <SPLIT distance="150" swimtime="00:01:25.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2090" number="1" reactiontime="+59" />
                    <RELAYPOSITION athleteid="2111" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="2141" number="3" reactiontime="+156" />
                    <RELAYPOSITION athleteid="2136" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1548" points="609" reactiontime="+68" swimtime="00:01:37.42" resultid="2164" heatid="9112" lane="5" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.08" />
                    <SPLIT distance="100" swimtime="00:00:50.10" />
                    <SPLIT distance="150" swimtime="00:01:13.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2111" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2141" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="2090" number="3" reactiontime="+164" />
                    <RELAYPOSITION athleteid="2136" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="253" reactiontime="+67" swimtime="00:02:22.93" resultid="2165" heatid="9033" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:14.21" />
                    <SPLIT distance="150" swimtime="00:01:51.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2152" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="2099" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2105" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2127" number="4" reactiontime="+105" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="304" reactiontime="+94" swimtime="00:02:02.80" resultid="2166" heatid="9111" lane="0" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:01:01.32" />
                    <SPLIT distance="150" swimtime="00:01:32.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2152" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="2099" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2105" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="2127" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="RZ" clubid="4228" name="Uks Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michaslik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="4279">
              <RESULTS>
                <RESULT eventid="1079" points="447" reactiontime="+80" swimtime="00:00:26.48" resultid="4280" heatid="8904" lane="8" entrytime="00:00:30.36" />
                <RESULT eventid="1113" points="367" reactiontime="+90" swimtime="00:02:33.04" resultid="4281" heatid="8926" lane="1" entrytime="00:02:50.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:57.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="455" reactiontime="+82" swimtime="00:00:58.40" resultid="4282" heatid="8994" lane="8" entrytime="00:01:04.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="409" reactiontime="+81" swimtime="00:01:08.20" resultid="4283" heatid="9016" lane="6" entrytime="00:01:12.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="416" reactiontime="+79" swimtime="00:00:29.19" resultid="4284" heatid="9066" lane="7" entrytime="00:00:32.64" />
                <RESULT eventid="1508" points="433" reactiontime="+82" swimtime="00:02:11.28" resultid="4285" heatid="9101" lane="4" entrytime="00:02:21.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="100" swimtime="00:01:02.48" />
                    <SPLIT distance="150" swimtime="00:01:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="358" reactiontime="+84" swimtime="00:01:08.21" resultid="4286" heatid="9132" lane="2" entrytime="00:01:20.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="405" reactiontime="+79" swimtime="00:00:34.12" resultid="4287" heatid="9169" lane="9" entrytime="00:00:36.28" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-04-09" firstname="Zbigniew" gender="M" lastname="Ramos" nation="POL" athleteid="4288">
              <RESULTS>
                <RESULT eventid="1307" points="270" reactiontime="+93" swimtime="00:01:18.29" resultid="4289" heatid="9013" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="275" reactiontime="+96" swimtime="00:01:25.43" resultid="4290" heatid="9049" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="253" reactiontime="+94" swimtime="00:00:34.44" resultid="4291" heatid="9065" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="4292" heatid="9167" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-17" firstname="Sławek" gender="M" lastname="Kowalski" nation="POL" athleteid="4229">
              <RESULTS>
                <RESULT eventid="1079" points="393" reactiontime="+81" swimtime="00:00:27.65" resultid="4230" heatid="8903" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1113" points="353" reactiontime="+78" swimtime="00:02:35.03" resultid="4231" heatid="8927" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="150" swimtime="00:01:57.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="357" reactiontime="+68" swimtime="00:02:49.77" resultid="4232" heatid="8976" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:18.59" />
                    <SPLIT distance="150" swimtime="00:02:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="354" reactiontime="+73" swimtime="00:01:11.58" resultid="4233" heatid="9016" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="386" reactiontime="+70" swimtime="00:01:16.36" resultid="4234" heatid="9051" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="334" reactiontime="+81" swimtime="00:00:31.41" resultid="4235" heatid="9066" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1681" points="376" reactiontime="+73" swimtime="00:00:34.98" resultid="4236" heatid="9171" lane="0" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-04-24" firstname="Renata" gender="F" lastname="Osmala" nation="POL" athleteid="4244">
              <RESULTS>
                <RESULT eventid="1147" points="375" reactiontime="+93" swimtime="00:11:04.62" resultid="4245" heatid="8939" lane="1" entrytime="00:11:20.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:01:14.61" />
                    <SPLIT distance="150" swimtime="00:01:54.99" />
                    <SPLIT distance="200" swimtime="00:02:35.71" />
                    <SPLIT distance="250" swimtime="00:03:16.83" />
                    <SPLIT distance="300" swimtime="00:03:58.19" />
                    <SPLIT distance="350" swimtime="00:04:39.64" />
                    <SPLIT distance="400" swimtime="00:05:21.30" />
                    <SPLIT distance="450" swimtime="00:06:03.46" />
                    <SPLIT distance="500" swimtime="00:06:46.09" />
                    <SPLIT distance="550" swimtime="00:07:28.77" />
                    <SPLIT distance="600" swimtime="00:08:11.89" />
                    <SPLIT distance="650" swimtime="00:08:55.54" />
                    <SPLIT distance="700" swimtime="00:09:39.18" />
                    <SPLIT distance="750" swimtime="00:10:22.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="304" reactiontime="+69" swimtime="00:00:38.15" resultid="4246" heatid="8951" lane="8" entrytime="00:00:38.60" />
                <RESULT eventid="1290" points="333" reactiontime="+84" swimtime="00:01:21.76" resultid="4247" heatid="9005" lane="7" entrytime="00:01:22.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="355" reactiontime="+84" swimtime="00:01:28.06" resultid="4248" heatid="9041" lane="6" entrytime="00:01:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="333" reactiontime="+69" swimtime="00:01:19.35" resultid="4249" heatid="9077" lane="9" entrytime="00:01:22.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="352" reactiontime="+78" swimtime="00:02:48.75" resultid="4250" heatid="9140" lane="4" entrytime="00:02:50.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                    <SPLIT distance="100" swimtime="00:01:22.55" />
                    <SPLIT distance="150" swimtime="00:02:06.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="395" reactiontime="+84" swimtime="00:05:19.56" resultid="4251" heatid="9181" lane="8" entrytime="00:05:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:16.17" />
                    <SPLIT distance="150" swimtime="00:01:56.99" />
                    <SPLIT distance="200" swimtime="00:02:38.01" />
                    <SPLIT distance="250" swimtime="00:03:19.16" />
                    <SPLIT distance="300" swimtime="00:04:00.20" />
                    <SPLIT distance="350" swimtime="00:04:40.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-15" firstname="Paweł" gender="M" lastname="Nowak" nation="POL" athleteid="4268">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="4269" heatid="8897" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1205" points="222" reactiontime="+67" swimtime="00:00:36.67" resultid="4270" heatid="8957" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1307" points="265" reactiontime="+81" swimtime="00:01:18.85" resultid="4271" heatid="9011" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="257" reactiontime="+81" swimtime="00:00:34.27" resultid="4272" heatid="9062" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="4273" heatid="9081" lane="5" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="4261">
              <RESULTS>
                <RESULT eventid="1062" points="394" reactiontime="+92" swimtime="00:00:31.69" resultid="4262" heatid="8890" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1256" points="368" reactiontime="+96" swimtime="00:01:11.14" resultid="4263" heatid="8983" lane="0" entrytime="00:01:10.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="346" reactiontime="+87" swimtime="00:01:20.71" resultid="4264" heatid="9005" lane="5" entrytime="00:01:21.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="297" reactiontime="+78" swimtime="00:00:36.52" resultid="4265" heatid="9057" lane="9" entrytime="00:00:37.20" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="4266" heatid="9076" lane="6" entrytime="00:01:25.00" />
                <RESULT eventid="1595" points="248" reactiontime="+86" swimtime="00:01:26.91" resultid="4267" heatid="9125" lane="2" entrytime="00:01:32.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="4237">
              <RESULTS>
                <RESULT eventid="1079" points="291" reactiontime="+81" swimtime="00:00:30.57" resultid="4238" heatid="8905" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1165" points="253" reactiontime="+89" swimtime="00:22:23.18" resultid="4239" heatid="8944" lane="1" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="150" swimtime="00:01:56.39" />
                    <SPLIT distance="200" swimtime="00:02:38.70" />
                    <SPLIT distance="250" swimtime="00:03:21.26" />
                    <SPLIT distance="300" swimtime="00:04:04.95" />
                    <SPLIT distance="350" swimtime="00:04:48.21" />
                    <SPLIT distance="400" swimtime="00:05:31.96" />
                    <SPLIT distance="450" swimtime="00:06:16.68" />
                    <SPLIT distance="500" swimtime="00:07:01.91" />
                    <SPLIT distance="550" swimtime="00:07:47.81" />
                    <SPLIT distance="600" swimtime="00:08:33.60" />
                    <SPLIT distance="650" swimtime="00:09:20.47" />
                    <SPLIT distance="700" swimtime="00:10:06.87" />
                    <SPLIT distance="750" swimtime="00:10:52.88" />
                    <SPLIT distance="800" swimtime="00:11:39.04" />
                    <SPLIT distance="850" swimtime="00:12:25.60" />
                    <SPLIT distance="900" swimtime="00:13:12.21" />
                    <SPLIT distance="950" swimtime="00:13:58.11" />
                    <SPLIT distance="1000" swimtime="00:14:44.74" />
                    <SPLIT distance="1050" swimtime="00:15:31.15" />
                    <SPLIT distance="1100" swimtime="00:16:17.33" />
                    <SPLIT distance="1150" swimtime="00:17:04.38" />
                    <SPLIT distance="1200" swimtime="00:17:51.21" />
                    <SPLIT distance="1250" swimtime="00:18:37.76" />
                    <SPLIT distance="1300" swimtime="00:19:24.51" />
                    <SPLIT distance="1350" swimtime="00:20:10.83" />
                    <SPLIT distance="1400" swimtime="00:20:57.71" />
                    <SPLIT distance="1450" swimtime="00:21:42.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="312" reactiontime="+78" swimtime="00:01:06.25" resultid="4240" heatid="8992" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="289" reactiontime="+81" swimtime="00:02:30.26" resultid="4241" heatid="9100" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="4242" heatid="9119" lane="8" entrytime="00:06:40.00" />
                <RESULT eventid="1744" points="271" reactiontime="+83" swimtime="00:05:27.95" resultid="4243" heatid="9187" lane="6" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:51.61" />
                    <SPLIT distance="200" swimtime="00:02:32.88" />
                    <SPLIT distance="250" swimtime="00:03:15.06" />
                    <SPLIT distance="300" swimtime="00:03:57.38" />
                    <SPLIT distance="350" swimtime="00:04:38.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="Szklarz" nation="POL" athleteid="4274">
              <RESULTS>
                <RESULT eventid="1079" points="368" reactiontime="+74" swimtime="00:00:28.26" resultid="4275" heatid="8906" lane="9" entrytime="00:00:29.50" />
                <RESULT eventid="1205" points="264" reactiontime="+70" swimtime="00:00:34.60" resultid="4276" heatid="8959" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1440" points="342" reactiontime="+82" swimtime="00:00:31.16" resultid="4277" heatid="9066" lane="3" entrytime="00:00:32.50" />
                <RESULT eventid="1681" points="348" reactiontime="+81" swimtime="00:00:35.89" resultid="4278" heatid="9168" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="4252">
              <RESULTS>
                <RESULT eventid="1062" points="365" reactiontime="+82" swimtime="00:00:32.50" resultid="4253" heatid="8890" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="1096" points="336" reactiontime="+81" swimtime="00:02:55.15" resultid="4254" heatid="8919" lane="8" entrytime="00:03:03.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:22.73" />
                    <SPLIT distance="150" swimtime="00:02:13.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="4255" heatid="8982" lane="5" entrytime="00:01:11.50" />
                <RESULT eventid="1290" points="346" reactiontime="+80" swimtime="00:01:20.69" resultid="4256" heatid="9006" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="340" reactiontime="+80" swimtime="00:01:29.29" resultid="4257" heatid="9040" lane="3" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="251" reactiontime="+81" swimtime="00:00:38.61" resultid="4258" heatid="9057" lane="1" entrytime="00:00:36.75" />
                <RESULT eventid="1595" points="259" reactiontime="+88" swimtime="00:01:25.59" resultid="4259" heatid="9125" lane="5" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="332" reactiontime="+76" swimtime="00:00:41.57" resultid="4260" heatid="9156" lane="3" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="349" reactiontime="+61" swimtime="00:02:08.52" resultid="4295" heatid="9034" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:11.85" />
                    <SPLIT distance="150" swimtime="00:01:42.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4268" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4229" number="2" reactiontime="+12" />
                    <RELAYPOSITION athleteid="4274" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="4279" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="394" reactiontime="+79" swimtime="00:01:52.61" resultid="4296" heatid="9111" lane="1" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="100" swimtime="00:00:54.56" />
                    <SPLIT distance="150" swimtime="00:01:22.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4279" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4274" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4229" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="4288" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="335" reactiontime="+83" swimtime="00:01:58.84" resultid="4293" heatid="8935" lane="0" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:00.99" />
                    <SPLIT distance="150" swimtime="00:01:32.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4229" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="4244" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="4261" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4279" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="316" reactiontime="+74" swimtime="00:02:12.75" resultid="4294" heatid="9175" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:12.22" />
                    <SPLIT distance="150" swimtime="00:01:41.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4244" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4229" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="4279" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="4261" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="DOL" clubid="2620" name="UKS Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www.plywanie-zgorzelec.pl" name="Kondracki Łukasz" phone="693852488" state="DOL" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="2621">
              <RESULTS>
                <RESULT eventid="1079" points="122" reactiontime="+87" swimtime="00:00:40.76" resultid="2622" heatid="8896" lane="2" entrytime="00:00:44.00" />
                <RESULT eventid="1165" points="96" reactiontime="+97" swimtime="00:30:55.89" resultid="2623" heatid="8941" lane="6" entrytime="00:32:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.90" />
                    <SPLIT distance="100" swimtime="00:01:52.63" />
                    <SPLIT distance="150" swimtime="00:02:54.83" />
                    <SPLIT distance="200" swimtime="00:03:55.35" />
                    <SPLIT distance="250" swimtime="00:04:57.75" />
                    <SPLIT distance="300" swimtime="00:05:58.50" />
                    <SPLIT distance="350" swimtime="00:07:00.97" />
                    <SPLIT distance="400" swimtime="00:08:02.07" />
                    <SPLIT distance="450" swimtime="00:09:01.98" />
                    <SPLIT distance="500" swimtime="00:10:02.70" />
                    <SPLIT distance="550" swimtime="00:11:03.58" />
                    <SPLIT distance="600" swimtime="00:12:05.57" />
                    <SPLIT distance="650" swimtime="00:13:07.28" />
                    <SPLIT distance="700" swimtime="00:14:08.98" />
                    <SPLIT distance="750" swimtime="00:15:10.83" />
                    <SPLIT distance="800" swimtime="00:16:13.01" />
                    <SPLIT distance="850" swimtime="00:17:15.63" />
                    <SPLIT distance="900" swimtime="00:18:19.26" />
                    <SPLIT distance="950" swimtime="00:19:21.89" />
                    <SPLIT distance="1000" swimtime="00:20:23.22" />
                    <SPLIT distance="1050" swimtime="00:21:24.89" />
                    <SPLIT distance="1100" swimtime="00:22:27.82" />
                    <SPLIT distance="1150" swimtime="00:23:30.62" />
                    <SPLIT distance="1200" swimtime="00:24:34.00" />
                    <SPLIT distance="1250" swimtime="00:25:37.37" />
                    <SPLIT distance="1300" swimtime="00:26:40.45" />
                    <SPLIT distance="1350" swimtime="00:27:44.40" />
                    <SPLIT distance="1400" swimtime="00:28:48.60" />
                    <SPLIT distance="1450" swimtime="00:29:51.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="93" reactiontime="+85" swimtime="00:00:48.96" resultid="2624" heatid="8956" lane="7" entrytime="00:00:49.93" />
                <RESULT eventid="1341" points="65" reactiontime="+85" swimtime="00:04:28.87" resultid="2625" heatid="9026" lane="9" entrytime="00:04:34.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.15" />
                    <SPLIT distance="100" swimtime="00:02:08.25" />
                    <SPLIT distance="150" swimtime="00:03:20.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="85" reactiontime="+84" swimtime="00:01:50.89" resultid="2626" heatid="9080" lane="3" entrytime="00:01:50.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="91" reactiontime="+95" swimtime="00:08:42.01" resultid="2627" heatid="9117" lane="0" entrytime="00:08:41.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.45" />
                    <SPLIT distance="100" swimtime="00:02:04.39" />
                    <SPLIT distance="150" swimtime="00:03:09.07" />
                    <SPLIT distance="200" swimtime="00:04:12.07" />
                    <SPLIT distance="250" swimtime="00:05:30.47" />
                    <SPLIT distance="300" swimtime="00:06:46.75" />
                    <SPLIT distance="350" swimtime="00:07:45.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="61" reactiontime="+90" swimtime="00:02:03.04" resultid="2628" heatid="9129" lane="6" entrytime="00:02:04.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="94" reactiontime="+82" swimtime="00:03:52.68" resultid="2629" heatid="9144" lane="5" entrytime="00:03:59.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.74" />
                    <SPLIT distance="100" swimtime="00:01:56.76" />
                    <SPLIT distance="150" swimtime="00:02:56.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5069" name="UKS Fala Nieporęt">
          <CONTACT email="bartoszkrawczak@wp.pl" name="Krawczak Bartosz" phone="530077078" />
          <ATHLETES>
            <ATHLETE birthdate="1986-05-14" firstname="Bartosz" gender="M" lastname="Krawczak" nation="POL" athleteid="5070">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="5071" heatid="8914" lane="2" entrytime="00:00:25.50" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="5072" heatid="9000" lane="0" entrytime="00:00:56.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="5073" heatid="9072" lane="0" entrytime="00:00:27.50" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="5074" heatid="9106" lane="2" entrytime="00:01:59.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="5075" heatid="9137" lane="0" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="026" nation="POL" clubid="2198" name="UKS FREGATA Kolbuszowa">
          <CONTACT name="Pietryka" phone="604620876" />
          <ATHLETES>
            <ATHLETE birthdate="1986-07-20" firstname="Bartosz" gender="M" lastname="Pietryka" nation="026" athleteid="2199">
              <RESULTS>
                <RESULT eventid="1165" points="360" reactiontime="+96" swimtime="00:19:54.90" resultid="2200" heatid="8947" lane="6" entrytime="00:19:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:13.32" />
                    <SPLIT distance="150" swimtime="00:01:50.77" />
                    <SPLIT distance="200" swimtime="00:02:29.03" />
                    <SPLIT distance="250" swimtime="00:03:07.94" />
                    <SPLIT distance="300" swimtime="00:03:47.91" />
                    <SPLIT distance="350" swimtime="00:04:27.39" />
                    <SPLIT distance="400" swimtime="00:05:07.55" />
                    <SPLIT distance="450" swimtime="00:05:47.62" />
                    <SPLIT distance="500" swimtime="00:06:28.32" />
                    <SPLIT distance="550" swimtime="00:07:08.37" />
                    <SPLIT distance="600" swimtime="00:07:48.87" />
                    <SPLIT distance="650" swimtime="00:08:29.98" />
                    <SPLIT distance="700" swimtime="00:09:11.11" />
                    <SPLIT distance="750" swimtime="00:09:51.46" />
                    <SPLIT distance="800" swimtime="00:10:31.89" />
                    <SPLIT distance="850" swimtime="00:11:12.10" />
                    <SPLIT distance="900" swimtime="00:11:52.27" />
                    <SPLIT distance="950" swimtime="00:12:31.82" />
                    <SPLIT distance="1000" swimtime="00:13:11.89" />
                    <SPLIT distance="1050" swimtime="00:13:53.06" />
                    <SPLIT distance="1100" swimtime="00:14:33.37" />
                    <SPLIT distance="1150" swimtime="00:15:14.22" />
                    <SPLIT distance="1200" swimtime="00:15:54.52" />
                    <SPLIT distance="1250" swimtime="00:16:35.44" />
                    <SPLIT distance="1300" swimtime="00:17:16.55" />
                    <SPLIT distance="1350" swimtime="00:17:56.87" />
                    <SPLIT distance="1400" swimtime="00:18:36.46" />
                    <SPLIT distance="1450" swimtime="00:19:17.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="2201" heatid="8962" lane="6" entrytime="00:00:31.20" entrycourse="SCM" />
                <RESULT eventid="1341" points="362" reactiontime="+87" swimtime="00:02:32.29" resultid="2202" heatid="9030" lane="7" entrytime="00:02:25.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                    <SPLIT distance="100" swimtime="00:01:07.05" />
                    <SPLIT distance="150" swimtime="00:01:45.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="2203" heatid="9071" lane="2" entrytime="00:00:27.90" entrycourse="SCM" />
                <RESULT eventid="1578" points="357" reactiontime="+93" swimtime="00:05:31.70" resultid="2204" heatid="9121" lane="5" entrytime="00:05:25.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:08.47" />
                    <SPLIT distance="150" swimtime="00:01:52.98" />
                    <SPLIT distance="200" swimtime="00:02:34.36" />
                    <SPLIT distance="250" swimtime="00:03:24.05" />
                    <SPLIT distance="300" swimtime="00:04:14.68" />
                    <SPLIT distance="350" swimtime="00:04:54.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="436" reactiontime="+86" swimtime="00:01:03.86" resultid="2205" heatid="9136" lane="2" entrytime="00:01:01.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2206" heatid="9191" lane="1" entrytime="00:04:45.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-11" firstname="Witold" gender="M" lastname="Rado" nation="026" athleteid="2207">
              <RESULTS>
                <RESULT eventid="1165" points="352" reactiontime="+109" swimtime="00:20:03.04" resultid="2208" heatid="8946" lane="1" entrytime="00:21:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:14.60" />
                    <SPLIT distance="150" swimtime="00:01:54.04" />
                    <SPLIT distance="200" swimtime="00:02:33.90" />
                    <SPLIT distance="250" swimtime="00:03:13.74" />
                    <SPLIT distance="300" swimtime="00:03:53.24" />
                    <SPLIT distance="350" swimtime="00:04:33.36" />
                    <SPLIT distance="400" swimtime="00:05:12.75" />
                    <SPLIT distance="450" swimtime="00:05:53.14" />
                    <SPLIT distance="500" swimtime="00:06:33.64" />
                    <SPLIT distance="550" swimtime="00:07:14.21" />
                    <SPLIT distance="600" swimtime="00:07:54.50" />
                    <SPLIT distance="650" swimtime="00:08:34.79" />
                    <SPLIT distance="700" swimtime="00:09:15.34" />
                    <SPLIT distance="750" swimtime="00:09:56.06" />
                    <SPLIT distance="800" swimtime="00:10:36.90" />
                    <SPLIT distance="850" swimtime="00:11:17.82" />
                    <SPLIT distance="900" swimtime="00:11:58.04" />
                    <SPLIT distance="950" swimtime="00:12:38.27" />
                    <SPLIT distance="1000" swimtime="00:13:19.01" />
                    <SPLIT distance="1050" swimtime="00:13:59.38" />
                    <SPLIT distance="1100" swimtime="00:14:39.86" />
                    <SPLIT distance="1150" swimtime="00:15:21.22" />
                    <SPLIT distance="1200" swimtime="00:16:02.04" />
                    <SPLIT distance="1250" swimtime="00:16:42.65" />
                    <SPLIT distance="1300" swimtime="00:17:23.15" />
                    <SPLIT distance="1350" swimtime="00:18:03.76" />
                    <SPLIT distance="1400" swimtime="00:18:43.68" />
                    <SPLIT distance="1450" swimtime="00:19:24.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="2209" heatid="8960" lane="7" entrytime="00:00:34.10" entrycourse="SCM" />
                <RESULT eventid="1341" points="333" reactiontime="+99" swimtime="00:02:36.57" resultid="2210" heatid="9029" lane="4" entrytime="00:02:40.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:01:53.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="307" reactiontime="+97" swimtime="00:00:32.29" resultid="2211" heatid="9067" lane="3" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1578" points="335" reactiontime="+103" swimtime="00:05:38.97" resultid="2212" heatid="9121" lane="8" entrytime="00:05:40.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:13.39" />
                    <SPLIT distance="150" swimtime="00:01:58.85" />
                    <SPLIT distance="200" swimtime="00:02:44.19" />
                    <SPLIT distance="250" swimtime="00:03:33.25" />
                    <SPLIT distance="300" swimtime="00:04:21.92" />
                    <SPLIT distance="350" swimtime="00:05:01.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="321" reactiontime="+99" swimtime="00:01:10.68" resultid="2213" heatid="9135" lane="1" entrytime="00:01:07.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2214" heatid="9189" lane="9" entrytime="00:05:10.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02214" nation="POL" clubid="2470" name="UKS JAGIELLONKA Warszawa">
          <CONTACT email="klipson@op.pl" name="Klepko" />
          <ATHLETES>
            <ATHLETE birthdate="1982-06-03" firstname="Piotr" gender="M" lastname="Fuliński" nation="POL" license="102214700157" athleteid="2471">
              <RESULTS>
                <RESULT eventid="1079" points="476" reactiontime="+86" swimtime="00:00:25.94" resultid="2472" heatid="8913" lane="4" entrytime="00:00:25.98" />
                <RESULT eventid="1273" points="472" reactiontime="+89" swimtime="00:00:57.68" resultid="2473" heatid="8999" lane="7" entrytime="00:00:57.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="467" reactiontime="+80" swimtime="00:02:08.02" resultid="2475" heatid="9104" lane="5" entrytime="00:02:09.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.30" />
                    <SPLIT distance="100" swimtime="00:01:00.86" />
                    <SPLIT distance="150" swimtime="00:01:34.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAL" clubid="2630" name="Uks Sp 8 Chrzanów">
          <CONTACT city="Chrzanów" email="abalp@poczta.onet.pl" name="Zabrzański Alfred" phone="692076808" street="Niepodległości 7/46" zip="32-500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="2631">
              <RESULTS>
                <RESULT eventid="1079" points="277" reactiontime="+83" swimtime="00:00:31.05" resultid="2632" heatid="8902" lane="4" entrytime="00:00:31.01" />
                <RESULT eventid="1205" points="164" reactiontime="+76" swimtime="00:00:40.55" resultid="2633" heatid="8957" lane="2" entrytime="00:00:41.50" />
                <RESULT eventid="1273" points="264" reactiontime="+91" swimtime="00:01:10.04" resultid="2634" heatid="8991" lane="0" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="205" reactiontime="+89" swimtime="00:01:34.19" resultid="2635" heatid="9046" lane="8" entrytime="00:01:35.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="2636" heatid="9098" lane="1" entrytime="00:02:48.00" />
                <RESULT eventid="1681" points="190" reactiontime="+89" swimtime="00:00:43.89" resultid="2637" heatid="9163" lane="1" entrytime="00:00:43.50" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2638" heatid="9185" lane="6" entrytime="00:06:14.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02914" nation="POL" region="MAZ" clubid="4619" name="UKS Victoria Józefów">
          <CONTACT email="ali90@o2.pl" name="kowalczyk alicja" />
          <ATHLETES>
            <ATHLETE birthdate="1966-03-01" firstname="Jan" gender="M" lastname="Kośmider" nation="POL" athleteid="4620">
              <RESULTS>
                <RESULT eventid="1113" points="301" reactiontime="+85" swimtime="00:02:43.42" resultid="4621" heatid="8927" lane="2" entrytime="00:02:45.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:19.22" />
                    <SPLIT distance="150" swimtime="00:02:04.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="296" reactiontime="+82" swimtime="00:03:00.68" resultid="4622" heatid="8976" lane="2" entrytime="00:03:02.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:25.08" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="4623" heatid="9014" lane="6" entrytime="00:01:16.88" />
                <RESULT eventid="1406" points="320" reactiontime="+79" swimtime="00:01:21.23" resultid="4624" heatid="9050" lane="4" entrytime="00:01:22.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="4625" heatid="9120" lane="3" entrytime="00:05:55.05" />
                <RESULT eventid="1681" points="352" reactiontime="+79" swimtime="00:00:35.74" resultid="4626" heatid="9170" lane="7" entrytime="00:00:34.55" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="4627" heatid="9189" lane="1" entrytime="00:05:05.09" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" region="SLA" clubid="5831" name="UKS Wodnik 29 Katowice">
          <CONTACT email="skoczyt@gmail.com" name="Skoczylas Tomasz" phone="662297707" />
          <ATHLETES>
            <ATHLETE birthdate="1937-11-14" firstname="Aleksander" gender="M" lastname="Aleksandrowicz" nation="POL" athleteid="5846">
              <RESULTS>
                <RESULT eventid="1079" points="92" reactiontime="+107" swimtime="00:00:44.74" resultid="5847" heatid="8896" lane="7" entrytime="00:00:44.49" />
                <RESULT eventid="1205" points="53" reactiontime="+79" swimtime="00:00:59.10" resultid="5848" heatid="8955" lane="5" entrytime="00:00:55.66" />
                <RESULT eventid="1239" points="56" reactiontime="+110" swimtime="00:05:13.59" resultid="5849" heatid="8972" lane="0" entrytime="00:04:50.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.04" />
                    <SPLIT distance="100" swimtime="00:02:28.88" />
                    <SPLIT distance="150" swimtime="00:03:52.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="58" reactiontime="+87" swimtime="00:02:22.86" resultid="5850" heatid="9044" lane="7" entrytime="00:02:13.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="49" reactiontime="+82" swimtime="00:02:13.09" resultid="5851" heatid="9080" lane="1" entrytime="00:02:01.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="5852" heatid="9160" lane="3" entrytime="00:00:59.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-08-30" firstname="Aleksandra" gender="F" lastname="Kącki" nation="POL" athleteid="5867">
              <RESULTS>
                <RESULT eventid="1062" points="191" reactiontime="+105" swimtime="00:00:40.29" resultid="5868" heatid="8888" lane="0" entrytime="00:00:39.78" />
                <RESULT eventid="1256" points="174" reactiontime="+109" swimtime="00:01:31.25" resultid="5869" heatid="8980" lane="1" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="132" reactiontime="+110" swimtime="00:00:47.86" resultid="5870" heatid="9054" lane="2" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="5871" heatid="9090" lane="0" entrytime="00:03:21.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-15" firstname="Andrzej" gender="M" lastname="Porszke" nation="POL" athleteid="5878">
              <RESULTS>
                <RESULT eventid="1239" points="220" reactiontime="+101" swimtime="00:03:19.51" resultid="5879" heatid="8975" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                    <SPLIT distance="100" swimtime="00:01:32.21" />
                    <SPLIT distance="150" swimtime="00:02:25.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="245" reactiontime="+72" swimtime="00:01:28.85" resultid="5880" heatid="9049" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="267" reactiontime="+100" swimtime="00:00:39.21" resultid="5881" heatid="9166" lane="1" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-09" firstname="Krystyna" gender="F" lastname="Nicpoń" nation="POL" athleteid="5887">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1096" points="80" reactiontime="+98" swimtime="00:04:41.89" resultid="5888" heatid="8916" lane="5" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.49" />
                    <SPLIT distance="100" swimtime="00:02:22.42" />
                    <SPLIT distance="150" swimtime="00:03:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="108" reactiontime="+78" swimtime="00:00:53.77" resultid="5889" heatid="8949" lane="9" entrytime="00:01:00.00" />
                <RESULT comment="Rekord Polski" eventid="1324" points="27" reactiontime="+104" swimtime="00:06:35.51" resultid="5890" heatid="9022" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.31" />
                    <SPLIT distance="100" swimtime="00:03:08.65" />
                    <SPLIT distance="150" swimtime="00:04:52.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1457" points="112" reactiontime="+82" swimtime="00:01:54.11" resultid="5891" heatid="9075" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.84" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1555" points="73" reactiontime="+105" swimtime="00:10:19.84" resultid="5892" heatid="9113" lane="1" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.33" />
                    <SPLIT distance="100" swimtime="00:03:10.88" />
                    <SPLIT distance="150" swimtime="00:04:12.43" />
                    <SPLIT distance="200" swimtime="00:05:15.20" />
                    <SPLIT distance="250" swimtime="00:06:41.83" />
                    <SPLIT distance="300" swimtime="00:08:02.58" />
                    <SPLIT distance="350" swimtime="00:09:10.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="113" reactiontime="+86" swimtime="00:04:06.56" resultid="5893" heatid="9139" lane="0" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.65" />
                    <SPLIT distance="100" swimtime="00:01:57.72" />
                    <SPLIT distance="150" swimtime="00:03:02.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="5843" />
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="5882">
              <RESULTS>
                <RESULT eventid="1079" points="346" reactiontime="+96" swimtime="00:00:28.84" resultid="5883" heatid="8907" lane="3" entrytime="00:00:28.75" />
                <RESULT eventid="1273" points="304" reactiontime="+104" swimtime="00:01:06.82" resultid="5884" heatid="8992" lane="2" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="315" reactiontime="+97" swimtime="00:00:32.01" resultid="5885" heatid="9067" lane="6" entrytime="00:00:31.20" />
                <RESULT eventid="1613" points="261" reactiontime="+107" swimtime="00:01:15.71" resultid="5886" heatid="9133" lane="6" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-19" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="5853">
              <RESULTS>
                <RESULT eventid="1079" points="239" reactiontime="+99" swimtime="00:00:32.62" resultid="5854" heatid="8901" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1273" points="212" reactiontime="+92" swimtime="00:01:15.33" resultid="5855" heatid="8989" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="117" reactiontime="+102" swimtime="00:03:41.45" resultid="5856" heatid="9027" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.66" />
                    <SPLIT distance="100" swimtime="00:01:44.74" />
                    <SPLIT distance="150" swimtime="00:02:46.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="238" reactiontime="+88" swimtime="00:00:35.13" resultid="5857" heatid="9064" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="5858" heatid="9097" lane="7" entrytime="00:02:59.50" />
                <RESULT eventid="1613" points="160" reactiontime="+96" swimtime="00:01:29.14" resultid="5859" heatid="9131" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="160" reactiontime="+105" swimtime="00:06:30.58" resultid="5860" heatid="9184" lane="1" entrytime="00:06:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:30.49" />
                    <SPLIT distance="150" swimtime="00:02:22.92" />
                    <SPLIT distance="200" swimtime="00:03:15.43" />
                    <SPLIT distance="250" swimtime="00:04:06.29" />
                    <SPLIT distance="300" swimtime="00:04:58.12" />
                    <SPLIT distance="350" swimtime="00:05:48.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-07-13" firstname="Szymon" gender="M" lastname="Warwas" nation="POL" athleteid="5872">
              <RESULTS>
                <RESULT eventid="1079" points="634" reactiontime="+64" swimtime="00:00:23.58" resultid="5873" heatid="8915" lane="4" entrytime="00:00:23.16" />
                <RESULT eventid="1205" points="505" reactiontime="+72" swimtime="00:00:27.90" resultid="5874" heatid="8965" lane="8" entrytime="00:00:27.90" />
                <RESULT eventid="1273" points="639" reactiontime="+64" swimtime="00:00:52.17" resultid="5875" heatid="9000" lane="4" entrytime="00:00:50.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="635" reactiontime="+67" swimtime="00:00:25.36" resultid="5876" heatid="9073" lane="6" entrytime="00:00:25.42" />
                <RESULT eventid="1613" points="609" reactiontime="+69" swimtime="00:00:57.12" resultid="5877" heatid="9137" lane="3" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="5861">
              <RESULTS>
                <RESULT eventid="1113" points="243" reactiontime="+87" swimtime="00:02:55.57" resultid="5862" heatid="8926" lane="0" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:20.24" />
                    <SPLIT distance="150" swimtime="00:02:08.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="311" reactiontime="+90" swimtime="00:02:57.64" resultid="5863" heatid="8977" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                    <SPLIT distance="150" swimtime="00:02:11.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="5864" heatid="9014" lane="3" entrytime="00:01:16.50" />
                <RESULT eventid="1406" points="357" reactiontime="+84" swimtime="00:01:18.32" resultid="5865" heatid="9051" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="380" reactiontime="+81" swimtime="00:00:34.85" resultid="5866" heatid="9169" lane="8" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01711" nation="POL" region="11" clubid="2403" name="UKS WODNIK Siemianowice Śląskie" shortname="UKS WODNIK Siemianowice Śląski">
          <CONTACT city="Siemianowice Śląskie" email="vivisektor@interia.pl" name="Małyszek" phone="534039934" state="ŚLĄSK" street="Mikołaja" zip="41-106" />
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="2404">
              <RESULTS>
                <RESULT eventid="1113" points="220" reactiontime="+86" swimtime="00:03:01.38" resultid="2405" heatid="8925" lane="3" entrytime="00:02:59.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:24.82" />
                    <SPLIT distance="150" swimtime="00:02:18.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="257" reactiontime="+88" swimtime="00:22:17.00" resultid="2406" heatid="8944" lane="4" entrytime="00:21:55.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:02:05.77" />
                    <SPLIT distance="200" swimtime="00:02:51.73" />
                    <SPLIT distance="250" swimtime="00:03:37.89" />
                    <SPLIT distance="300" swimtime="00:04:23.38" />
                    <SPLIT distance="350" swimtime="00:05:09.40" />
                    <SPLIT distance="400" swimtime="00:05:54.61" />
                    <SPLIT distance="450" swimtime="00:06:39.49" />
                    <SPLIT distance="500" swimtime="00:07:24.31" />
                    <SPLIT distance="550" swimtime="00:08:09.88" />
                    <SPLIT distance="600" swimtime="00:08:55.46" />
                    <SPLIT distance="650" swimtime="00:09:40.25" />
                    <SPLIT distance="700" swimtime="00:10:26.03" />
                    <SPLIT distance="750" swimtime="00:11:11.43" />
                    <SPLIT distance="800" swimtime="00:11:56.20" />
                    <SPLIT distance="850" swimtime="00:12:40.94" />
                    <SPLIT distance="900" swimtime="00:13:26.39" />
                    <SPLIT distance="950" swimtime="00:14:11.01" />
                    <SPLIT distance="1000" swimtime="00:14:55.33" />
                    <SPLIT distance="1050" swimtime="00:15:40.53" />
                    <SPLIT distance="1100" swimtime="00:16:25.32" />
                    <SPLIT distance="1150" swimtime="00:17:10.68" />
                    <SPLIT distance="1200" swimtime="00:17:54.57" />
                    <SPLIT distance="1250" swimtime="00:18:39.25" />
                    <SPLIT distance="1300" swimtime="00:19:23.32" />
                    <SPLIT distance="1350" swimtime="00:20:08.24" />
                    <SPLIT distance="1400" swimtime="00:20:52.84" />
                    <SPLIT distance="1450" swimtime="00:21:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="2407" heatid="9027" lane="4" entrytime="00:03:15.60" />
                <RESULT eventid="1508" points="222" reactiontime="+90" swimtime="00:02:43.89" resultid="2408" heatid="9098" lane="4" entrytime="00:02:41.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                    <SPLIT distance="100" swimtime="00:01:18.30" />
                    <SPLIT distance="150" swimtime="00:02:01.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="205" reactiontime="+87" swimtime="00:06:39.04" resultid="2409" heatid="9119" lane="5" entrytime="00:06:25.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                    <SPLIT distance="100" swimtime="00:01:36.47" />
                    <SPLIT distance="150" swimtime="00:02:27.64" />
                    <SPLIT distance="200" swimtime="00:03:20.58" />
                    <SPLIT distance="250" swimtime="00:04:16.28" />
                    <SPLIT distance="300" swimtime="00:05:12.26" />
                    <SPLIT distance="350" swimtime="00:05:56.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="2410" heatid="9132" lane="8" entrytime="00:01:22.60" />
                <RESULT eventid="1744" points="219" reactiontime="+98" swimtime="00:05:51.78" resultid="2411" heatid="9187" lane="0" entrytime="00:05:36.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                    <SPLIT distance="100" swimtime="00:02:05.98" />
                    <SPLIT distance="200" swimtime="00:02:51.30" />
                    <SPLIT distance="250" swimtime="00:03:36.72" />
                    <SPLIT distance="300" swimtime="00:04:23.17" />
                    <SPLIT distance="350" swimtime="00:05:08.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" nation="POL" region="WAR" clubid="2932" name="Ursynów Masters">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1942-03-23" firstname="Ryszard" gender="M" lastname="Rybarczyk" nation="POL" athleteid="2951">
              <RESULTS>
                <RESULT eventid="1079" points="118" reactiontime="+92" swimtime="00:00:41.29" resultid="2952" heatid="8897" lane="9" entrytime="00:00:40.89" />
                <RESULT eventid="1205" points="60" reactiontime="+129" swimtime="00:00:56.57" resultid="2953" heatid="8956" lane="0" entrytime="00:00:53.57" />
                <RESULT eventid="1239" reactiontime="+99" status="DNF" swimtime="00:00:00.00" resultid="2954" heatid="8972" lane="3" entrytime="00:03:57.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="130" reactiontime="+124" swimtime="00:01:49.70" resultid="2955" heatid="9045" lane="1" entrytime="00:01:47.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="2956" heatid="9080" lane="0" entrytime="00:02:06.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="2957" heatid="9144" lane="1" entrytime="00:04:32.00" />
                <RESULT eventid="1681" points="122" reactiontime="+98" swimtime="00:00:50.90" resultid="2958" heatid="9162" lane="8" entrytime="00:00:47.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="Nowak" nation="POL" athleteid="2936">
              <RESULTS>
                <RESULT eventid="1113" points="205" reactiontime="+84" swimtime="00:03:05.76" resultid="2937" heatid="8925" lane="9" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:01:33.33" />
                    <SPLIT distance="150" swimtime="00:02:23.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="249" reactiontime="+85" swimtime="00:03:11.38" resultid="2938" heatid="8975" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                    <SPLIT distance="100" swimtime="00:01:29.96" />
                    <SPLIT distance="150" swimtime="00:02:19.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="257" reactiontime="+83" swimtime="00:01:19.61" resultid="2939" heatid="9012" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="287" reactiontime="+80" swimtime="00:01:24.27" resultid="2940" heatid="9049" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="167" reactiontime="+86" swimtime="00:07:06.81" resultid="2941" heatid="9118" lane="3" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.39" />
                    <SPLIT distance="100" swimtime="00:01:45.08" />
                    <SPLIT distance="150" swimtime="00:02:42.25" />
                    <SPLIT distance="200" swimtime="00:03:41.28" />
                    <SPLIT distance="250" swimtime="00:04:35.59" />
                    <SPLIT distance="300" swimtime="00:05:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="332" reactiontime="+89" swimtime="00:00:36.44" resultid="2942" heatid="9168" lane="1" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-06-01" firstname="Robert" gender="M" lastname="Zieliński" nation="POL" athleteid="2959">
              <RESULTS>
                <RESULT eventid="1079" points="235" reactiontime="+85" swimtime="00:00:32.79" resultid="2960" heatid="8902" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="1205" points="143" reactiontime="+75" swimtime="00:00:42.43" resultid="2961" heatid="8958" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="1273" points="245" reactiontime="+88" swimtime="00:01:11.75" resultid="2962" heatid="8989" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="177" reactiontime="+80" swimtime="00:00:38.77" resultid="2963" heatid="9063" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="2964" heatid="9097" lane="6" entrytime="00:02:58.00" />
                <RESULT eventid="1647" points="137" reactiontime="+77" swimtime="00:03:25.52" resultid="2965" heatid="9145" lane="8" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:39.01" />
                    <SPLIT distance="150" swimtime="00:02:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="174" reactiontime="+86" swimtime="00:00:45.16" resultid="2966" heatid="9161" lane="5" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="Rybarczyk" nation="POL" athleteid="2943">
              <RESULTS>
                <RESULT eventid="1079" points="313" reactiontime="+84" swimtime="00:00:29.82" resultid="2944" heatid="8905" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1205" points="158" reactiontime="+77" swimtime="00:00:41.04" resultid="2945" heatid="8957" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1273" points="323" reactiontime="+77" swimtime="00:01:05.47" resultid="2946" heatid="8990" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="262" reactiontime="+80" swimtime="00:00:34.04" resultid="2947" heatid="9064" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1508" points="267" reactiontime="+92" swimtime="00:02:34.31" resultid="2948" heatid="9099" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="150" swimtime="00:01:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="171" reactiontime="+86" swimtime="00:01:27.16" resultid="2949" heatid="9131" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="128" reactiontime="+84" swimtime="00:03:30.24" resultid="2950" heatid="9145" lane="1" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.89" />
                    <SPLIT distance="100" swimtime="00:01:43.05" />
                    <SPLIT distance="150" swimtime="00:02:38.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="204" reactiontime="+69" swimtime="00:02:33.63" resultid="2967" heatid="9033" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:01:52.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2959" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2936" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="2943" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2951" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1548" points="225" reactiontime="+83" swimtime="00:02:15.67" resultid="2968" heatid="9109" lane="5" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:01:46.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2959" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2951" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="2936" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2943" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="031" nation="POL" region="LOD" clubid="3485" name="UTW &quot;Masters&quot; Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1976-09-03" firstname="Arkadiusz" gender="M" lastname="Bilski" nation="POL" license="503105700042" athleteid="3532">
              <RESULTS>
                <RESULT eventid="1205" points="294" reactiontime="+81" swimtime="00:00:33.40" resultid="3533" heatid="8963" lane="0" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1239" points="383" reactiontime="+73" swimtime="00:02:45.78" resultid="3534" heatid="8977" lane="3" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:19.92" />
                    <SPLIT distance="150" swimtime="00:02:03.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="400" reactiontime="+74" swimtime="00:01:15.42" resultid="3535" heatid="9052" lane="5" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="3536" heatid="9085" lane="1" entrytime="00:01:10.00" entrycourse="SCM" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="3537" heatid="9148" lane="7" entrytime="00:02:40.00" entrycourse="SCM" />
                <RESULT eventid="1681" points="396" reactiontime="+67" swimtime="00:00:34.36" resultid="3538" heatid="9171" lane="6" entrytime="00:00:33.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-23" firstname="Tomasz" gender="M" lastname="Cajdler" nation="POL" license="503105700035" athleteid="3578">
              <RESULTS>
                <RESULT eventid="1079" points="245" reactiontime="+103" swimtime="00:00:32.37" resultid="3579" heatid="8901" lane="2" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="222" reactiontime="+94" swimtime="00:01:14.14" resultid="3580" heatid="8990" lane="8" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="131" reactiontime="+79" swimtime="00:00:42.84" resultid="3581" heatid="9062" lane="9" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="1681" points="216" reactiontime="+85" swimtime="00:00:42.08" resultid="3582" heatid="9164" lane="9" entrytime="00:00:42.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-16" firstname="Adrian" gender="M" lastname="Styrzyński" nation="POL" license="503105700033" athleteid="3592">
              <RESULTS>
                <RESULT eventid="1113" points="565" reactiontime="+74" swimtime="00:02:12.56" resultid="3593" heatid="8931" lane="6" entrytime="00:02:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.20" />
                    <SPLIT distance="100" swimtime="00:01:01.71" />
                    <SPLIT distance="150" swimtime="00:01:39.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="606" reactiontime="+74" swimtime="00:00:59.84" resultid="3594" heatid="9021" lane="7" entrytime="00:01:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="594" reactiontime="+74" swimtime="00:01:58.19" resultid="3595" heatid="9106" lane="7" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                    <SPLIT distance="100" swimtime="00:00:58.01" />
                    <SPLIT distance="150" swimtime="00:01:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="3596" heatid="9137" lane="2" entrytime="00:00:57.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-07-18" firstname="Tomasz" gender="M" lastname="Niedżwiedż" nation="POL" license="503105700038" athleteid="3583">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="3584" heatid="8899" lane="3" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1113" points="146" reactiontime="+110" swimtime="00:03:28.05" resultid="3585" heatid="8923" lane="1" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.61" />
                    <SPLIT distance="100" swimtime="00:01:45.50" />
                    <SPLIT distance="150" swimtime="00:02:43.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="3586" heatid="9010" lane="3" entrytime="00:01:35.00" entrycourse="SCM" />
                <RESULT eventid="1341" points="103" reactiontime="+113" swimtime="00:03:51.56" resultid="3587" heatid="9027" lane="0" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.06" />
                    <SPLIT distance="100" swimtime="00:01:49.80" />
                    <SPLIT distance="150" swimtime="00:02:51.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="3588" heatid="9081" lane="9" entrytime="00:01:50.00" entrycourse="SCM" />
                <RESULT eventid="1578" points="137" reactiontime="+112" swimtime="00:07:36.50" resultid="3589" heatid="9117" lane="4" entrytime="00:07:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.64" />
                    <SPLIT distance="100" swimtime="00:01:50.25" />
                    <SPLIT distance="150" swimtime="00:02:51.96" />
                    <SPLIT distance="200" swimtime="00:03:54.61" />
                    <SPLIT distance="250" swimtime="00:04:55.97" />
                    <SPLIT distance="300" swimtime="00:05:57.94" />
                    <SPLIT distance="350" swimtime="00:06:48.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="3590" heatid="9130" lane="7" entrytime="00:01:45.00" entrycourse="SCM" />
                <RESULT eventid="1647" points="97" reactiontime="+101" swimtime="00:03:50.47" resultid="3591" heatid="9145" lane="0" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.24" />
                    <SPLIT distance="100" swimtime="00:01:53.51" />
                    <SPLIT distance="150" swimtime="00:02:52.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105700038" athleteid="3566">
              <RESULTS>
                <RESULT eventid="1239" points="170" reactiontime="+116" swimtime="00:03:37.21" resultid="3567" heatid="8973" lane="2" entrytime="00:03:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                    <SPLIT distance="100" swimtime="00:01:43.36" />
                    <SPLIT distance="150" swimtime="00:02:41.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="3568" heatid="9011" lane="1" entrytime="00:01:30.00" entrycourse="SCM" />
                <RESULT eventid="1406" points="206" reactiontime="+109" swimtime="00:01:34.04" resultid="3569" heatid="9046" lane="2" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="237" reactiontime="+106" swimtime="00:00:40.75" resultid="3570" heatid="9164" lane="6" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-10" firstname="Sonia" gender="F" lastname="Bochyńska" nation="POL" license="503105600046" athleteid="3571">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="3572" heatid="8893" lane="1" entrytime="00:00:28.48" entrycourse="SCM" />
                <RESULT eventid="1187" points="550" reactiontime="+71" swimtime="00:00:31.33" resultid="3573" heatid="8953" lane="4" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1290" points="530" reactiontime="+72" swimtime="00:01:10.04" resultid="3574" heatid="9007" lane="4" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="516" reactiontime="+73" swimtime="00:00:30.39" resultid="3575" heatid="9059" lane="6" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1457" points="508" reactiontime="+69" swimtime="00:01:08.93" resultid="3576" heatid="9078" lane="4" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="502" reactiontime="+74" swimtime="00:02:29.99" resultid="3577" heatid="9141" lane="5" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="150" swimtime="00:01:52.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-08" firstname="Ewa" gender="F" lastname="Zimna-Walendzik" nation="POL" license="503105600019" athleteid="3615">
              <RESULTS>
                <RESULT eventid="1062" points="166" reactiontime="+100" swimtime="00:00:42.26" resultid="3616" heatid="8887" lane="2" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1096" points="125" reactiontime="+95" swimtime="00:04:03.28" resultid="3617" heatid="8917" lane="8" entrytime="00:03:48.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.50" />
                    <SPLIT distance="100" swimtime="00:01:57.38" />
                    <SPLIT distance="150" swimtime="00:03:05.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="144" reactiontime="+97" swimtime="00:01:37.27" resultid="3618" heatid="8979" lane="4" entrytime="00:01:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="149" reactiontime="+98" swimtime="00:01:46.81" resultid="3619" heatid="9002" lane="7" entrytime="00:01:46.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="112" reactiontime="+101" swimtime="00:00:50.46" resultid="3620" heatid="9055" lane="0" entrytime="00:00:49.00" entrycourse="SCM" />
                <RESULT eventid="1491" points="137" reactiontime="+97" swimtime="00:03:34.61" resultid="3621" heatid="9089" lane="6" entrytime="00:03:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="100" swimtime="00:01:40.32" />
                    <SPLIT distance="150" swimtime="00:02:36.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="99" reactiontime="+101" swimtime="00:01:57.68" resultid="3622" heatid="9124" lane="0" entrytime="00:02:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700027" athleteid="3499">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="3500" heatid="8903" lane="1" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1113" points="258" reactiontime="+86" swimtime="00:02:52.08" resultid="3501" heatid="8926" lane="9" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:20.32" />
                    <SPLIT distance="150" swimtime="00:02:13.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="255" reactiontime="+74" swimtime="00:00:35.00" resultid="3502" heatid="8959" lane="5" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1341" points="194" reactiontime="+93" swimtime="00:03:07.45" resultid="3503" heatid="9028" lane="3" entrytime="00:03:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:29.86" />
                    <SPLIT distance="150" swimtime="00:02:19.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="3504" heatid="9082" lane="5" entrytime="00:01:20.00" entrycourse="SCM" />
                <RESULT eventid="1508" points="290" reactiontime="+89" swimtime="00:02:30.11" resultid="3505" heatid="9100" lane="4" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:12.40" />
                    <SPLIT distance="150" swimtime="00:01:51.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="3506" heatid="9147" lane="0" entrytime="00:03:00.00" entrycourse="SCM" />
                <RESULT eventid="1744" points="278" reactiontime="+95" swimtime="00:05:24.98" resultid="3507" heatid="9187" lane="4" entrytime="00:05:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:15.45" />
                    <SPLIT distance="150" swimtime="00:01:55.58" />
                    <SPLIT distance="200" swimtime="00:02:37.32" />
                    <SPLIT distance="250" swimtime="00:03:19.52" />
                    <SPLIT distance="300" swimtime="00:04:01.75" />
                    <SPLIT distance="350" swimtime="00:04:44.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105600018" athleteid="3546">
              <RESULTS>
                <RESULT eventid="1062" points="529" reactiontime="+79" swimtime="00:00:28.72" resultid="3547" heatid="8893" lane="9" entrytime="00:00:29.50" entrycourse="SCM" />
                <RESULT eventid="1187" points="486" reactiontime="+77" swimtime="00:00:32.64" resultid="3548" heatid="8953" lane="7" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT comment="Rekord Polski" eventid="1290" points="511" reactiontime="+87" swimtime="00:01:10.91" resultid="3549" heatid="9007" lane="5" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="480" reactiontime="+70" swimtime="00:01:10.26" resultid="3550" heatid="9078" lane="5" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1555" points="451" reactiontime="+95" swimtime="00:05:38.63" resultid="3551" heatid="9115" lane="6" entrytime="00:05:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:15.92" />
                    <SPLIT distance="150" swimtime="00:02:00.12" />
                    <SPLIT distance="200" swimtime="00:02:42.76" />
                    <SPLIT distance="250" swimtime="00:03:30.65" />
                    <SPLIT distance="300" swimtime="00:04:19.16" />
                    <SPLIT distance="350" swimtime="00:04:59.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="440" reactiontime="+71" swimtime="00:02:36.72" resultid="3552" heatid="9141" lane="7" entrytime="00:02:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:01:56.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="503105700036" athleteid="3597">
              <RESULTS>
                <RESULT eventid="1079" points="470" reactiontime="+91" swimtime="00:00:26.04" resultid="3598" heatid="8914" lane="0" entrytime="00:00:25.95" entrycourse="SCM" />
                <RESULT eventid="1205" points="374" reactiontime="+80" swimtime="00:00:30.84" resultid="3599" heatid="8964" lane="0" entrytime="00:00:29.99" entrycourse="SCM" />
                <RESULT eventid="1474" points="368" reactiontime="+80" swimtime="00:01:08.24" resultid="3600" heatid="9086" lane="7" entrytime="00:01:05.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="415" reactiontime="+86" swimtime="00:00:33.84" resultid="3601" heatid="9170" lane="4" entrytime="00:00:34.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-16" firstname="Krzysztof" gender="M" lastname="Gawłowicz" nation="POL" license="503105700049" athleteid="3612">
              <RESULTS>
                <RESULT eventid="1079" points="548" reactiontime="+68" swimtime="00:00:24.75" resultid="3613" heatid="8914" lane="6" entrytime="00:00:25.00" entrycourse="SCM" />
                <RESULT eventid="1440" points="551" reactiontime="+69" swimtime="00:00:26.58" resultid="3614" heatid="9073" lane="8" entrytime="00:00:26.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-04-11" firstname="Jakub" gender="M" lastname="Jurek" nation="POL" license="503105700047" athleteid="3553">
              <RESULTS>
                <RESULT eventid="1079" points="374" reactiontime="+66" swimtime="00:00:28.10" resultid="3554" heatid="8907" lane="5" entrytime="00:00:28.50" entrycourse="SCM" />
                <RESULT eventid="1113" points="315" reactiontime="+87" swimtime="00:02:41.10" resultid="3555" heatid="8928" lane="0" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:02:05.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="302" reactiontime="+72" swimtime="00:00:33.09" resultid="3556" heatid="8961" lane="7" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1307" points="353" reactiontime="+78" swimtime="00:01:11.67" resultid="3557" heatid="9017" lane="5" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="302" reactiontime="+69" swimtime="00:01:12.87" resultid="3558" heatid="9084" lane="2" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="3559" heatid="9100" lane="1" entrytime="00:02:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-06" firstname="Wojciech" gender="M" lastname="Szymański" nation="POL" license="503105700037" athleteid="3608">
              <RESULTS>
                <RESULT eventid="1165" points="68" reactiontime="+119" swimtime="00:34:32.75" resultid="3609" heatid="8941" lane="9" entrytime="00:36:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.54" />
                    <SPLIT distance="100" swimtime="00:01:53.98" />
                    <SPLIT distance="150" swimtime="00:02:59.06" />
                    <SPLIT distance="200" swimtime="00:04:04.99" />
                    <SPLIT distance="250" swimtime="00:05:12.65" />
                    <SPLIT distance="300" swimtime="00:06:22.73" />
                    <SPLIT distance="350" swimtime="00:07:32.38" />
                    <SPLIT distance="400" swimtime="00:08:42.74" />
                    <SPLIT distance="450" swimtime="00:09:52.72" />
                    <SPLIT distance="500" swimtime="00:11:01.45" />
                    <SPLIT distance="550" swimtime="00:12:10.83" />
                    <SPLIT distance="600" swimtime="00:13:19.94" />
                    <SPLIT distance="650" swimtime="00:14:30.12" />
                    <SPLIT distance="700" swimtime="00:15:37.98" />
                    <SPLIT distance="750" swimtime="00:16:47.42" />
                    <SPLIT distance="800" swimtime="00:17:58.12" />
                    <SPLIT distance="850" swimtime="00:19:07.26" />
                    <SPLIT distance="900" swimtime="00:20:17.87" />
                    <SPLIT distance="950" swimtime="00:21:27.88" />
                    <SPLIT distance="1000" swimtime="00:22:38.80" />
                    <SPLIT distance="1050" swimtime="00:23:49.90" />
                    <SPLIT distance="1100" swimtime="00:25:00.72" />
                    <SPLIT distance="1150" swimtime="00:26:11.85" />
                    <SPLIT distance="1200" swimtime="00:27:22.88" />
                    <SPLIT distance="1250" swimtime="00:28:34.56" />
                    <SPLIT distance="1300" swimtime="00:29:47.50" />
                    <SPLIT distance="1350" swimtime="00:30:59.53" />
                    <SPLIT distance="1400" swimtime="00:32:14.96" />
                    <SPLIT distance="1450" swimtime="00:33:26.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="3610" heatid="9095" lane="1" entrytime="00:04:00.00" entrycourse="SCM" />
                <RESULT eventid="1744" points="66" reactiontime="+106" swimtime="00:08:42.93" resultid="3611" heatid="9182" lane="6" entrytime="00:09:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.84" />
                    <SPLIT distance="100" swimtime="00:01:51.71" />
                    <SPLIT distance="150" swimtime="00:02:56.25" />
                    <SPLIT distance="200" swimtime="00:04:04.01" />
                    <SPLIT distance="250" swimtime="00:05:12.28" />
                    <SPLIT distance="300" swimtime="00:06:21.74" />
                    <SPLIT distance="350" swimtime="00:07:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="3539">
              <RESULTS>
                <RESULT eventid="1096" points="447" reactiontime="+93" swimtime="00:02:39.31" resultid="3540" heatid="8920" lane="7" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:14.80" />
                    <SPLIT distance="150" swimtime="00:02:01.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1324" points="396" reactiontime="+93" swimtime="00:02:42.85" resultid="3541" heatid="9024" lane="5" entrytime="00:02:49.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:16.04" />
                    <SPLIT distance="150" swimtime="00:01:58.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="401" reactiontime="+98" swimtime="00:01:24.50" resultid="3542" heatid="9042" lane="1" entrytime="00:01:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="433" reactiontime="+87" swimtime="00:00:32.21" resultid="3543" heatid="9058" lane="4" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1595" points="444" reactiontime="+95" swimtime="00:01:11.56" resultid="3544" heatid="9127" lane="2" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="390" reactiontime="+94" swimtime="00:00:39.41" resultid="3545" heatid="9158" lane="6" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" license="503105600029" athleteid="3520">
              <RESULTS>
                <RESULT eventid="1062" points="374" reactiontime="+75" swimtime="00:00:32.23" resultid="3521" heatid="8891" lane="6" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1290" points="332" reactiontime="+75" swimtime="00:01:21.86" resultid="3522" heatid="9006" lane="1" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="344" reactiontime="+78" swimtime="00:01:28.97" resultid="3523" heatid="9042" lane="8" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="402" reactiontime="+71" swimtime="00:00:39.01" resultid="3524" heatid="9157" lane="3" entrytime="00:00:39.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700034" athleteid="3486">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="3487" heatid="8898" lane="8" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1239" points="165" reactiontime="+107" swimtime="00:03:39.66" resultid="3488" heatid="8973" lane="1" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.23" />
                    <SPLIT distance="100" swimtime="00:01:47.14" />
                    <SPLIT distance="150" swimtime="00:02:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="187" reactiontime="+103" swimtime="00:01:37.18" resultid="3489" heatid="9046" lane="7" entrytime="00:01:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="211" reactiontime="+108" swimtime="00:00:42.38" resultid="3490" heatid="9164" lane="0" entrytime="00:00:41.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1922-01-04" firstname="Kazimierz" gender="M" lastname="Mrówczyński" nation="POL" license="503105700021" athleteid="3515">
              <RESULTS>
                <RESULT eventid="1079" points="40" reactiontime="+120" swimtime="00:00:58.81" resultid="3516" heatid="8895" lane="6" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="32" reactiontime="+128" swimtime="00:02:20.30" resultid="3517" heatid="8986" lane="2" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="31" swimtime="00:05:13.41" resultid="3518" heatid="9095" lane="0" entrytime="00:04:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.35" />
                    <SPLIT distance="100" swimtime="00:02:31.91" />
                    <SPLIT distance="150" swimtime="00:03:54.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="39" reactiontime="+116" swimtime="00:01:13.88" resultid="3519" heatid="9160" lane="8" entrytime="00:01:12.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="3508">
              <RESULTS>
                <RESULT eventid="1079" points="242" swimtime="00:00:32.49" resultid="3509" heatid="8900" lane="5" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1113" points="126" reactiontime="+110" swimtime="00:03:38.43" resultid="3510" heatid="8923" lane="5" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                    <SPLIT distance="100" swimtime="00:01:54.18" />
                    <SPLIT distance="150" swimtime="00:02:57.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="203" reactiontime="+106" swimtime="00:01:16.44" resultid="3511" heatid="8988" lane="5" entrytime="00:01:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="142" reactiontime="+98" swimtime="00:01:37.09" resultid="3512" heatid="9010" lane="7" entrytime="00:01:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="179" reactiontime="+109" swimtime="00:00:38.67" resultid="3513" heatid="9063" lane="0" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="1613" points="97" reactiontime="+103" swimtime="00:01:45.24" resultid="3514" heatid="9130" lane="8" entrytime="00:01:47.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="3525">
              <RESULTS>
                <RESULT eventid="1062" points="373" reactiontime="+90" swimtime="00:00:32.28" resultid="3526" heatid="8890" lane="4" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1187" points="337" reactiontime="+75" swimtime="00:00:36.86" resultid="3527" heatid="8951" lane="4" entrytime="00:00:36.30" entrycourse="SCM" />
                <RESULT eventid="1256" points="296" reactiontime="+96" swimtime="00:01:16.50" resultid="3528" heatid="8982" lane="9" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="363" reactiontime="+95" swimtime="00:00:34.17" resultid="3529" heatid="9057" lane="3" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1457" points="269" reactiontime="+81" swimtime="00:01:25.20" resultid="3530" heatid="9076" lane="7" entrytime="00:01:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="266" reactiontime="+91" swimtime="00:01:24.82" resultid="3531" heatid="9126" lane="7" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-07-06" firstname="Alicja" gender="F" lastname="Michalak" nation="POL" license="503105600044" athleteid="3602">
              <RESULTS>
                <RESULT eventid="1222" points="353" reactiontime="+79" swimtime="00:03:10.40" resultid="3603" heatid="8970" lane="2" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                    <SPLIT distance="100" swimtime="00:01:29.46" />
                    <SPLIT distance="150" swimtime="00:02:18.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="360" reactiontime="+78" swimtime="00:01:19.65" resultid="3604" heatid="9006" lane="0" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="363" reactiontime="+74" swimtime="00:01:27.38" resultid="3605" heatid="9041" lane="7" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="338" reactiontime="+74" swimtime="00:02:38.95" resultid="3606" heatid="9092" lane="8" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="100" swimtime="00:01:17.78" />
                    <SPLIT distance="150" swimtime="00:01:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="409" reactiontime="+75" swimtime="00:00:38.77" resultid="3607" heatid="9157" lane="4" entrytime="00:00:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-20" firstname="Bogdan" gender="M" lastname="Wąsik" nation="POL" license="503105700025" athleteid="3560">
              <RESULTS>
                <RESULT eventid="1239" points="239" reactiontime="+100" swimtime="00:03:13.89" resultid="3561" heatid="8975" lane="0" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:31.88" />
                    <SPLIT distance="150" swimtime="00:02:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="137" reactiontime="+98" swimtime="00:03:30.46" resultid="3562" heatid="9027" lane="3" entrytime="00:03:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                    <SPLIT distance="100" swimtime="00:01:41.88" />
                    <SPLIT distance="150" swimtime="00:02:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="226" reactiontime="+99" swimtime="00:01:31.29" resultid="3563" heatid="9046" lane="3" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="168" reactiontime="+99" swimtime="00:07:06.76" resultid="3564" heatid="9116" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                    <SPLIT distance="100" swimtime="00:01:41.08" />
                    <SPLIT distance="150" swimtime="00:02:37.08" />
                    <SPLIT distance="200" swimtime="00:03:35.10" />
                    <SPLIT distance="250" swimtime="00:04:28.40" />
                    <SPLIT distance="300" swimtime="00:05:23.28" />
                    <SPLIT distance="350" swimtime="00:06:16.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="242" reactiontime="+96" swimtime="00:00:40.48" resultid="3565" heatid="9163" lane="5" entrytime="00:00:42.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-31" firstname="Mateusz" gender="M" lastname="Sass" nation="POL" license="503105700047" athleteid="3491">
              <RESULTS>
                <RESULT eventid="1079" points="479" reactiontime="+77" swimtime="00:00:25.89" resultid="3492" heatid="8914" lane="8" entrytime="00:00:25.90" entrycourse="SCM" />
                <RESULT eventid="1113" points="402" reactiontime="+84" swimtime="00:02:28.52" resultid="3493" heatid="8930" lane="2" entrytime="00:02:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="331" reactiontime="+65" swimtime="00:00:32.12" resultid="3494" heatid="8962" lane="9" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1307" points="462" reactiontime="+86" swimtime="00:01:05.52" resultid="3495" heatid="9020" lane="0" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="453" reactiontime="+78" swimtime="00:01:12.38" resultid="3496" heatid="9052" lane="4" entrytime="00:01:12.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="354" reactiontime="+87" swimtime="00:05:32.87" resultid="3497" heatid="9122" lane="0" entrytime="00:05:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:10.67" />
                    <SPLIT distance="200" swimtime="00:02:40.93" />
                    <SPLIT distance="250" swimtime="00:03:27.43" />
                    <SPLIT distance="300" swimtime="00:04:15.22" />
                    <SPLIT distance="350" swimtime="00:04:55.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="498" reactiontime="+81" swimtime="00:00:31.84" resultid="3498" heatid="9172" lane="1" entrytime="00:00:32.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="531" reactiontime="+74" swimtime="00:01:51.72" resultid="3628" heatid="9035" lane="8" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="100" swimtime="00:01:01.57" />
                    <SPLIT distance="150" swimtime="00:01:27.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3597" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="3491" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3592" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3612" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1548" points="564" reactiontime="+73" swimtime="00:01:39.93" resultid="3629" heatid="9112" lane="1" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.48" />
                    <SPLIT distance="100" swimtime="00:00:50.29" />
                    <SPLIT distance="150" swimtime="00:01:15.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3592" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3597" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="3491" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3612" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="252" reactiontime="+69" swimtime="00:02:23.26" resultid="3630" heatid="9033" lane="7" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:14.01" />
                    <SPLIT distance="150" swimtime="00:01:43.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3553" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3566" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3532" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3486" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="259" reactiontime="+70" swimtime="00:02:09.43" resultid="3631" heatid="9110" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:01:06.54" />
                    <SPLIT distance="150" swimtime="00:01:41.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3532" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="3486" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3566" number="3" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3553" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="3">
              <RESULTS>
                <RESULT comment="K15 - Brak dotknięcia ściany obydwoma rozłączonymi dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 13:31)" eventid="1381" reactiontime="+78" status="DSQ" swimtime="00:02:27.07" resultid="3632" heatid="9033" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:19.00" />
                    <SPLIT distance="150" swimtime="00:01:59.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3499" number="1" reactiontime="+78" status="DSQ" />
                    <RELAYPOSITION athleteid="3560" number="2" reactiontime="+80" status="DSQ" />
                    <RELAYPOSITION athleteid="3508" number="3" reactiontime="+67" status="DSQ" />
                    <RELAYPOSITION athleteid="3578" number="4" reactiontime="+71" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="225" reactiontime="+111" swimtime="00:02:15.69" resultid="3633" heatid="9110" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:00.39" />
                    <SPLIT distance="150" swimtime="00:01:26.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3508" number="1" reactiontime="+111" />
                    <RELAYPOSITION athleteid="3560" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3578" number="3" />
                    <RELAYPOSITION athleteid="3499" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1358" points="468" reactiontime="+68" swimtime="00:02:13.94" resultid="3626" heatid="9031" lane="5" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:12.68" />
                    <SPLIT distance="150" swimtime="00:01:45.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3546" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3539" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3520" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3571" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1525" points="463" reactiontime="+89" swimtime="00:02:01.74" resultid="3627" heatid="9108" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="100" swimtime="00:01:01.61" />
                    <SPLIT distance="150" swimtime="00:01:32.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3546" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3520" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="3539" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="3571" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="433" reactiontime="+79" swimtime="00:01:49.10" resultid="3623" heatid="8935" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.82" />
                    <SPLIT distance="100" swimtime="00:00:54.19" />
                    <SPLIT distance="150" swimtime="00:01:24.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3592" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="3546" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3539" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3612" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1698" points="436" reactiontime="+68" swimtime="00:01:59.31" resultid="3624" heatid="9176" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:04.16" />
                    <SPLIT distance="150" swimtime="00:01:31.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3546" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3491" number="2" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3592" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3571" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="221" reactiontime="+86" swimtime="00:02:16.58" resultid="3625" heatid="8934" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:09.76" />
                    <SPLIT distance="150" swimtime="00:01:44.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3525" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="3486" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3508" number="3" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3520" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1698" points="224" reactiontime="+72" swimtime="00:02:28.85" resultid="3634" heatid="9175" lane="8" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:19.32" />
                    <SPLIT distance="150" swimtime="00:01:55.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3525" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="3486" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="3520" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="3508" number="4" reactiontime="+91" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WAR" clubid="2878" name="Victory Masters Elbląg">
          <CONTACT name="Latecki Grzegorz" state="WAR" street="Łokietka 45" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1965-03-12" firstname="Grzegorz" gender="M" lastname="Latecki" nation="POL" athleteid="6149">
              <RESULTS>
                <RESULT eventid="1079" points="366" reactiontime="+78" swimtime="00:00:28.30" resultid="6150" heatid="8907" lane="6" entrytime="00:00:28.80" />
                <RESULT eventid="1205" points="259" reactiontime="+78" swimtime="00:00:34.83" resultid="6151" heatid="8960" lane="1" entrytime="00:00:34.50" />
                <RESULT eventid="1307" points="354" reactiontime="+80" swimtime="00:01:11.61" resultid="6152" heatid="9016" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="376" reactiontime="+86" swimtime="00:00:30.18" resultid="6153" heatid="9068" lane="2" entrytime="00:00:30.50" />
                <RESULT eventid="1578" points="289" reactiontime="+81" swimtime="00:05:56.00" resultid="6154" heatid="9120" lane="9" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:19.07" />
                    <SPLIT distance="150" swimtime="00:02:05.96" />
                    <SPLIT distance="200" swimtime="00:02:51.32" />
                    <SPLIT distance="250" swimtime="00:03:42.04" />
                    <SPLIT distance="300" swimtime="00:04:33.15" />
                    <SPLIT distance="350" swimtime="00:05:15.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="315" reactiontime="+85" swimtime="00:00:37.11" resultid="6155" heatid="9165" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1744" points="292" reactiontime="+82" swimtime="00:05:19.58" resultid="6156" heatid="9188" lane="9" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:54.19" />
                    <SPLIT distance="200" swimtime="00:02:35.61" />
                    <SPLIT distance="250" swimtime="00:03:17.50" />
                    <SPLIT distance="300" swimtime="00:03:59.38" />
                    <SPLIT distance="350" swimtime="00:04:41.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karas" nation="POL" athleteid="6143">
              <RESULTS>
                <RESULT eventid="1147" points="167" reactiontime="+108" swimtime="00:14:30.27" resultid="6144" heatid="8937" lane="0" entrytime="00:14:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.87" />
                    <SPLIT distance="100" swimtime="00:01:45.06" />
                    <SPLIT distance="150" swimtime="00:02:39.42" />
                    <SPLIT distance="200" swimtime="00:03:34.56" />
                    <SPLIT distance="250" swimtime="00:04:30.80" />
                    <SPLIT distance="300" swimtime="00:05:26.38" />
                    <SPLIT distance="350" swimtime="00:06:22.01" />
                    <SPLIT distance="400" swimtime="00:07:16.95" />
                    <SPLIT distance="450" swimtime="00:08:12.63" />
                    <SPLIT distance="500" swimtime="00:09:07.78" />
                    <SPLIT distance="550" swimtime="00:10:02.95" />
                    <SPLIT distance="600" swimtime="00:10:57.65" />
                    <SPLIT distance="650" swimtime="00:11:52.22" />
                    <SPLIT distance="700" swimtime="00:12:46.06" />
                    <SPLIT distance="750" swimtime="00:13:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="107" reactiontime="+112" swimtime="00:04:11.80" resultid="6145" heatid="9023" lane="6" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                    <SPLIT distance="100" swimtime="00:01:59.27" />
                    <SPLIT distance="150" swimtime="00:03:05.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="124" reactiontime="+107" swimtime="00:08:40.20" resultid="6146" heatid="9113" lane="6" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.57" />
                    <SPLIT distance="100" swimtime="00:01:57.71" />
                    <SPLIT distance="150" swimtime="00:03:10.69" />
                    <SPLIT distance="200" swimtime="00:04:18.29" />
                    <SPLIT distance="250" swimtime="00:05:35.42" />
                    <SPLIT distance="300" swimtime="00:06:54.15" />
                    <SPLIT distance="350" swimtime="00:07:48.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="98" reactiontime="+107" swimtime="00:01:58.39" resultid="6147" heatid="9124" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="164" reactiontime="+115" swimtime="00:07:08.16" resultid="6148" heatid="9178" lane="2" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.15" />
                    <SPLIT distance="100" swimtime="00:01:43.70" />
                    <SPLIT distance="150" swimtime="00:02:37.74" />
                    <SPLIT distance="200" swimtime="00:03:32.81" />
                    <SPLIT distance="250" swimtime="00:04:27.62" />
                    <SPLIT distance="300" swimtime="00:05:22.23" />
                    <SPLIT distance="350" swimtime="00:06:16.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-04" firstname="Karol" gender="M" lastname="Sosna" nation="POL" athleteid="6157">
              <RESULTS>
                <RESULT eventid="1079" points="284" reactiontime="+86" swimtime="00:00:30.82" resultid="6158" heatid="8904" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1406" points="303" reactiontime="+84" swimtime="00:01:22.71" resultid="6159" heatid="9049" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="351" reactiontime="+85" swimtime="00:00:35.79" resultid="6160" heatid="9168" lane="5" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-21" firstname="Tomasz" gender="M" lastname="Wysocki" nation="POL" athleteid="6129">
              <RESULTS>
                <RESULT eventid="1205" points="454" reactiontime="+76" swimtime="00:00:28.89" resultid="6130" heatid="8964" lane="7" entrytime="00:00:29.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner Mateusiak" nation="POL" athleteid="6161">
              <RESULTS>
                <RESULT eventid="1147" points="75" reactiontime="+131" swimtime="00:18:55.51" resultid="6162" heatid="8936" lane="2" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.23" />
                    <SPLIT distance="100" swimtime="00:02:06.90" />
                    <SPLIT distance="150" swimtime="00:03:18.96" />
                    <SPLIT distance="200" swimtime="00:04:31.93" />
                    <SPLIT distance="250" swimtime="00:05:44.18" />
                    <SPLIT distance="300" swimtime="00:06:56.61" />
                    <SPLIT distance="350" swimtime="00:08:08.31" />
                    <SPLIT distance="400" swimtime="00:09:19.97" />
                    <SPLIT distance="450" swimtime="00:10:31.66" />
                    <SPLIT distance="500" swimtime="00:11:43.99" />
                    <SPLIT distance="550" swimtime="00:12:55.92" />
                    <SPLIT distance="600" swimtime="00:14:08.05" />
                    <SPLIT distance="650" swimtime="00:15:20.25" />
                    <SPLIT distance="700" swimtime="00:16:32.37" />
                    <SPLIT distance="750" swimtime="00:17:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="57" reactiontime="+94" swimtime="00:01:06.59" resultid="6163" heatid="8948" lane="5" entrytime="00:01:20.00" />
                <RESULT comment="K13 - Stopy niezwrócone na zewnątrz w trakcie napędzającej części ruchu nóg (Time: 9:47), K-14" eventid="1222" reactiontime="+111" status="DSQ" swimtime="00:05:32.47" resultid="6164" heatid="8967" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.39" />
                    <SPLIT distance="100" swimtime="00:02:43.30" />
                    <SPLIT distance="150" swimtime="00:04:08.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="51" reactiontime="+122" swimtime="00:02:47.40" resultid="6165" heatid="9037" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="49" reactiontime="+86" swimtime="00:02:29.70" resultid="6166" heatid="9074" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="69" reactiontime="+117" swimtime="00:09:30.74" resultid="6167" heatid="9177" lane="4" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.31" />
                    <SPLIT distance="100" swimtime="00:02:11.30" />
                    <SPLIT distance="150" swimtime="00:03:26.01" />
                    <SPLIT distance="200" swimtime="00:04:39.63" />
                    <SPLIT distance="250" swimtime="00:05:53.40" />
                    <SPLIT distance="300" swimtime="00:07:07.21" />
                    <SPLIT distance="350" swimtime="00:08:21.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-06" firstname="Andrzej" gender="M" lastname="Pasieczny" nation="POL" athleteid="6131">
              <RESULTS>
                <RESULT eventid="1079" points="390" reactiontime="+92" swimtime="00:00:27.73" resultid="6132" heatid="8906" lane="7" entrytime="00:00:29.33" />
                <RESULT eventid="1341" points="410" reactiontime="+93" swimtime="00:02:26.13" resultid="6133" heatid="9030" lane="6" entrytime="00:02:23.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:06.65" />
                    <SPLIT distance="150" swimtime="00:01:43.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="457" reactiontime="+87" swimtime="00:02:09.00" resultid="6134" heatid="9105" lane="8" entrytime="00:02:08.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                    <SPLIT distance="100" swimtime="00:01:03.00" />
                    <SPLIT distance="150" swimtime="00:01:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="440" reactiontime="+91" swimtime="00:01:03.64" resultid="6135" heatid="9136" lane="9" entrytime="00:01:04.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1744" points="464" reactiontime="+99" swimtime="00:04:34.09" resultid="6136" heatid="9192" lane="0" entrytime="00:04:37.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:06.16" />
                    <SPLIT distance="150" swimtime="00:01:40.71" />
                    <SPLIT distance="200" swimtime="00:02:15.68" />
                    <SPLIT distance="250" swimtime="00:02:50.19" />
                    <SPLIT distance="300" swimtime="00:03:24.88" />
                    <SPLIT distance="350" swimtime="00:04:00.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="6137">
              <RESULTS>
                <RESULT eventid="1062" points="172" reactiontime="+107" swimtime="00:00:41.78" resultid="6138" heatid="8887" lane="1" entrytime="00:00:42.81" />
                <RESULT eventid="1147" reactiontime="+117" status="DNF" swimtime="00:00:00.00" resultid="6139" heatid="8937" lane="7" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.03" />
                    <SPLIT distance="100" swimtime="00:02:38.56" />
                    <SPLIT distance="150" swimtime="00:03:32.94" />
                    <SPLIT distance="200" swimtime="00:04:27.67" />
                    <SPLIT distance="250" swimtime="00:06:14.44" />
                    <SPLIT distance="300" swimtime="00:08:02.69" />
                    <SPLIT distance="350" swimtime="00:08:56.22" />
                    <SPLIT distance="400" swimtime="00:09:50.54" />
                    <SPLIT distance="450" swimtime="00:11:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="171" reactiontime="+110" swimtime="00:01:31.88" resultid="6140" heatid="8980" lane="0" entrytime="00:01:32.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="175" reactiontime="+102" swimtime="00:03:17.84" resultid="6141" heatid="9090" lane="9" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.53" />
                    <SPLIT distance="100" swimtime="00:01:39.44" />
                    <SPLIT distance="150" swimtime="00:02:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="177" reactiontime="+104" swimtime="00:06:57.35" resultid="6142" heatid="9178" lane="5" entrytime="00:06:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.56" />
                    <SPLIT distance="100" swimtime="00:01:43.11" />
                    <SPLIT distance="150" swimtime="00:02:36.32" />
                    <SPLIT distance="200" swimtime="00:03:28.96" />
                    <SPLIT distance="250" swimtime="00:04:22.16" />
                    <SPLIT distance="300" swimtime="00:05:15.09" />
                    <SPLIT distance="350" swimtime="00:06:07.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="406" reactiontime="+75" swimtime="00:02:02.15" resultid="6168" heatid="9034" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="100" swimtime="00:01:04.23" />
                    <SPLIT distance="150" swimtime="00:01:34.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6129" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="6157" number="2" reactiontime="+79" />
                    <RELAYPOSITION athleteid="6131" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="6149" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WMT" nation="POL" region="MAZ" clubid="3788" name="Warsaw Masters team">
          <CONTACT city="Warszawa" email="wojciech.kaluzynski@gmail.com" name="Kałużyński Wojciech" phone="607 45 4444" state="MAZ" />
          <ATHLETES>
            <ATHLETE birthdate="1975-10-20" firstname="Norbert" gender="M" lastname="Stablewski" nation="POL" athleteid="3955">
              <RESULTS>
                <RESULT eventid="1273" points="313" reactiontime="+92" swimtime="00:01:06.12" resultid="3956" heatid="8993" lane="0" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="301" reactiontime="+89" swimtime="00:02:28.24" resultid="3957" heatid="9099" lane="4" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:49.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-06-02" firstname="Wojciech" gender="M" lastname="Czupryn" nation="POL" athleteid="3988">
              <RESULTS>
                <RESULT eventid="1165" points="139" reactiontime="+105" swimtime="00:27:18.13" resultid="3989" heatid="8942" lane="1" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:36.52" />
                    <SPLIT distance="150" swimtime="00:02:30.14" />
                    <SPLIT distance="200" swimtime="00:03:24.27" />
                    <SPLIT distance="250" swimtime="00:04:18.21" />
                    <SPLIT distance="300" swimtime="00:05:12.93" />
                    <SPLIT distance="350" swimtime="00:06:07.13" />
                    <SPLIT distance="400" swimtime="00:07:00.12" />
                    <SPLIT distance="450" swimtime="00:07:53.62" />
                    <SPLIT distance="500" swimtime="00:08:47.16" />
                    <SPLIT distance="550" swimtime="00:09:40.07" />
                    <SPLIT distance="600" swimtime="00:10:34.54" />
                    <SPLIT distance="650" swimtime="00:11:30.14" />
                    <SPLIT distance="700" swimtime="00:12:26.22" />
                    <SPLIT distance="750" swimtime="00:13:21.93" />
                    <SPLIT distance="800" swimtime="00:14:17.84" />
                    <SPLIT distance="850" swimtime="00:15:13.47" />
                    <SPLIT distance="900" swimtime="00:16:08.46" />
                    <SPLIT distance="950" swimtime="00:17:04.27" />
                    <SPLIT distance="1000" swimtime="00:18:00.44" />
                    <SPLIT distance="1050" swimtime="00:18:55.76" />
                    <SPLIT distance="1100" swimtime="00:19:51.67" />
                    <SPLIT distance="1150" swimtime="00:20:46.86" />
                    <SPLIT distance="1200" swimtime="00:21:42.71" />
                    <SPLIT distance="1250" swimtime="00:22:38.31" />
                    <SPLIT distance="1300" swimtime="00:23:33.91" />
                    <SPLIT distance="1350" swimtime="00:24:29.90" />
                    <SPLIT distance="1400" swimtime="00:25:26.77" />
                    <SPLIT distance="1450" swimtime="00:26:23.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="95" reactiontime="+90" swimtime="00:00:48.61" resultid="3990" heatid="8956" lane="6" entrytime="00:00:48.00" />
                <RESULT eventid="1307" points="125" reactiontime="+85" swimtime="00:01:41.30" resultid="3991" heatid="9010" lane="9" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="124" reactiontime="+92" swimtime="00:01:51.23" resultid="3992" heatid="9045" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="98" reactiontime="+93" swimtime="00:01:45.85" resultid="3993" heatid="9080" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="93" reactiontime="+87" swimtime="00:03:53.99" resultid="3994" heatid="9145" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.29" />
                    <SPLIT distance="100" swimtime="00:01:52.44" />
                    <SPLIT distance="150" swimtime="00:02:53.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="131" reactiontime="+101" swimtime="00:06:57.19" resultid="3995" heatid="9184" lane="7" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="100" swimtime="00:01:32.48" />
                    <SPLIT distance="150" swimtime="00:02:22.57" />
                    <SPLIT distance="200" swimtime="00:03:14.54" />
                    <SPLIT distance="300" swimtime="00:05:07.91" />
                    <SPLIT distance="350" swimtime="00:06:03.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-28" firstname="Paweł" gender="M" lastname="Rogosz" nation="POL" athleteid="3909">
              <RESULTS>
                <RESULT eventid="1113" points="374" reactiontime="+96" swimtime="00:02:32.07" resultid="3910" heatid="8928" lane="5" entrytime="00:02:38.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="150" swimtime="00:01:56.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="333" reactiontime="+100" swimtime="00:20:26.41" resultid="3911" heatid="8945" lane="6" entrytime="00:21:15.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:14.05" />
                    <SPLIT distance="150" swimtime="00:01:53.29" />
                    <SPLIT distance="200" swimtime="00:02:33.68" />
                    <SPLIT distance="250" swimtime="00:03:13.64" />
                    <SPLIT distance="300" swimtime="00:03:53.80" />
                    <SPLIT distance="350" swimtime="00:04:33.90" />
                    <SPLIT distance="400" swimtime="00:05:13.61" />
                    <SPLIT distance="450" swimtime="00:05:53.99" />
                    <SPLIT distance="500" swimtime="00:06:34.47" />
                    <SPLIT distance="550" swimtime="00:07:15.70" />
                    <SPLIT distance="600" swimtime="00:07:56.67" />
                    <SPLIT distance="650" swimtime="00:08:37.96" />
                    <SPLIT distance="700" swimtime="00:09:19.19" />
                    <SPLIT distance="750" swimtime="00:10:00.18" />
                    <SPLIT distance="800" swimtime="00:10:41.23" />
                    <SPLIT distance="850" swimtime="00:11:22.12" />
                    <SPLIT distance="900" swimtime="00:12:04.36" />
                    <SPLIT distance="950" swimtime="00:12:45.69" />
                    <SPLIT distance="1000" swimtime="00:13:27.32" />
                    <SPLIT distance="1050" swimtime="00:14:08.77" />
                    <SPLIT distance="1100" swimtime="00:14:50.62" />
                    <SPLIT distance="1150" swimtime="00:15:33.41" />
                    <SPLIT distance="1200" swimtime="00:16:16.31" />
                    <SPLIT distance="1250" swimtime="00:16:58.60" />
                    <SPLIT distance="1300" swimtime="00:17:41.33" />
                    <SPLIT distance="1350" swimtime="00:18:23.81" />
                    <SPLIT distance="1400" swimtime="00:19:05.39" />
                    <SPLIT distance="1450" swimtime="00:19:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="361" reactiontime="+97" swimtime="00:02:49.18" resultid="3912" heatid="8977" lane="8" entrytime="00:02:55.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:05.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="329" reactiontime="+103" swimtime="00:02:37.15" resultid="3913" heatid="9029" lane="8" entrytime="00:02:48.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:15.81" />
                    <SPLIT distance="150" swimtime="00:01:56.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-17" firstname="Waldemar" gender="M" lastname="de Makay" nation="POL" athleteid="3814">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 16:35)" eventid="1079" reactiontime="+55" status="DSQ" swimtime="00:00:32.49" resultid="3815" heatid="8901" lane="8" entrytime="00:00:32.00" />
                <RESULT comment="Rekord Polski" eventid="1165" points="233" reactiontime="+121" swimtime="00:23:01.16" resultid="3816" heatid="8944" lane="0" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:01:25.64" />
                    <SPLIT distance="150" swimtime="00:02:10.70" />
                    <SPLIT distance="200" swimtime="00:02:55.56" />
                    <SPLIT distance="250" swimtime="00:03:40.73" />
                    <SPLIT distance="300" swimtime="00:04:26.02" />
                    <SPLIT distance="350" swimtime="00:05:12.15" />
                    <SPLIT distance="400" swimtime="00:05:58.44" />
                    <SPLIT distance="450" swimtime="00:06:45.14" />
                    <SPLIT distance="500" swimtime="00:07:31.50" />
                    <SPLIT distance="550" swimtime="00:08:17.68" />
                    <SPLIT distance="600" swimtime="00:09:04.20" />
                    <SPLIT distance="650" swimtime="00:09:50.46" />
                    <SPLIT distance="700" swimtime="00:10:37.30" />
                    <SPLIT distance="750" swimtime="00:11:23.61" />
                    <SPLIT distance="800" swimtime="00:12:10.11" />
                    <SPLIT distance="850" swimtime="00:12:56.55" />
                    <SPLIT distance="900" swimtime="00:13:42.72" />
                    <SPLIT distance="950" swimtime="00:14:29.11" />
                    <SPLIT distance="1000" swimtime="00:15:15.27" />
                    <SPLIT distance="1050" swimtime="00:16:01.73" />
                    <SPLIT distance="1100" swimtime="00:16:48.02" />
                    <SPLIT distance="1150" swimtime="00:17:34.20" />
                    <SPLIT distance="1200" swimtime="00:18:20.29" />
                    <SPLIT distance="1250" swimtime="00:19:07.09" />
                    <SPLIT distance="1300" swimtime="00:19:53.90" />
                    <SPLIT distance="1350" swimtime="00:20:40.51" />
                    <SPLIT distance="1400" swimtime="00:21:27.86" />
                    <SPLIT distance="1450" swimtime="00:22:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="139" reactiontime="+78" swimtime="00:00:42.85" resultid="3817" heatid="8958" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1273" points="220" reactiontime="+110" swimtime="00:01:14.34" resultid="3818" heatid="8990" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="149" reactiontime="+74" swimtime="00:01:32.16" resultid="3819" heatid="9082" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="217" reactiontime="+115" swimtime="00:02:45.15" resultid="3820" heatid="9099" lane="7" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="150" swimtime="00:02:01.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="151" reactiontime="+84" swimtime="00:03:19.01" resultid="3821" heatid="9146" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                    <SPLIT distance="100" swimtime="00:01:36.17" />
                    <SPLIT distance="150" swimtime="00:02:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="225" reactiontime="+114" swimtime="00:05:48.49" resultid="3822" heatid="9187" lane="9" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:01:21.56" />
                    <SPLIT distance="150" swimtime="00:02:05.42" />
                    <SPLIT distance="200" swimtime="00:02:49.63" />
                    <SPLIT distance="250" swimtime="00:03:34.22" />
                    <SPLIT distance="300" swimtime="00:04:19.63" />
                    <SPLIT distance="350" swimtime="00:05:04.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-31" firstname="Katharina" gender="F" lastname="Szymańska" nation="POL" athleteid="4014">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="4015" heatid="8887" lane="4" entrytime="00:00:39.99" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="4016" heatid="8950" lane="8" entrytime="00:00:45.99" />
                <RESULT eventid="1290" points="164" reactiontime="+79" swimtime="00:01:43.44" resultid="4017" heatid="9002" lane="2" entrytime="00:01:45.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="120" reactiontime="+82" swimtime="00:00:49.32" resultid="4018" heatid="9055" lane="3" entrytime="00:00:46.99" />
                <RESULT eventid="1664" points="194" reactiontime="+90" swimtime="00:00:49.70" resultid="4019" heatid="9154" lane="8" entrytime="00:00:48.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-10" firstname="Tomasz" gender="M" lastname="Porada" nation="POL" athleteid="3855">
              <RESULTS>
                <RESULT eventid="1113" points="394" reactiontime="+79" swimtime="00:02:29.43" resultid="3856" heatid="8929" lane="6" entrytime="00:02:31.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:53.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="397" reactiontime="+90" swimtime="00:19:16.63" resultid="3857" heatid="8947" lane="7" entrytime="00:19:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:12.12" />
                    <SPLIT distance="150" swimtime="00:01:50.25" />
                    <SPLIT distance="200" swimtime="00:02:29.08" />
                    <SPLIT distance="250" swimtime="00:03:07.62" />
                    <SPLIT distance="300" swimtime="00:03:46.69" />
                    <SPLIT distance="350" swimtime="00:04:25.77" />
                    <SPLIT distance="400" swimtime="00:05:04.75" />
                    <SPLIT distance="450" swimtime="00:05:43.31" />
                    <SPLIT distance="550" swimtime="00:07:00.90" />
                    <SPLIT distance="600" swimtime="00:07:39.58" />
                    <SPLIT distance="650" swimtime="00:08:17.92" />
                    <SPLIT distance="700" swimtime="00:08:56.01" />
                    <SPLIT distance="750" swimtime="00:09:34.53" />
                    <SPLIT distance="800" swimtime="00:10:13.02" />
                    <SPLIT distance="850" swimtime="00:10:51.26" />
                    <SPLIT distance="900" swimtime="00:11:29.98" />
                    <SPLIT distance="950" swimtime="00:12:08.31" />
                    <SPLIT distance="1000" swimtime="00:12:47.60" />
                    <SPLIT distance="1050" swimtime="00:13:25.81" />
                    <SPLIT distance="1100" swimtime="00:14:04.60" />
                    <SPLIT distance="1150" swimtime="00:14:43.60" />
                    <SPLIT distance="1200" swimtime="00:15:22.82" />
                    <SPLIT distance="1250" swimtime="00:16:02.19" />
                    <SPLIT distance="1300" swimtime="00:17:20.46" />
                    <SPLIT distance="1350" swimtime="00:17:59.87" />
                    <SPLIT distance="1400" swimtime="00:18:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="431" reactiontime="+87" swimtime="00:02:39.42" resultid="3858" heatid="8978" lane="1" entrytime="00:02:38.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:01:57.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3859" heatid="8997" lane="7" entrytime="00:01:00.44" />
                <RESULT eventid="1406" points="427" reactiontime="+74" swimtime="00:01:13.81" resultid="3860" heatid="9053" lane="9" entrytime="00:01:12.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="413" reactiontime="+79" swimtime="00:05:16.04" resultid="3861" heatid="9122" lane="8" entrytime="00:05:18.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="150" swimtime="00:01:56.18" />
                    <SPLIT distance="200" swimtime="00:02:39.51" />
                    <SPLIT distance="250" swimtime="00:03:21.09" />
                    <SPLIT distance="300" swimtime="00:04:03.70" />
                    <SPLIT distance="350" swimtime="00:04:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="432" reactiontime="+72" swimtime="00:00:33.38" resultid="3862" heatid="9171" lane="2" entrytime="00:00:33.70" />
                <RESULT eventid="1744" points="415" reactiontime="+85" swimtime="00:04:44.44" resultid="3863" heatid="9191" lane="8" entrytime="00:04:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:43.72" />
                    <SPLIT distance="200" swimtime="00:02:56.86" />
                    <SPLIT distance="250" swimtime="00:03:32.92" />
                    <SPLIT distance="300" swimtime="00:04:09.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-05" firstname="Bartłomiej" gender="M" lastname="Pawłowski" nation="POL" athleteid="3934">
              <RESULTS>
                <RESULT eventid="1079" points="389" reactiontime="+81" swimtime="00:00:27.74" resultid="3935" heatid="8906" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1273" points="339" reactiontime="+86" swimtime="00:01:04.45" resultid="3936" heatid="8994" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="339" reactiontime="+85" swimtime="00:01:19.70" resultid="3937" heatid="9049" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="399" reactiontime="+82" swimtime="00:00:34.28" resultid="3938" heatid="9168" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-18" firstname="Jacek" gender="M" lastname="Czupryn" nation="POL" athleteid="3996" />
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="3949">
              <RESULTS>
                <RESULT eventid="1239" points="201" reactiontime="+110" swimtime="00:03:25.36" resultid="3950" heatid="8974" lane="1" entrytime="00:03:21.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="100" swimtime="00:01:36.12" />
                    <SPLIT distance="150" swimtime="00:02:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="106" reactiontime="+108" swimtime="00:03:48.73" resultid="3951" heatid="9026" lane="3" entrytime="00:04:09.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="100" swimtime="00:01:45.54" />
                    <SPLIT distance="150" swimtime="00:02:46.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="202" reactiontime="+101" swimtime="00:01:34.63" resultid="3952" heatid="9046" lane="5" entrytime="00:01:31.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="122" reactiontime="+105" swimtime="00:01:37.48" resultid="3953" heatid="9130" lane="4" entrytime="00:01:35.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="209" reactiontime="+100" swimtime="00:00:42.52" resultid="3954" heatid="9163" lane="6" entrytime="00:00:42.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-22" firstname="Daniel" gender="M" lastname="Żółtowski" nation="POL" athleteid="3901">
              <RESULTS>
                <RESULT eventid="1079" points="368" reactiontime="+78" swimtime="00:00:28.27" resultid="3902" heatid="8908" lane="0" entrytime="00:00:28.20" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="3903" heatid="8945" lane="9" entrytime="00:21:55.00" />
                <RESULT eventid="1205" points="279" reactiontime="+69" swimtime="00:00:34.00" resultid="3904" heatid="8961" lane="8" entrytime="00:00:33.20" />
                <RESULT eventid="1273" points="375" reactiontime="+84" swimtime="00:01:02.30" resultid="3905" heatid="8997" lane="8" entrytime="00:01:00.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="334" reactiontime="+83" swimtime="00:00:31.41" resultid="3906" heatid="9067" lane="2" entrytime="00:00:31.40" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="3907" heatid="9102" lane="2" entrytime="00:02:18.90" />
                <RESULT eventid="1744" points="335" reactiontime="+86" swimtime="00:05:05.33" resultid="3908" heatid="9188" lane="4" entrytime="00:05:10.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:09.06" />
                    <SPLIT distance="150" swimtime="00:01:46.82" />
                    <SPLIT distance="200" swimtime="00:02:25.27" />
                    <SPLIT distance="250" swimtime="00:03:04.57" />
                    <SPLIT distance="300" swimtime="00:03:44.68" />
                    <SPLIT distance="350" swimtime="00:04:24.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="3832">
              <RESULTS>
                <RESULT eventid="1113" points="420" reactiontime="+85" swimtime="00:02:26.38" resultid="3833" heatid="8929" lane="1" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                    <SPLIT distance="150" swimtime="00:01:52.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="385" reactiontime="+85" swimtime="00:00:30.52" resultid="3834" heatid="8962" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1307" points="450" reactiontime="+82" swimtime="00:01:06.07" resultid="3835" heatid="9019" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="417" reactiontime="+71" swimtime="00:01:05.47" resultid="3836" heatid="9085" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="436" reactiontime="+84" swimtime="00:02:11.00" resultid="3837" heatid="9103" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:04.84" />
                    <SPLIT distance="150" swimtime="00:01:38.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="392" reactiontime="+76" swimtime="00:02:24.96" resultid="3838" heatid="9149" lane="0" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:09.00" />
                    <SPLIT distance="150" swimtime="00:01:46.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="4020">
              <RESULTS>
                <RESULT eventid="1290" points="270" reactiontime="+93" swimtime="00:01:27.65" resultid="4021" heatid="9004" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="253" reactiontime="+86" swimtime="00:00:38.53" resultid="4022" heatid="9056" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1491" points="286" reactiontime="+90" swimtime="00:02:48.00" resultid="4023" heatid="9091" lane="1" entrytime="00:02:53.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="150" swimtime="00:02:06.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="211" reactiontime="+88" swimtime="00:01:31.70" resultid="4024" heatid="9125" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-14" firstname="Wojciech" gender="M" lastname="Kałużyński" nation="POL" athleteid="3939">
              <RESULTS>
                <RESULT eventid="1079" points="293" reactiontime="+86" swimtime="00:00:30.50" resultid="3940" heatid="8904" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1113" points="252" reactiontime="+94" swimtime="00:02:53.44" resultid="3941" heatid="8925" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:22.57" />
                    <SPLIT distance="150" swimtime="00:02:12.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="288" reactiontime="+88" swimtime="00:01:16.69" resultid="3942" heatid="9014" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="262" reactiontime="+85" swimtime="00:00:34.04" resultid="3943" heatid="9064" lane="8" entrytime="00:00:35.57" />
                <RESULT eventid="1508" points="281" reactiontime="+86" swimtime="00:02:31.68" resultid="3944" heatid="9100" lane="9" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:13.43" />
                    <SPLIT distance="150" swimtime="00:01:52.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="268" reactiontime="+90" swimtime="00:05:29.16" resultid="3945" heatid="9187" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.75" />
                    <SPLIT distance="100" swimtime="00:01:57.99" />
                    <SPLIT distance="150" swimtime="00:02:39.49" />
                    <SPLIT distance="250" swimtime="00:03:21.71" />
                    <SPLIT distance="300" swimtime="00:04:04.99" />
                    <SPLIT distance="350" swimtime="00:04:47.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-02-17" firstname="Piotr" gender="M" lastname="Barski" nation="POL" athleteid="3883">
              <RESULTS>
                <RESULT eventid="1079" points="435" reactiontime="+80" swimtime="00:00:26.73" resultid="3884" heatid="8909" lane="6" entrytime="00:00:27.90" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="3885" heatid="8972" lane="5" entrytime="00:03:50.00" />
                <RESULT eventid="1273" points="447" reactiontime="+77" swimtime="00:00:58.76" resultid="3886" heatid="8998" lane="9" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="407" reactiontime="+72" swimtime="00:01:15.02" resultid="3887" heatid="9048" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="405" reactiontime="+79" swimtime="00:00:29.46" resultid="3888" heatid="9070" lane="3" entrytime="00:00:28.50" />
                <RESULT comment="Rekord Polski" eventid="1681" points="420" reactiontime="+87" swimtime="00:00:33.69" resultid="3889" heatid="9170" lane="0" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-09" firstname="Tomasz" gender="M" lastname="Makomaski" nation="POL" athleteid="3890">
              <RESULTS>
                <RESULT eventid="1273" points="382" reactiontime="+76" swimtime="00:01:01.91" resultid="3891" heatid="8995" lane="8" entrytime="00:01:02.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="376" reactiontime="+74" swimtime="00:01:16.98" resultid="3892" heatid="9052" lane="9" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="389" reactiontime="+76" swimtime="00:00:34.56" resultid="3893" heatid="9170" lane="6" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="Barbara" gender="F" lastname="Łowkis" nation="POL" athleteid="3928">
              <RESULTS>
                <RESULT eventid="1062" points="172" reactiontime="+99" swimtime="00:00:41.72" resultid="3929" heatid="8887" lane="9" entrytime="00:00:43.59" />
                <RESULT eventid="1187" points="146" reactiontime="+93" swimtime="00:00:48.65" resultid="3930" heatid="8949" lane="2" entrytime="00:00:50.70" />
                <RESULT eventid="1256" points="121" reactiontime="+114" swimtime="00:01:43.01" resultid="3931" heatid="8979" lane="6" entrytime="00:01:42.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="89" reactiontime="+110" swimtime="00:00:54.51" resultid="3932" heatid="9054" lane="1" />
                <RESULT eventid="1457" points="121" reactiontime="+90" swimtime="00:01:51.10" resultid="3933" heatid="9075" lane="2" entrytime="00:01:53.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="4003">
              <RESULTS>
                <RESULT eventid="1062" points="110" reactiontime="+103" swimtime="00:00:48.44" resultid="4004" heatid="8886" lane="6" entrytime="00:00:49.43" />
                <RESULT eventid="1147" points="119" reactiontime="+108" swimtime="00:16:12.70" resultid="4005" heatid="8936" lane="5" entrytime="00:16:55.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.55" />
                    <SPLIT distance="100" swimtime="00:01:54.47" />
                    <SPLIT distance="150" swimtime="00:02:57.82" />
                    <SPLIT distance="200" swimtime="00:03:59.73" />
                    <SPLIT distance="250" swimtime="00:05:03.27" />
                    <SPLIT distance="300" swimtime="00:06:06.69" />
                    <SPLIT distance="350" swimtime="00:07:07.72" />
                    <SPLIT distance="400" swimtime="00:08:08.69" />
                    <SPLIT distance="450" swimtime="00:09:10.46" />
                    <SPLIT distance="500" swimtime="00:10:11.73" />
                    <SPLIT distance="550" swimtime="00:11:12.19" />
                    <SPLIT distance="600" swimtime="00:12:13.48" />
                    <SPLIT distance="650" swimtime="00:13:14.32" />
                    <SPLIT distance="700" swimtime="00:14:14.56" />
                    <SPLIT distance="750" swimtime="00:15:14.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="98" reactiontime="+94" swimtime="00:03:59.70" resultid="4006" heatid="9089" lane="8" entrytime="00:04:04.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.42" />
                    <SPLIT distance="100" swimtime="00:01:54.46" />
                    <SPLIT distance="150" swimtime="00:02:57.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="98" reactiontime="+106" swimtime="00:08:27.74" resultid="4007" heatid="9178" lane="0" entrytime="00:08:07.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.76" />
                    <SPLIT distance="150" swimtime="00:03:05.17" />
                    <SPLIT distance="200" swimtime="00:04:10.89" />
                    <SPLIT distance="250" swimtime="00:05:15.56" />
                    <SPLIT distance="300" swimtime="00:06:22.38" />
                    <SPLIT distance="350" swimtime="00:07:26.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="3975">
              <RESULTS>
                <RESULT eventid="1079" points="402" reactiontime="+78" swimtime="00:00:27.43" resultid="3976" heatid="8909" lane="4" entrytime="00:00:27.80" />
                <RESULT eventid="1165" points="353" reactiontime="+85" swimtime="00:20:02.55" resultid="3977" heatid="8944" lane="6" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:12.76" />
                    <SPLIT distance="150" swimtime="00:01:51.28" />
                    <SPLIT distance="200" swimtime="00:02:30.63" />
                    <SPLIT distance="250" swimtime="00:03:09.66" />
                    <SPLIT distance="300" swimtime="00:03:49.18" />
                    <SPLIT distance="350" swimtime="00:04:29.18" />
                    <SPLIT distance="400" swimtime="00:05:09.41" />
                    <SPLIT distance="450" swimtime="00:05:49.65" />
                    <SPLIT distance="500" swimtime="00:06:30.07" />
                    <SPLIT distance="550" swimtime="00:07:10.56" />
                    <SPLIT distance="600" swimtime="00:07:50.83" />
                    <SPLIT distance="650" swimtime="00:08:31.60" />
                    <SPLIT distance="700" swimtime="00:09:11.97" />
                    <SPLIT distance="750" swimtime="00:09:52.40" />
                    <SPLIT distance="800" swimtime="00:10:33.61" />
                    <SPLIT distance="850" swimtime="00:11:14.19" />
                    <SPLIT distance="900" swimtime="00:11:54.88" />
                    <SPLIT distance="950" swimtime="00:12:35.47" />
                    <SPLIT distance="1000" swimtime="00:13:16.12" />
                    <SPLIT distance="1050" swimtime="00:13:57.23" />
                    <SPLIT distance="1100" swimtime="00:14:38.34" />
                    <SPLIT distance="1150" swimtime="00:15:19.71" />
                    <SPLIT distance="1200" swimtime="00:16:01.40" />
                    <SPLIT distance="1250" swimtime="00:16:43.06" />
                    <SPLIT distance="1300" swimtime="00:17:24.62" />
                    <SPLIT distance="1350" swimtime="00:18:05.74" />
                    <SPLIT distance="1400" swimtime="00:18:45.62" />
                    <SPLIT distance="1450" swimtime="00:19:21.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="381" reactiontime="+80" swimtime="00:01:01.94" resultid="3978" heatid="8995" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="354" reactiontime="+81" swimtime="00:00:30.79" resultid="3979" heatid="9068" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1508" points="376" reactiontime="+87" swimtime="00:02:17.58" resultid="3980" heatid="9102" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="100" swimtime="00:01:07.19" />
                    <SPLIT distance="150" swimtime="00:01:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="351" reactiontime="+77" swimtime="00:05:00.81" resultid="3981" heatid="9189" lane="8" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:11.11" />
                    <SPLIT distance="150" swimtime="00:01:48.98" />
                    <SPLIT distance="200" swimtime="00:02:27.41" />
                    <SPLIT distance="250" swimtime="00:03:06.68" />
                    <SPLIT distance="300" swimtime="00:03:45.53" />
                    <SPLIT distance="350" swimtime="00:04:24.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-28" firstname="Krzysztof" gender="M" lastname="Olszewski" nation="POL" athleteid="3848">
              <RESULTS>
                <RESULT eventid="1113" points="371" reactiontime="+71" swimtime="00:02:32.47" resultid="3849" heatid="8929" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:11.37" />
                    <SPLIT distance="150" swimtime="00:01:54.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="381" reactiontime="+81" swimtime="00:02:46.09" resultid="3850" heatid="8977" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="150" swimtime="00:02:01.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="442" reactiontime="+82" swimtime="00:01:06.48" resultid="3851" heatid="9019" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="418" reactiontime="+79" swimtime="00:01:14.36" resultid="3852" heatid="9052" lane="2" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="369" reactiontime="+80" swimtime="00:01:08.18" resultid="3853" heatid="9085" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="452" reactiontime="+73" swimtime="00:00:32.90" resultid="3854" heatid="9171" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="3969">
              <RESULTS>
                <RESULT eventid="1222" points="363" reactiontime="+85" swimtime="00:03:08.59" resultid="3970" heatid="8970" lane="6" entrytime="00:03:11.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                    <SPLIT distance="100" swimtime="00:01:31.60" />
                    <SPLIT distance="150" swimtime="00:02:19.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="366" reactiontime="+86" swimtime="00:01:27.16" resultid="3971" heatid="9042" lane="0" entrytime="00:01:28.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="298" reactiontime="+83" swimtime="00:02:45.81" resultid="3972" heatid="9091" lane="2" entrytime="00:02:50.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:22.45" />
                    <SPLIT distance="150" swimtime="00:02:04.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="350" reactiontime="+83" swimtime="00:00:40.84" resultid="3973" heatid="9157" lane="1" entrytime="00:00:40.28" />
                <RESULT eventid="1721" points="300" reactiontime="+83" swimtime="00:05:50.10" resultid="3974" heatid="9180" lane="6" entrytime="00:05:49.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:25.43" />
                    <SPLIT distance="150" swimtime="00:02:10.69" />
                    <SPLIT distance="200" swimtime="00:02:55.58" />
                    <SPLIT distance="250" swimtime="00:03:38.40" />
                    <SPLIT distance="300" swimtime="00:04:22.58" />
                    <SPLIT distance="350" swimtime="00:05:07.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-07" firstname="Paulina" gender="F" lastname="Mroczek" nation="POL" athleteid="3946">
              <RESULTS>
                <RESULT eventid="1256" points="346" reactiontime="+84" swimtime="00:01:12.62" resultid="3947" heatid="8983" lane="9" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="305" reactiontime="+87" swimtime="00:02:44.45" resultid="3948" heatid="9092" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:16.98" />
                    <SPLIT distance="150" swimtime="00:02:00.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="F" lastname="Nawrocka" nation="POL" athleteid="3809">
              <RESULTS>
                <RESULT eventid="1290" points="465" reactiontime="+87" swimtime="00:01:13.15" resultid="3810" heatid="9007" lane="1" entrytime="00:01:13.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="399" reactiontime="+87" swimtime="00:01:24.68" resultid="3811" heatid="9042" lane="6" entrytime="00:01:23.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="3812" heatid="9126" lane="3" entrytime="00:01:19.80" />
                <RESULT eventid="1664" points="388" reactiontime="+81" swimtime="00:00:39.48" resultid="3813" heatid="9158" lane="9" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" athleteid="3982">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1062" points="620" reactiontime="+73" swimtime="00:00:27.25" resultid="3983" heatid="8885" lane="3" />
                <RESULT comment="Rekord Polski" eventid="1096" points="559" reactiontime="+78" swimtime="00:02:27.85" resultid="3984" heatid="8916" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                    <SPLIT distance="100" swimtime="00:01:10.31" />
                    <SPLIT distance="150" swimtime="00:01:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1324" points="491" reactiontime="+69" swimtime="00:02:31.53" resultid="3985" heatid="9022" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:09.30" />
                    <SPLIT distance="150" swimtime="00:01:48.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="564" reactiontime="+74" swimtime="00:00:29.50" resultid="3986" heatid="9059" lane="5" entrytime="00:00:29.80" />
                <RESULT eventid="1595" points="591" reactiontime="+74" swimtime="00:01:05.05" resultid="3987" heatid="9127" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-10" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="4008">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="4009" heatid="8914" lane="4" entrytime="00:00:24.50" />
                <RESULT eventid="1307" points="504" reactiontime="+78" swimtime="00:01:03.65" resultid="4010" heatid="9021" lane="8" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="482" reactiontime="+74" swimtime="00:00:27.79" resultid="4011" heatid="9072" lane="8" entrytime="00:00:27.50" />
                <RESULT eventid="1578" points="386" reactiontime="+84" swimtime="00:05:23.40" resultid="4012" heatid="9122" lane="9" entrytime="00:05:20.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                    <SPLIT distance="150" swimtime="00:01:52.38" />
                    <SPLIT distance="200" swimtime="00:02:33.90" />
                    <SPLIT distance="250" swimtime="00:03:19.46" />
                    <SPLIT distance="300" swimtime="00:04:05.49" />
                    <SPLIT distance="350" swimtime="00:04:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="459" reactiontime="+86" swimtime="00:00:32.71" resultid="4013" heatid="9171" lane="1" entrytime="00:00:33.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="3839">
              <RESULTS>
                <RESULT eventid="1079" points="152" reactiontime="+101" swimtime="00:00:37.89" resultid="3840" heatid="8898" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1165" points="105" reactiontime="+102" swimtime="00:29:58.06" resultid="3841" heatid="8941" lane="3" entrytime="00:32:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.17" />
                    <SPLIT distance="100" swimtime="00:01:47.25" />
                    <SPLIT distance="150" swimtime="00:02:45.67" />
                    <SPLIT distance="200" swimtime="00:03:46.08" />
                    <SPLIT distance="250" swimtime="00:04:46.08" />
                    <SPLIT distance="300" swimtime="00:05:45.74" />
                    <SPLIT distance="350" swimtime="00:06:46.51" />
                    <SPLIT distance="400" swimtime="00:07:48.42" />
                    <SPLIT distance="450" swimtime="00:08:48.40" />
                    <SPLIT distance="500" swimtime="00:09:49.21" />
                    <SPLIT distance="550" swimtime="00:10:49.62" />
                    <SPLIT distance="600" swimtime="00:11:51.66" />
                    <SPLIT distance="650" swimtime="00:12:52.07" />
                    <SPLIT distance="700" swimtime="00:13:53.04" />
                    <SPLIT distance="750" swimtime="00:14:53.94" />
                    <SPLIT distance="800" swimtime="00:15:54.00" />
                    <SPLIT distance="850" swimtime="00:16:54.34" />
                    <SPLIT distance="900" swimtime="00:17:55.22" />
                    <SPLIT distance="950" swimtime="00:18:54.71" />
                    <SPLIT distance="1000" swimtime="00:19:55.86" />
                    <SPLIT distance="1050" swimtime="00:20:57.39" />
                    <SPLIT distance="1100" swimtime="00:21:57.99" />
                    <SPLIT distance="1150" swimtime="00:22:59.72" />
                    <SPLIT distance="1200" swimtime="00:23:59.59" />
                    <SPLIT distance="1250" swimtime="00:24:59.95" />
                    <SPLIT distance="1300" swimtime="00:26:00.14" />
                    <SPLIT distance="1350" swimtime="00:27:00.27" />
                    <SPLIT distance="1400" swimtime="00:28:02.13" />
                    <SPLIT distance="1450" swimtime="00:29:04.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O7 - Przeszkadzanie innemu zawodnikowi (przez wypłynięcie na tor zajmowany przez innego zawodnika lub w inny sposób) (Time: 9:17)" eventid="1205" reactiontime="+78" status="DSQ" swimtime="00:00:52.45" resultid="3842" heatid="8954" lane="5" entrytime="00:01:50.00" />
                <RESULT eventid="1273" points="145" reactiontime="+91" swimtime="00:01:25.52" resultid="3843" heatid="8988" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="78" reactiontime="+74" swimtime="00:01:54.13" resultid="3844" heatid="9080" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="120" reactiontime="+86" swimtime="00:03:21.35" resultid="3845" heatid="9096" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="100" swimtime="00:01:32.69" />
                    <SPLIT distance="150" swimtime="00:02:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="110" reactiontime="+81" swimtime="00:00:52.56" resultid="3846" heatid="9161" lane="9" entrytime="00:00:53.00" />
                <RESULT eventid="1744" points="110" reactiontime="+92" swimtime="00:07:22.39" resultid="3847" heatid="9183" lane="2" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                    <SPLIT distance="100" swimtime="00:01:42.96" />
                    <SPLIT distance="150" swimtime="00:02:39.30" />
                    <SPLIT distance="200" swimtime="00:03:36.73" />
                    <SPLIT distance="250" swimtime="00:04:34.58" />
                    <SPLIT distance="300" swimtime="00:05:32.10" />
                    <SPLIT distance="350" swimtime="00:06:30.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="3914">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1079" points="486" reactiontime="+69" swimtime="00:00:25.76" resultid="3915" heatid="8911" lane="4" entrytime="00:00:26.50" />
                <RESULT eventid="1113" points="449" reactiontime="+82" swimtime="00:02:23.14" resultid="3916" heatid="8930" lane="1" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:01:07.93" />
                    <SPLIT distance="150" swimtime="00:01:49.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="445" reactiontime="+62" swimtime="00:00:29.09" resultid="3917" heatid="8963" lane="4" entrytime="00:00:30.00" />
                <RESULT comment="Rekord Polski" eventid="1341" points="441" reactiontime="+94" swimtime="00:02:22.58" resultid="3918" heatid="9030" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:08.62" />
                    <SPLIT distance="150" swimtime="00:01:45.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1440" points="513" reactiontime="+73" swimtime="00:00:27.23" resultid="3919" heatid="9071" lane="6" entrytime="00:00:27.90" />
                <RESULT eventid="1474" points="454" reactiontime="+61" swimtime="00:01:03.64" resultid="3920" heatid="9086" lane="5" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1613" points="488" reactiontime="+76" swimtime="00:01:01.49" resultid="3921" heatid="9136" lane="7" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="3869">
              <RESULTS>
                <RESULT eventid="1079" points="123" reactiontime="+116" swimtime="00:00:40.71" resultid="3870" heatid="8897" lane="1" entrytime="00:00:40.18" />
                <RESULT eventid="1165" points="159" reactiontime="+118" swimtime="00:26:09.10" resultid="3871" heatid="8942" lane="2" entrytime="00:26:33.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.63" />
                    <SPLIT distance="100" swimtime="00:01:37.21" />
                    <SPLIT distance="150" swimtime="00:02:31.96" />
                    <SPLIT distance="200" swimtime="00:03:25.77" />
                    <SPLIT distance="250" swimtime="00:04:19.68" />
                    <SPLIT distance="300" swimtime="00:05:12.95" />
                    <SPLIT distance="350" swimtime="00:06:06.01" />
                    <SPLIT distance="400" swimtime="00:06:58.92" />
                    <SPLIT distance="450" swimtime="00:07:51.61" />
                    <SPLIT distance="500" swimtime="00:08:44.22" />
                    <SPLIT distance="550" swimtime="00:09:36.92" />
                    <SPLIT distance="600" swimtime="00:10:28.29" />
                    <SPLIT distance="650" swimtime="00:11:20.67" />
                    <SPLIT distance="700" swimtime="00:12:12.43" />
                    <SPLIT distance="750" swimtime="00:13:03.90" />
                    <SPLIT distance="800" swimtime="00:13:56.93" />
                    <SPLIT distance="850" swimtime="00:14:49.01" />
                    <SPLIT distance="900" swimtime="00:15:41.47" />
                    <SPLIT distance="950" swimtime="00:16:34.28" />
                    <SPLIT distance="1000" swimtime="00:17:26.42" />
                    <SPLIT distance="1050" swimtime="00:18:19.20" />
                    <SPLIT distance="1100" swimtime="00:19:12.76" />
                    <SPLIT distance="1150" swimtime="00:20:06.69" />
                    <SPLIT distance="1200" swimtime="00:20:59.41" />
                    <SPLIT distance="1250" swimtime="00:21:51.51" />
                    <SPLIT distance="1300" swimtime="00:22:44.23" />
                    <SPLIT distance="1350" swimtime="00:23:37.92" />
                    <SPLIT distance="1400" swimtime="00:24:30.24" />
                    <SPLIT distance="1450" swimtime="00:25:22.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="134" reactiontime="+113" swimtime="00:01:27.63" resultid="3872" heatid="8987" lane="5" entrytime="00:01:28.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="90" reactiontime="+114" swimtime="00:00:48.53" resultid="3873" heatid="9061" lane="8" entrytime="00:00:47.45" />
                <RESULT eventid="1508" points="151" reactiontime="+114" swimtime="00:03:06.50" resultid="3874" heatid="9096" lane="4" entrytime="00:03:08.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                    <SPLIT distance="100" swimtime="00:01:31.31" />
                    <SPLIT distance="150" swimtime="00:02:20.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="164" reactiontime="+113" swimtime="00:06:27.39" resultid="3875" heatid="9184" lane="6" entrytime="00:06:45.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                    <SPLIT distance="100" swimtime="00:01:31.11" />
                    <SPLIT distance="150" swimtime="00:02:20.70" />
                    <SPLIT distance="200" swimtime="00:03:09.98" />
                    <SPLIT distance="250" swimtime="00:03:59.58" />
                    <SPLIT distance="300" swimtime="00:04:49.82" />
                    <SPLIT distance="350" swimtime="00:05:39.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka - Skorykow" nation="POL" athleteid="3922">
              <RESULTS>
                <RESULT eventid="1062" points="391" reactiontime="+86" swimtime="00:00:31.78" resultid="3923" heatid="8890" lane="7" entrytime="00:00:32.71" />
                <RESULT eventid="1222" points="351" reactiontime="+90" swimtime="00:03:10.62" resultid="3924" heatid="8969" lane="8" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.46" />
                    <SPLIT distance="100" swimtime="00:01:31.36" />
                    <SPLIT distance="150" swimtime="00:02:20.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="341" reactiontime="+85" swimtime="00:01:21.10" resultid="3925" heatid="9004" lane="6" entrytime="00:01:25.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="374" reactiontime="+87" swimtime="00:01:26.53" resultid="3926" heatid="9041" lane="2" entrytime="00:01:29.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="405" reactiontime="+82" swimtime="00:00:38.92" resultid="3927" heatid="9156" lane="4" entrytime="00:00:41.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-19" firstname="Marcin" gender="M" lastname="Giejsztowt" nation="POL" athleteid="3876">
              <RESULTS>
                <RESULT eventid="1079" points="334" reactiontime="+76" swimtime="00:00:29.20" resultid="3877" heatid="8903" lane="4" entrytime="00:00:30.65" />
                <RESULT eventid="1165" points="354" reactiontime="+82" swimtime="00:20:00.88" resultid="3878" heatid="8944" lane="5" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:13.73" />
                    <SPLIT distance="150" swimtime="00:01:52.31" />
                    <SPLIT distance="200" swimtime="00:02:31.54" />
                    <SPLIT distance="250" swimtime="00:03:11.52" />
                    <SPLIT distance="300" swimtime="00:03:51.47" />
                    <SPLIT distance="350" swimtime="00:04:31.84" />
                    <SPLIT distance="400" swimtime="00:05:12.30" />
                    <SPLIT distance="450" swimtime="00:05:52.91" />
                    <SPLIT distance="500" swimtime="00:06:33.82" />
                    <SPLIT distance="550" swimtime="00:07:14.52" />
                    <SPLIT distance="600" swimtime="00:07:55.04" />
                    <SPLIT distance="650" swimtime="00:08:35.98" />
                    <SPLIT distance="700" swimtime="00:09:16.10" />
                    <SPLIT distance="750" swimtime="00:09:57.14" />
                    <SPLIT distance="800" swimtime="00:10:37.58" />
                    <SPLIT distance="850" swimtime="00:11:18.84" />
                    <SPLIT distance="900" swimtime="00:11:59.09" />
                    <SPLIT distance="950" swimtime="00:12:40.03" />
                    <SPLIT distance="1000" swimtime="00:13:20.71" />
                    <SPLIT distance="1050" swimtime="00:14:01.57" />
                    <SPLIT distance="1100" swimtime="00:14:42.23" />
                    <SPLIT distance="1150" swimtime="00:15:23.54" />
                    <SPLIT distance="1200" swimtime="00:16:04.05" />
                    <SPLIT distance="1250" swimtime="00:16:44.49" />
                    <SPLIT distance="1300" swimtime="00:17:25.82" />
                    <SPLIT distance="1350" swimtime="00:18:06.63" />
                    <SPLIT distance="1400" swimtime="00:18:46.05" />
                    <SPLIT distance="1450" swimtime="00:19:25.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="344" reactiontime="+79" swimtime="00:01:04.13" resultid="3879" heatid="8993" lane="1" entrytime="00:01:06.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="322" reactiontime="+84" swimtime="00:00:31.78" resultid="3880" heatid="9066" lane="2" entrytime="00:00:32.55" />
                <RESULT eventid="1508" points="343" reactiontime="+77" swimtime="00:02:21.95" resultid="3881" heatid="9101" lane="9" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:08.78" />
                    <SPLIT distance="150" swimtime="00:01:46.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="339" reactiontime="+84" swimtime="00:05:04.33" resultid="3882" heatid="9188" lane="8" entrytime="00:05:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:10.13" />
                    <SPLIT distance="150" swimtime="00:01:48.67" />
                    <SPLIT distance="200" swimtime="00:02:27.64" />
                    <SPLIT distance="250" swimtime="00:03:06.92" />
                    <SPLIT distance="300" swimtime="00:03:46.18" />
                    <SPLIT distance="350" swimtime="00:04:25.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-07" firstname="Andrzej" gender="M" lastname="Lewandowski" nation="POL" athleteid="3894">
              <RESULTS>
                <RESULT eventid="1079" points="231" reactiontime="+85" swimtime="00:00:33.00" resultid="3895" heatid="8902" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="1205" points="176" reactiontime="+74" swimtime="00:00:39.63" resultid="3896" heatid="8957" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1273" points="225" reactiontime="+87" swimtime="00:01:13.87" resultid="3897" heatid="8990" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="271" reactiontime="+97" swimtime="00:01:25.87" resultid="3898" heatid="9046" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="183" reactiontime="+89" swimtime="00:02:54.94" resultid="3899" heatid="9094" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="324" reactiontime="+85" swimtime="00:00:36.76" resultid="3900" heatid="9167" lane="9" entrytime="00:00:38.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-12-28" firstname="Giovanni" gender="M" lastname="Moreno" nation="POL" athleteid="3795">
              <RESULTS>
                <RESULT eventid="1307" points="298" reactiontime="+83" swimtime="00:01:15.78" resultid="3796" heatid="9014" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="351" reactiontime="+77" swimtime="00:01:18.80" resultid="3797" heatid="9051" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="258" reactiontime="+75" swimtime="00:00:34.20" resultid="3798" heatid="9065" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1681" points="388" reactiontime="+77" swimtime="00:00:34.60" resultid="3799" heatid="9169" lane="0" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="3963">
              <RESULTS>
                <RESULT eventid="1113" points="309" reactiontime="+88" swimtime="00:02:42.03" resultid="3964" heatid="8927" lane="8" entrytime="00:02:48.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:15.14" />
                    <SPLIT distance="150" swimtime="00:02:06.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="344" reactiontime="+95" swimtime="00:01:04.08" resultid="3965" heatid="8989" lane="0" entrytime="00:01:15.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="317" reactiontime="+91" swimtime="00:01:14.25" resultid="3966" heatid="9014" lane="4" entrytime="00:01:15.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="350" reactiontime="+95" swimtime="00:02:21.00" resultid="3967" heatid="9101" lane="2" entrytime="00:02:22.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:44.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="301" reactiontime="+76" swimtime="00:02:38.20" resultid="3968" heatid="9147" lane="4" entrytime="00:02:42.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:17.47" />
                    <SPLIT distance="150" swimtime="00:01:57.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="3823">
              <RESULTS>
                <RESULT eventid="1079" points="49" reactiontime="+121" swimtime="00:00:55.05" resultid="3824" heatid="8895" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1113" points="48" reactiontime="+121" swimtime="00:05:00.11" resultid="3825" heatid="8921" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.09" />
                    <SPLIT distance="100" swimtime="00:02:38.92" />
                    <SPLIT distance="150" swimtime="00:03:49.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="63" reactiontime="+123" swimtime="00:05:01.65" resultid="3826" heatid="8972" lane="9" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.39" />
                    <SPLIT distance="100" swimtime="00:02:30.09" />
                    <SPLIT distance="150" swimtime="00:03:49.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="56" reactiontime="+122" swimtime="00:02:12.33" resultid="3827" heatid="9008" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="62" reactiontime="+123" swimtime="00:02:20.00" resultid="3828" heatid="9044" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="29" reactiontime="+120" swimtime="00:01:10.75" resultid="3829" heatid="9060" lane="8" entrytime="00:01:30.00" />
                <RESULT eventid="1647" points="42" reactiontime="+81" swimtime="00:05:04.27" resultid="3830" heatid="9143" lane="3" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.16" />
                    <SPLIT distance="100" swimtime="00:02:31.25" />
                    <SPLIT distance="150" swimtime="00:03:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="85" reactiontime="+130" swimtime="00:00:57.21" resultid="3831" heatid="9160" lane="7" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-10" firstname="Katarzyna" gender="F" lastname="Czarnecka" nation="POL" athleteid="3864">
              <RESULTS>
                <RESULT eventid="1062" points="373" reactiontime="+74" swimtime="00:00:32.27" resultid="3865" heatid="8889" lane="4" entrytime="00:00:33.70" />
                <RESULT eventid="1222" points="309" reactiontime="+75" swimtime="00:03:18.89" resultid="3866" heatid="8969" lane="5" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.05" />
                    <SPLIT distance="100" swimtime="00:01:37.27" />
                    <SPLIT distance="150" swimtime="00:02:29.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="348" reactiontime="+74" swimtime="00:01:28.58" resultid="3867" heatid="9040" lane="5" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="413" reactiontime="+74" swimtime="00:00:38.66" resultid="3868" heatid="9157" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-10-19" firstname="Emilia" gender="F" lastname="Sączyńska" nation="POL" athleteid="3958">
              <RESULTS>
                <RESULT eventid="1187" points="337" reactiontime="+79" swimtime="00:00:36.86" resultid="3959" heatid="8952" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1324" points="255" reactiontime="+98" swimtime="00:03:08.51" resultid="3960" heatid="9024" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:27.57" />
                    <SPLIT distance="150" swimtime="00:02:18.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="328" reactiontime="+77" swimtime="00:01:19.75" resultid="3961" heatid="9077" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="366" reactiontime="+77" swimtime="00:02:46.67" resultid="3962" heatid="9140" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:20.58" />
                    <SPLIT distance="150" swimtime="00:02:04.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="3789">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1079" points="456" reactiontime="+73" swimtime="00:00:26.31" resultid="3790" heatid="8910" lane="4" entrytime="00:00:26.81" />
                <RESULT comment="Rekord Polski" eventid="1273" points="481" reactiontime="+76" swimtime="00:00:57.33" resultid="3791" heatid="8987" lane="4" entrytime="00:01:28.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1307" points="440" reactiontime="+79" swimtime="00:01:06.59" resultid="3792" heatid="9019" lane="1" entrytime="00:01:07.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="439" reactiontime="+80" swimtime="00:02:10.69" resultid="3793" heatid="9104" lane="3" entrytime="00:02:09.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                    <SPLIT distance="150" swimtime="00:01:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1681" points="412" reactiontime="+80" swimtime="00:00:33.91" resultid="3794" heatid="9170" lane="3" entrytime="00:00:34.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-25" firstname="Barbara" gender="F" lastname="Ropa" nation="POL" athleteid="3800" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="1381" points="417" reactiontime="+79" swimtime="00:02:01.06" resultid="8606" heatid="9035" lane="0" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:07.39" />
                    <SPLIT distance="150" swimtime="00:01:34.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3901" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="3848" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="4008" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="3890" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="10">
              <RESULTS>
                <RESULT eventid="1381" points="337" reactiontime="+92" swimtime="00:02:10.05" resultid="8607" heatid="9033" lane="5" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                    <SPLIT distance="100" swimtime="00:01:11.37" />
                    <SPLIT distance="150" swimtime="00:01:42.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3939" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="3795" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="3876" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="3934" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="13">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1548" points="491" reactiontime="+73" swimtime="00:01:44.66" resultid="8610" heatid="9112" lane="9" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.02" />
                    <SPLIT distance="100" swimtime="00:00:51.91" />
                    <SPLIT distance="150" swimtime="00:01:18.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4008" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3832" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="3855" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="3914" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="14">
              <RESULTS>
                <RESULT eventid="1548" points="388" reactiontime="+83" swimtime="00:01:53.24" resultid="8611" heatid="9111" lane="7" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                    <SPLIT distance="100" swimtime="00:00:56.21" />
                    <SPLIT distance="150" swimtime="00:01:26.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3934" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="3901" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3996" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3890" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="15">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="8612" heatid="9110" lane="7" entrytime="00:02:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3814" number="1" />
                    <RELAYPOSITION athleteid="3988" number="2" />
                    <RELAYPOSITION athleteid="3939" number="3" />
                    <RELAYPOSITION athleteid="3909" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="7">
              <RESULTS>
                <RESULT eventid="1358" points="285" reactiontime="+76" swimtime="00:02:38.09" resultid="8604" heatid="9031" lane="4" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                    <SPLIT distance="100" swimtime="00:01:27.57" />
                    <SPLIT distance="150" swimtime="00:02:06.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3958" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4014" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="3946" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4020" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="11">
              <RESULTS>
                <RESULT eventid="1525" points="430" reactiontime="+79" swimtime="00:02:04.85" resultid="8608" heatid="9108" lane="2" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:03.24" />
                    <SPLIT distance="150" swimtime="00:01:37.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3864" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="3922" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4020" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3982" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="296" reactiontime="+78" swimtime="00:02:03.89" resultid="8599" heatid="8934" lane="5" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                    <SPLIT distance="100" swimtime="00:01:07.65" />
                    <SPLIT distance="150" swimtime="00:01:39.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3855" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4014" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3864" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4008" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="3">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1698" points="392" reactiontime="+88" swimtime="00:02:03.58" resultid="8600" heatid="9176" lane="1" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:01:08.28" />
                    <SPLIT distance="150" swimtime="00:01:37.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4008" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3922" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3982" number="3" reactiontime="+10" />
                    <RELAYPOSITION athleteid="3789" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1698" points="307" reactiontime="+85" swimtime="00:02:14.07" resultid="8601" heatid="9176" lane="6" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="100" swimtime="00:01:12.50" />
                    <SPLIT distance="150" swimtime="00:01:43.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3958" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="3890" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="3901" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="3809" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="1698" points="245" reactiontime="+80" swimtime="00:02:24.57" resultid="8603" heatid="9175" lane="2" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:05.41" />
                    <SPLIT distance="150" swimtime="00:01:44.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3832" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3795" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4020" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="4014" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="4982" name="Weteran  Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" phone="604 522 654" street="ŚW.JANA   4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE birthdate="1947-05-23" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" license="502611100004" athleteid="6362">
              <RESULTS>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="6363" heatid="8949" lane="8" entrytime="00:00:56.00" />
                <RESULT eventid="1664" points="176" reactiontime="+91" swimtime="00:00:51.36" resultid="6364" heatid="9153" lane="8" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-11-06" firstname="Joanna" gender="F" lastname="Sulewska - Bielak" nation="POL" athleteid="6406">
              <RESULTS>
                <RESULT eventid="1290" points="341" reactiontime="+91" swimtime="00:01:21.12" resultid="6407" heatid="9005" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="6408" heatid="9057" lane="8" entrytime="00:00:36.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="502611200005" athleteid="6358">
              <RESULTS>
                <RESULT eventid="1079" points="120" reactiontime="+108" swimtime="00:00:41.05" resultid="6359" heatid="8897" lane="3" entrytime="00:00:39.65" />
                <RESULT eventid="1205" points="70" reactiontime="+85" swimtime="00:00:53.84" resultid="6360" heatid="8955" lane="4" entrytime="00:00:54.00" />
                <RESULT eventid="1440" points="88" reactiontime="+101" swimtime="00:00:48.83" resultid="6361" heatid="9061" lane="3" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="502611200008" athleteid="6374">
              <RESULTS>
                <RESULT eventid="1079" points="282" reactiontime="+80" swimtime="00:00:30.88" resultid="6375" heatid="8902" lane="1" entrytime="00:00:31.50" />
                <RESULT eventid="1205" points="195" reactiontime="+74" swimtime="00:00:38.29" resultid="6376" heatid="8958" lane="3" entrytime="00:00:38.69" />
                <RESULT eventid="1440" points="213" reactiontime="+86" swimtime="00:00:36.45" resultid="6377" heatid="9065" lane="3" entrytime="00:00:33.50" />
                <RESULT eventid="1474" points="190" reactiontime="+89" swimtime="00:01:25.02" resultid="6378" heatid="9082" lane="2" entrytime="00:01:25.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="193" reactiontime="+64" swimtime="00:03:03.48" resultid="6379" heatid="9146" lane="7" entrytime="00:03:14.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:01:28.87" />
                    <SPLIT distance="150" swimtime="00:02:16.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-07-16" firstname="Ewald" gender="M" lastname="Bastek" nation="POL" license="502611200001" athleteid="6380">
              <RESULTS>
                <RESULT eventid="1113" points="132" reactiontime="+122" swimtime="00:03:34.81" resultid="6381" heatid="8922" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.38" />
                    <SPLIT distance="100" swimtime="00:01:48.26" />
                    <SPLIT distance="150" swimtime="00:02:47.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="150" reactiontime="+116" swimtime="00:01:35.18" resultid="6382" heatid="9010" lane="0" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1578" points="136" reactiontime="+114" swimtime="00:07:37.27" resultid="6383" heatid="9117" lane="1" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.64" />
                    <SPLIT distance="100" swimtime="00:01:57.44" />
                    <SPLIT distance="150" swimtime="00:02:59.18" />
                    <SPLIT distance="200" swimtime="00:03:58.60" />
                    <SPLIT distance="250" swimtime="00:05:00.56" />
                    <SPLIT distance="300" swimtime="00:06:02.78" />
                    <SPLIT distance="350" swimtime="00:06:52.45" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1744" points="152" reactiontime="+99" swimtime="00:06:37.09" resultid="6384" heatid="9184" lane="8" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                    <SPLIT distance="150" swimtime="00:02:22.59" />
                    <SPLIT distance="200" swimtime="00:03:14.31" />
                    <SPLIT distance="250" swimtime="00:04:05.15" />
                    <SPLIT distance="300" swimtime="00:04:57.38" />
                    <SPLIT distance="350" swimtime="00:05:48.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="502611100009" athleteid="6391">
              <RESULTS>
                <RESULT eventid="1147" points="464" reactiontime="+88" swimtime="00:10:19.11" resultid="6392" heatid="8939" lane="3" entrytime="00:10:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:50.17" />
                    <SPLIT distance="200" swimtime="00:02:29.00" />
                    <SPLIT distance="250" swimtime="00:03:07.89" />
                    <SPLIT distance="300" swimtime="00:03:46.71" />
                    <SPLIT distance="350" swimtime="00:04:25.77" />
                    <SPLIT distance="400" swimtime="00:05:04.83" />
                    <SPLIT distance="450" swimtime="00:05:44.21" />
                    <SPLIT distance="500" swimtime="00:06:23.55" />
                    <SPLIT distance="550" swimtime="00:07:03.12" />
                    <SPLIT distance="600" swimtime="00:07:42.51" />
                    <SPLIT distance="650" swimtime="00:08:21.72" />
                    <SPLIT distance="700" swimtime="00:09:01.50" />
                    <SPLIT distance="750" swimtime="00:09:41.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="411" reactiontime="+92" swimtime="00:03:00.99" resultid="6393" heatid="8970" lane="4" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:01:26.67" />
                    <SPLIT distance="150" swimtime="00:02:13.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="420" reactiontime="+88" swimtime="00:01:23.23" resultid="6394" heatid="9042" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="443" reactiontime="+95" swimtime="00:02:25.32" resultid="6395" heatid="9093" lane="1" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:10.33" />
                    <SPLIT distance="150" swimtime="00:01:48.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="454" reactiontime="+97" swimtime="00:05:05.03" resultid="6396" heatid="9181" lane="2" entrytime="00:05:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:01:50.76" />
                    <SPLIT distance="200" swimtime="00:02:29.76" />
                    <SPLIT distance="250" swimtime="00:03:08.87" />
                    <SPLIT distance="300" swimtime="00:03:48.14" />
                    <SPLIT distance="350" swimtime="00:04:26.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="502611100001" athleteid="6385">
              <RESULTS>
                <RESULT eventid="1062" points="248" reactiontime="+86" swimtime="00:00:36.96" resultid="6386" heatid="8888" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1187" points="190" reactiontime="+70" swimtime="00:00:44.58" resultid="6387" heatid="8950" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1256" points="214" reactiontime="+81" swimtime="00:01:25.27" resultid="6388" heatid="8981" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="122" reactiontime="+87" swimtime="00:00:49.07" resultid="6389" heatid="9055" lane="1" entrytime="00:00:48.00" />
                <RESULT eventid="1630" points="151" reactiontime="+71" swimtime="00:03:43.70" resultid="6390" heatid="9139" lane="7" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.09" />
                    <SPLIT distance="100" swimtime="00:01:50.67" />
                    <SPLIT distance="150" swimtime="00:02:48.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="502611100002" athleteid="6369">
              <RESULTS>
                <RESULT eventid="1222" points="183" reactiontime="+115" swimtime="00:03:56.93" resultid="6370" heatid="8968" lane="1" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.13" />
                    <SPLIT distance="100" swimtime="00:01:54.74" />
                    <SPLIT distance="150" swimtime="00:02:56.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="177" reactiontime="+105" swimtime="00:01:50.92" resultid="6371" heatid="9039" lane="0" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="121" reactiontime="+98" swimtime="00:01:50.24" resultid="6372" heatid="9124" lane="4" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="162" reactiontime="+99" swimtime="00:00:52.74" resultid="6373" heatid="9154" lane="9" entrytime="00:00:49.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" license="502611200004" athleteid="6354">
              <RESULTS>
                <RESULT eventid="1205" points="147" reactiontime="+71" swimtime="00:00:42.05" resultid="6355" heatid="8957" lane="6" entrytime="00:00:41.46" />
                <RESULT eventid="1474" points="123" reactiontime="+72" swimtime="00:01:38.26" resultid="6356" heatid="9081" lane="1" entrytime="00:01:37.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="117" reactiontime="+72" swimtime="00:03:36.72" resultid="6357" heatid="9145" lane="6" entrytime="00:03:39.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                    <SPLIT distance="100" swimtime="00:01:43.79" />
                    <SPLIT distance="150" swimtime="00:02:40.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="502611200002" athleteid="6365">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1239" points="189" reactiontime="+107" swimtime="00:03:29.62" resultid="6366" heatid="8973" lane="6" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.62" />
                    <SPLIT distance="100" swimtime="00:01:41.59" />
                    <SPLIT distance="150" swimtime="00:02:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="184" reactiontime="+99" swimtime="00:01:37.67" resultid="6367" heatid="9046" lane="0" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="170" reactiontime="+95" swimtime="00:00:45.52" resultid="6368" heatid="9163" lane="9" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-28" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="502611200007" athleteid="6397">
              <RESULTS>
                <RESULT eventid="1079" points="178" reactiontime="+88" swimtime="00:00:36.01" resultid="6398" heatid="8903" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1273" points="200" reactiontime="+90" swimtime="00:01:16.72" resultid="6399" heatid="8989" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="238" reactiontime="+89" swimtime="00:00:35.17" resultid="6400" heatid="9064" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-09-27" firstname="Przemysław" gender="M" lastname="Pindor" nation="POL" athleteid="6412">
              <RESULTS>
                <RESULT eventid="1508" points="281" reactiontime="+74" swimtime="00:02:31.58" resultid="6413" heatid="9100" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="233" reactiontime="+82" swimtime="00:05:44.51" resultid="6414" heatid="9190" lane="1" entrytime="00:04:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:16.81" />
                    <SPLIT distance="150" swimtime="00:01:59.70" />
                    <SPLIT distance="200" swimtime="00:02:43.70" />
                    <SPLIT distance="250" swimtime="00:03:29.63" />
                    <SPLIT distance="300" swimtime="00:04:16.05" />
                    <SPLIT distance="350" swimtime="00:05:02.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-05" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" license="502611100005" athleteid="6401">
              <RESULTS>
                <RESULT eventid="1062" points="178" reactiontime="+100" swimtime="00:00:41.27" resultid="6402" heatid="8887" lane="7" entrytime="00:00:42.50" />
                <RESULT eventid="1256" points="148" reactiontime="+105" swimtime="00:01:36.43" resultid="6403" heatid="8980" lane="9" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="105" reactiontime="+106" swimtime="00:03:54.22" resultid="6404" heatid="9089" lane="5" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.49" />
                    <SPLIT distance="100" swimtime="00:01:52.28" />
                    <SPLIT distance="150" swimtime="00:02:53.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="82" reactiontime="+87" swimtime="00:04:33.36" resultid="6405" heatid="9138" lane="3" entrytime="00:04:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.37" />
                    <SPLIT distance="100" swimtime="00:02:15.30" />
                    <SPLIT distance="150" swimtime="00:03:26.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-02-18" firstname="Genowefa" gender="F" lastname="Drużyńska" nation="POL" athleteid="6409">
              <RESULTS>
                <RESULT eventid="1388" points="111" reactiontime="+98" swimtime="00:02:09.41" resultid="6410" heatid="9038" lane="0" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="140" reactiontime="+105" swimtime="00:00:55.37" resultid="6411" heatid="9152" lane="4" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="158" reactiontime="+88" swimtime="00:02:47.14" resultid="6418" heatid="9032" lane="6" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.33" />
                    <SPLIT distance="100" swimtime="00:01:31.70" />
                    <SPLIT distance="150" swimtime="00:02:07.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6380" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="6365" number="2" reactiontime="+84" />
                    <RELAYPOSITION athleteid="6397" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="6358" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1548" points="170" reactiontime="+93" swimtime="00:02:29.02" resultid="6420" heatid="9109" lane="6" entrytime="00:02:34.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:17.34" />
                    <SPLIT distance="150" swimtime="00:01:55.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6358" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="6365" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="6380" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="6397" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="217" reactiontime="+70" swimtime="00:02:52.97" resultid="6417" heatid="9031" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:37.30" />
                    <SPLIT distance="150" swimtime="00:02:12.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6385" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="6369" number="2" />
                    <RELAYPOSITION athleteid="6391" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="6401" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="5">
              <RESULTS>
                <RESULT eventid="1525" points="196" reactiontime="+86" swimtime="00:02:42.00" resultid="6419" heatid="9108" lane="7" entrytime="00:02:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:26.34" />
                    <SPLIT distance="150" swimtime="00:02:08.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6385" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="6369" number="2" reactiontime="+74" />
                    <RELAYPOSITION athleteid="6401" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="6391" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="137" reactiontime="+83" swimtime="00:02:40.00" resultid="6415" heatid="8933" lane="8" entrytime="00:02:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:01:22.73" />
                    <SPLIT distance="150" swimtime="00:02:00.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6385" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="6362" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="6380" number="3" reactiontime="+90" />
                    <RELAYPOSITION athleteid="6358" number="4" reactiontime="+78" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="207" reactiontime="+90" swimtime="00:02:19.54" resultid="6416" heatid="8933" lane="0" entrytime="00:02:47.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:11.64" />
                    <SPLIT distance="150" swimtime="00:01:47.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6397" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="6401" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="6354" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="6391" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="1698" points="148" reactiontime="+76" swimtime="00:02:50.76" resultid="6421" heatid="9174" lane="6" entrytime="00:02:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                    <SPLIT distance="100" swimtime="00:01:38.19" />
                    <SPLIT distance="150" swimtime="00:02:13.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6385" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="6369" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="6397" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="6380" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WKSSLA" nation="POL" region="DOL" clubid="5772" name="WKS ŚlĄSK">
          <CONTACT city="BIELANY WROCLAWSK" email="BIURO@PLYWANIEWROCLAW.PL" name="wERESZCZYŃSKI" phone="723897862" state="DOL" street="KŁODZKA" zip="55-040" />
          <ATHLETES>
            <ATHLETE birthdate="1975-01-13" firstname="Cezary" gender="M" lastname="Wereszczyński" nation="POL" athleteid="5798">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="5799" heatid="8910" lane="3" entrytime="00:00:26.98" />
                <RESULT eventid="1440" points="349" reactiontime="+84" swimtime="00:00:30.96" resultid="5800" heatid="9070" lane="8" entrytime="00:00:29.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-03-17" firstname="Maciej" gender="M" lastname="Dąbrowski" nation="POL" athleteid="5814">
              <RESULTS>
                <RESULT eventid="1079" points="317" reactiontime="+98" swimtime="00:00:29.69" resultid="5815" heatid="8907" lane="7" entrytime="00:00:28.95" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="5816" heatid="8927" lane="7" entrytime="00:02:47.00" />
                <RESULT eventid="1205" points="281" reactiontime="+79" swimtime="00:00:33.91" resultid="5817" heatid="8961" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1307" points="305" reactiontime="+98" swimtime="00:01:15.22" resultid="5818" heatid="9015" lane="3" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="279" reactiontime="+93" swimtime="00:00:33.36" resultid="5819" heatid="9065" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="5820" heatid="9083" lane="6" entrytime="00:01:17.00" />
                <RESULT eventid="1613" points="224" reactiontime="+114" swimtime="00:01:19.74" resultid="5821" heatid="9132" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="251" reactiontime="+84" swimtime="00:02:48.16" resultid="5822" heatid="9147" lane="2" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                    <SPLIT distance="100" swimtime="00:01:22.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Wojciech" gender="M" lastname="Sobczak" nation="POL" athleteid="5807">
              <RESULTS>
                <RESULT eventid="1113" points="186" reactiontime="+91" swimtime="00:03:11.96" resultid="5808" heatid="8924" lane="9" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:33.33" />
                    <SPLIT distance="150" swimtime="00:02:29.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="218" reactiontime="+117" swimtime="00:23:31.21" resultid="5809" heatid="8943" lane="1" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:22.38" />
                    <SPLIT distance="150" swimtime="00:02:06.55" />
                    <SPLIT distance="200" swimtime="00:02:51.58" />
                    <SPLIT distance="250" swimtime="00:03:37.99" />
                    <SPLIT distance="300" swimtime="00:04:24.77" />
                    <SPLIT distance="350" swimtime="00:05:11.42" />
                    <SPLIT distance="400" swimtime="00:05:57.87" />
                    <SPLIT distance="450" swimtime="00:06:45.02" />
                    <SPLIT distance="500" swimtime="00:07:33.38" />
                    <SPLIT distance="550" swimtime="00:08:21.44" />
                    <SPLIT distance="600" swimtime="00:09:09.28" />
                    <SPLIT distance="650" swimtime="00:09:58.56" />
                    <SPLIT distance="700" swimtime="00:10:45.91" />
                    <SPLIT distance="750" swimtime="00:11:33.70" />
                    <SPLIT distance="800" swimtime="00:12:22.45" />
                    <SPLIT distance="850" swimtime="00:13:10.09" />
                    <SPLIT distance="900" swimtime="00:13:57.40" />
                    <SPLIT distance="950" swimtime="00:14:45.62" />
                    <SPLIT distance="1000" swimtime="00:15:33.41" />
                    <SPLIT distance="1050" swimtime="00:16:21.13" />
                    <SPLIT distance="1100" swimtime="00:17:08.30" />
                    <SPLIT distance="1150" swimtime="00:17:56.21" />
                    <SPLIT distance="1200" swimtime="00:18:43.16" />
                    <SPLIT distance="1250" swimtime="00:19:31.16" />
                    <SPLIT distance="1300" swimtime="00:20:18.31" />
                    <SPLIT distance="1350" swimtime="00:21:06.90" />
                    <SPLIT distance="1400" swimtime="00:21:55.46" />
                    <SPLIT distance="1450" swimtime="00:22:44.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="194" reactiontime="+114" swimtime="00:03:27.79" resultid="5810" heatid="8973" lane="0" entrytime="00:03:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.68" />
                    <SPLIT distance="100" swimtime="00:01:40.46" />
                    <SPLIT distance="150" swimtime="00:02:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="116" reactiontime="+93" swimtime="00:03:42.13" resultid="5811" heatid="9027" lane="9" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                    <SPLIT distance="100" swimtime="00:01:44.82" />
                    <SPLIT distance="150" swimtime="00:02:47.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="118" reactiontime="+107" swimtime="00:01:38.67" resultid="5812" heatid="9130" lane="2" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="227" reactiontime="+98" swimtime="00:05:47.60" resultid="5813" heatid="9186" lane="8" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:20.65" />
                    <SPLIT distance="150" swimtime="00:02:03.61" />
                    <SPLIT distance="200" swimtime="00:02:47.95" />
                    <SPLIT distance="250" swimtime="00:03:32.59" />
                    <SPLIT distance="300" swimtime="00:04:18.03" />
                    <SPLIT distance="350" swimtime="00:05:03.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-09-15" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="5790">
              <RESULTS>
                <RESULT eventid="1062" points="218" reactiontime="+90" swimtime="00:00:38.59" resultid="5791" heatid="8888" lane="7" entrytime="00:00:38.88" />
                <RESULT eventid="1096" points="152" reactiontime="+86" swimtime="00:03:47.93" resultid="5792" heatid="8917" lane="1" entrytime="00:03:47.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.43" />
                    <SPLIT distance="100" swimtime="00:01:49.97" />
                    <SPLIT distance="150" swimtime="00:02:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="5793" heatid="8968" lane="2" entrytime="00:03:52.72" />
                <RESULT eventid="1290" points="201" reactiontime="+83" swimtime="00:01:36.66" resultid="5794" heatid="9002" lane="5" entrytime="00:01:41.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="209" reactiontime="+90" swimtime="00:01:45.01" resultid="5795" heatid="9039" lane="5" entrytime="00:01:41.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="157" reactiontime="+94" swimtime="00:03:25.31" resultid="5796" heatid="9090" lane="1" entrytime="00:03:18.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                    <SPLIT distance="100" swimtime="00:01:37.37" />
                    <SPLIT distance="150" swimtime="00:02:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="267" reactiontime="+83" swimtime="00:00:44.71" resultid="5797" heatid="9154" lane="4" entrytime="00:00:46.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-23" firstname="Agata" gender="F" lastname="Sobczak" nation="POL" athleteid="5784">
              <RESULTS>
                <RESULT eventid="1147" points="183" reactiontime="+119" swimtime="00:14:02.90" resultid="5785" heatid="8937" lane="2" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.99" />
                    <SPLIT distance="100" swimtime="00:01:37.39" />
                    <SPLIT distance="150" swimtime="00:02:29.27" />
                    <SPLIT distance="200" swimtime="00:03:21.49" />
                    <SPLIT distance="250" swimtime="00:04:12.98" />
                    <SPLIT distance="300" swimtime="00:06:00.28" />
                    <SPLIT distance="350" swimtime="00:06:54.99" />
                    <SPLIT distance="400" swimtime="00:07:48.98" />
                    <SPLIT distance="450" swimtime="00:08:42.55" />
                    <SPLIT distance="500" swimtime="00:09:36.92" />
                    <SPLIT distance="550" swimtime="00:10:30.35" />
                    <SPLIT distance="600" swimtime="00:11:23.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="129" reactiontime="+104" swimtime="00:03:56.57" resultid="5786" heatid="9023" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.66" />
                    <SPLIT distance="100" swimtime="00:01:52.12" />
                    <SPLIT distance="150" swimtime="00:02:55.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="183" reactiontime="+101" swimtime="00:03:14.87" resultid="5787" heatid="9090" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                    <SPLIT distance="100" swimtime="00:01:35.11" />
                    <SPLIT distance="150" swimtime="00:02:26.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="121" reactiontime="+107" swimtime="00:01:50.14" resultid="5788" heatid="9124" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="188" reactiontime="+89" swimtime="00:06:48.94" resultid="5789" heatid="9178" lane="3" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.10" />
                    <SPLIT distance="100" swimtime="00:01:38.16" />
                    <SPLIT distance="150" swimtime="00:02:29.87" />
                    <SPLIT distance="200" swimtime="00:03:22.11" />
                    <SPLIT distance="250" swimtime="00:04:14.59" />
                    <SPLIT distance="300" swimtime="00:05:07.30" />
                    <SPLIT distance="350" swimtime="00:05:59.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-19" firstname="Kinga" gender="F" lastname="Murawska" nation="POL" athleteid="5777">
              <RESULTS>
                <RESULT eventid="1096" points="168" reactiontime="+92" swimtime="00:03:40.46" resultid="5778" heatid="8917" lane="0" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                    <SPLIT distance="100" swimtime="00:01:47.08" />
                    <SPLIT distance="150" swimtime="00:02:48.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="184" reactiontime="+87" swimtime="00:03:56.37" resultid="5779" heatid="8967" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.19" />
                    <SPLIT distance="100" swimtime="00:01:54.28" />
                    <SPLIT distance="150" swimtime="00:02:55.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="163" reactiontime="+86" swimtime="00:01:43.70" resultid="5780" heatid="9003" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="173" reactiontime="+89" swimtime="00:07:45.48" resultid="5781" heatid="9113" lane="3" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.04" />
                    <SPLIT distance="100" swimtime="00:01:54.31" />
                    <SPLIT distance="150" swimtime="00:02:51.08" />
                    <SPLIT distance="200" swimtime="00:03:47.45" />
                    <SPLIT distance="250" swimtime="00:04:51.49" />
                    <SPLIT distance="300" swimtime="00:05:56.76" />
                    <SPLIT distance="350" swimtime="00:06:52.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="122" reactiontime="+89" swimtime="00:01:50.03" resultid="5782" heatid="9125" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="177" reactiontime="+90" swimtime="00:06:57.42" resultid="5783" heatid="9178" lane="6" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                    <SPLIT distance="100" swimtime="00:01:40.34" />
                    <SPLIT distance="150" swimtime="00:02:33.00" />
                    <SPLIT distance="200" swimtime="00:03:25.97" />
                    <SPLIT distance="250" swimtime="00:04:20.24" />
                    <SPLIT distance="300" swimtime="00:05:14.04" />
                    <SPLIT distance="350" swimtime="00:06:07.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-07" firstname="Radosław" gender="M" lastname="Stefurak" nation="POL" athleteid="5773">
              <RESULTS>
                <RESULT eventid="1239" points="285" reactiontime="+86" swimtime="00:03:02.94" resultid="5774" heatid="8976" lane="3" entrytime="00:03:00.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:25.12" />
                    <SPLIT distance="150" swimtime="00:02:13.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="284" reactiontime="+91" swimtime="00:01:24.60" resultid="5775" heatid="9049" lane="1" entrytime="00:01:25.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="232" reactiontime="+101" swimtime="00:02:41.55" resultid="5776" heatid="9098" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:01:59.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-23" firstname="Anna" gender="F" lastname="Głowiak" nation="POL" athleteid="5801">
              <RESULTS>
                <RESULT eventid="1062" points="358" reactiontime="+85" swimtime="00:00:32.71" resultid="5802" heatid="8890" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1290" points="259" reactiontime="+85" swimtime="00:01:28.85" resultid="5803" heatid="9004" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="272" reactiontime="+86" swimtime="00:01:36.14" resultid="5804" heatid="9039" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="5805" heatid="9126" lane="4" entrytime="00:01:16.00" />
                <RESULT eventid="1664" points="302" reactiontime="+87" swimtime="00:00:42.88" resultid="5806" heatid="9155" lane="4" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="299" reactiontime="+81" swimtime="00:02:03.47" resultid="5823" heatid="9110" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                    <SPLIT distance="100" swimtime="00:01:00.30" />
                    <SPLIT distance="150" swimtime="00:01:33.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5798" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="5773" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5807" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="5814" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="273" reactiontime="+86" swimtime="00:02:19.51" resultid="5824" heatid="9033" lane="3" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:52.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5814" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="5773" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="5807" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="5798" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1525" points="225" reactiontime="+86" swimtime="00:02:34.76" resultid="5825" heatid="9108" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:12.25" />
                    <SPLIT distance="150" swimtime="00:01:53.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5801" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="5790" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="5777" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="5784" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1358" points="203" reactiontime="+82" swimtime="00:02:56.92" resultid="5826" heatid="9031" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:25.79" />
                    <SPLIT distance="150" swimtime="00:02:17.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5801" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="5790" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="5777" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="5784" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="241" reactiontime="+102" swimtime="00:02:12.58" resultid="5827" heatid="8934" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:04.53" />
                    <SPLIT distance="150" swimtime="00:01:43.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5807" number="1" reactiontime="+102" />
                    <RELAYPOSITION athleteid="5801" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="5790" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="5814" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="205" reactiontime="+83" swimtime="00:02:33.43" resultid="5830" heatid="9174" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:28.68" />
                    <SPLIT distance="150" swimtime="00:02:01.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5801" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="5790" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="5814" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="5798" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="5828" heatid="8933" lane="6" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5807" number="1" />
                    <RELAYPOSITION athleteid="5777" number="2" />
                    <RELAYPOSITION athleteid="5784" number="3" />
                    <RELAYPOSITION athleteid="5773" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="5829" heatid="9174" lane="7" entrytime="00:02:45.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5807" number="1" />
                    <RELAYPOSITION athleteid="5773" number="2" />
                    <RELAYPOSITION athleteid="5777" number="3" />
                    <RELAYPOSITION athleteid="5784" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WIE" nation="POL" region="WIE" clubid="4968" name="Wojewódzki Sztab Wojskowy Poznań" shortname="Wojewódzki Sztab Wojskowy Pozn">
          <CONTACT city="Świdnica" email="horbacz.marcin@wp.pl" name="Horbacz" phone="603672717" state="LUB" street="Buchałów 12c" zip="66-008" />
          <ATHLETES>
            <ATHLETE birthdate="1981-01-01" firstname="Małgorzata" gender="F" lastname="Matkowska" nation="POL" athleteid="4969">
              <RESULTS>
                <RESULT eventid="1096" points="212" reactiontime="+98" swimtime="00:03:24.29" resultid="4970" heatid="8917" lane="6" entrytime="00:03:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:34.34" />
                    <SPLIT distance="150" swimtime="00:02:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="160" reactiontime="+107" swimtime="00:03:40.01" resultid="4971" heatid="9023" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                    <SPLIT distance="100" swimtime="00:01:47.63" />
                    <SPLIT distance="150" swimtime="00:02:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="192" reactiontime="+101" swimtime="00:07:29.92" resultid="4972" heatid="9113" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:01:37.00" />
                    <SPLIT distance="150" swimtime="00:02:39.35" />
                    <SPLIT distance="200" swimtime="00:03:39.56" />
                    <SPLIT distance="250" swimtime="00:04:42.28" />
                    <SPLIT distance="300" swimtime="00:05:45.67" />
                    <SPLIT distance="350" swimtime="00:06:39.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="4973" heatid="9123" lane="5" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="4974" heatid="9177" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2068" name="WOPR Tczew">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="2069">
              <RESULTS>
                <RESULT eventid="1079" points="449" reactiontime="+83" swimtime="00:00:26.44" resultid="2070" heatid="8913" lane="8" entrytime="00:00:26.00" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="2071" heatid="8929" lane="5" entrytime="00:02:30.00" />
                <RESULT eventid="1273" points="460" reactiontime="+82" swimtime="00:00:58.18" resultid="2072" heatid="8998" lane="7" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="455" reactiontime="+96" swimtime="00:01:12.25" resultid="2073" heatid="9053" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="418" reactiontime="+83" swimtime="00:02:12.80" resultid="2074" heatid="9104" lane="9" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:04.67" />
                    <SPLIT distance="150" swimtime="00:01:39.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="458" reactiontime="+90" swimtime="00:00:32.74" resultid="2075" heatid="9172" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="2076" heatid="9190" lane="6" entrytime="00:04:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-18" firstname="Marek" gender="M" lastname="Stuczyński" nation="POL" athleteid="2084">
              <RESULTS>
                <RESULT eventid="1079" points="517" reactiontime="+78" swimtime="00:00:25.23" resultid="2085" heatid="8913" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1307" points="491" reactiontime="+75" swimtime="00:01:04.21" resultid="2086" heatid="9019" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="504" reactiontime="+80" swimtime="00:01:09.87" resultid="2087" heatid="9053" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="535" reactiontime="+79" swimtime="00:00:31.09" resultid="2088" heatid="9172" lane="6" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="2077">
              <RESULTS>
                <RESULT eventid="1062" points="362" reactiontime="+96" swimtime="00:00:32.60" resultid="2078" heatid="8891" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1187" points="226" reactiontime="+89" swimtime="00:00:42.13" resultid="2079" heatid="8950" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1256" points="309" reactiontime="+102" swimtime="00:01:15.43" resultid="2080" heatid="8981" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="2081" heatid="9076" lane="0" entrytime="00:01:32.00" />
                <RESULT eventid="1491" points="262" reactiontime="+101" swimtime="00:02:53.01" resultid="2082" heatid="9091" lane="8" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:01:22.25" />
                    <SPLIT distance="150" swimtime="00:02:08.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="237" reactiontime="+89" swimtime="00:03:12.54" resultid="2083" heatid="9139" lane="3" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="100" swimtime="00:01:34.99" />
                    <SPLIT distance="150" swimtime="00:02:24.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOPRWL" nation="POL" region="LBS" clubid="2727" name="WOPR Województwa Lubuskiego">
          <CONTACT city="Zielona Góra" email="kifertnat@gmail.com" internet="www.woprlubuski.pl" name="Kifert Natalia" state="LUBUS" street="Lisowskiego 1" zip="65-072" />
          <ATHLETES>
            <ATHLETE birthdate="1975-05-25" firstname="Mieszko" gender="M" lastname="Bencych" nation="POL" athleteid="2728">
              <RESULTS>
                <RESULT eventid="1239" points="330" reactiontime="+89" swimtime="00:02:54.24" resultid="2729" heatid="8978" lane="8" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:20.74" />
                    <SPLIT distance="150" swimtime="00:02:06.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="359" reactiontime="+89" swimtime="00:01:18.19" resultid="2730" heatid="9051" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="358" reactiontime="+88" swimtime="00:00:35.53" resultid="2731" heatid="9167" lane="6" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-02" firstname="Natalia" gender="F" lastname="Kifert" nation="POL" athleteid="2739">
              <RESULTS>
                <RESULT eventid="1187" points="309" reactiontime="+66" swimtime="00:00:37.94" resultid="2740" heatid="8951" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1457" points="299" reactiontime="+66" swimtime="00:01:22.24" resultid="2741" heatid="9077" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="2742" heatid="9140" lane="5" entrytime="00:02:55.00" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="2743" heatid="9155" lane="7" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-20" firstname="Kalina" gender="F" lastname="Chęcińska" nation="POL" athleteid="2732">
              <RESULTS>
                <RESULT eventid="1062" points="376" reactiontime="+85" swimtime="00:00:32.18" resultid="2733" heatid="8890" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1096" points="298" reactiontime="+91" swimtime="00:03:02.39" resultid="2734" heatid="8918" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:26.58" />
                    <SPLIT distance="150" swimtime="00:02:20.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="330" reactiontime="+91" swimtime="00:01:21.99" resultid="2735" heatid="9004" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="274" reactiontime="+87" swimtime="00:00:37.52" resultid="2736" heatid="9056" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1555" points="278" reactiontime="+94" swimtime="00:06:38.09" resultid="2737" heatid="9114" lane="8" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                    <SPLIT distance="100" swimtime="00:01:35.19" />
                    <SPLIT distance="150" swimtime="00:02:27.36" />
                    <SPLIT distance="200" swimtime="00:03:18.57" />
                    <SPLIT distance="250" swimtime="00:04:14.18" />
                    <SPLIT distance="300" swimtime="00:05:09.29" />
                    <SPLIT distance="350" swimtime="00:05:55.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="235" reactiontime="+92" swimtime="00:01:28.39" resultid="2738" heatid="9125" lane="0" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-12-07" firstname="Wojciech" gender="M" lastname="Oczkoś" nation="POL" athleteid="2744">
              <RESULTS>
                <RESULT eventid="1079" points="345" reactiontime="+84" swimtime="00:00:28.88" resultid="2745" heatid="8908" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1165" points="189" reactiontime="+90" swimtime="00:24:40.96" resultid="2746" heatid="8944" lane="3" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                    <SPLIT distance="100" swimtime="00:01:20.37" />
                    <SPLIT distance="150" swimtime="00:02:05.52" />
                    <SPLIT distance="200" swimtime="00:02:52.33" />
                    <SPLIT distance="250" swimtime="00:03:40.39" />
                    <SPLIT distance="300" swimtime="00:04:28.71" />
                    <SPLIT distance="350" swimtime="00:05:17.87" />
                    <SPLIT distance="400" swimtime="00:06:06.82" />
                    <SPLIT distance="450" swimtime="00:06:56.55" />
                    <SPLIT distance="500" swimtime="00:07:46.82" />
                    <SPLIT distance="550" swimtime="00:08:36.81" />
                    <SPLIT distance="600" swimtime="00:09:26.37" />
                    <SPLIT distance="650" swimtime="00:10:16.84" />
                    <SPLIT distance="700" swimtime="00:11:06.96" />
                    <SPLIT distance="750" swimtime="00:11:56.52" />
                    <SPLIT distance="800" swimtime="00:12:46.51" />
                    <SPLIT distance="850" swimtime="00:13:37.25" />
                    <SPLIT distance="900" swimtime="00:14:27.90" />
                    <SPLIT distance="950" swimtime="00:15:18.82" />
                    <SPLIT distance="1000" swimtime="00:16:09.79" />
                    <SPLIT distance="1050" swimtime="00:17:00.56" />
                    <SPLIT distance="1100" swimtime="00:17:51.71" />
                    <SPLIT distance="1150" swimtime="00:18:42.55" />
                    <SPLIT distance="1200" swimtime="00:19:33.88" />
                    <SPLIT distance="1250" swimtime="00:20:25.47" />
                    <SPLIT distance="1300" swimtime="00:21:16.88" />
                    <SPLIT distance="1350" swimtime="00:22:08.00" />
                    <SPLIT distance="1400" swimtime="00:22:59.62" />
                    <SPLIT distance="1450" swimtime="00:23:51.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="322" reactiontime="+83" swimtime="00:01:05.52" resultid="2747" heatid="8993" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="325" reactiontime="+87" swimtime="00:01:13.64" resultid="2748" heatid="9015" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="267" reactiontime="+92" swimtime="00:01:26.29" resultid="2749" heatid="9045" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="297" reactiontime="+87" swimtime="00:00:32.64" resultid="2750" heatid="9069" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1681" points="288" reactiontime="+93" swimtime="00:00:38.21" resultid="2751" heatid="9167" lane="1" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="293" reactiontime="+89" swimtime="00:02:04.25" resultid="2752" heatid="8934" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:01.41" />
                    <SPLIT distance="150" swimtime="00:01:36.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2732" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="2728" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2739" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2744" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="283" reactiontime="+68" swimtime="00:02:17.73" resultid="2753" heatid="9175" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:13.31" />
                    <SPLIT distance="150" swimtime="00:01:45.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2739" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2744" number="2" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2728" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2732" number="4" reactiontime="+5" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="LUB" nation="POL" region="LBS" clubid="4975" name="ZKS Jorge Drzonków">
          <CONTACT city="Świdnica" email="horbacz.marcin@wp.pl" name="Horbacz" phone="603672717" state="LUB" street="Buchałów 12c" zip="66-008" />
          <ATHLETES>
            <ATHLETE birthdate="1971-05-11" firstname="Grzegorz" gender="M" lastname="Sądel" nation="POL" athleteid="4976">
              <RESULTS>
                <RESULT eventid="1165" points="294" reactiontime="+96" swimtime="00:21:17.42" resultid="4977" heatid="8946" lane="3" entrytime="00:20:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="150" swimtime="00:01:55.24" />
                    <SPLIT distance="200" swimtime="00:02:36.20" />
                    <SPLIT distance="250" swimtime="00:03:17.60" />
                    <SPLIT distance="300" swimtime="00:03:59.22" />
                    <SPLIT distance="350" swimtime="00:04:41.68" />
                    <SPLIT distance="400" swimtime="00:05:24.21" />
                    <SPLIT distance="450" swimtime="00:06:06.87" />
                    <SPLIT distance="500" swimtime="00:06:50.01" />
                    <SPLIT distance="550" swimtime="00:07:32.51" />
                    <SPLIT distance="600" swimtime="00:08:15.92" />
                    <SPLIT distance="650" swimtime="00:08:58.40" />
                    <SPLIT distance="700" swimtime="00:09:42.08" />
                    <SPLIT distance="750" swimtime="00:10:25.11" />
                    <SPLIT distance="800" swimtime="00:11:08.49" />
                    <SPLIT distance="850" swimtime="00:11:51.92" />
                    <SPLIT distance="900" swimtime="00:12:35.20" />
                    <SPLIT distance="950" swimtime="00:13:18.97" />
                    <SPLIT distance="1000" swimtime="00:14:03.20" />
                    <SPLIT distance="1050" swimtime="00:14:46.65" />
                    <SPLIT distance="1100" swimtime="00:15:30.52" />
                    <SPLIT distance="1150" swimtime="00:16:14.15" />
                    <SPLIT distance="1200" swimtime="00:16:57.82" />
                    <SPLIT distance="1250" swimtime="00:17:41.33" />
                    <SPLIT distance="1300" swimtime="00:18:24.76" />
                    <SPLIT distance="1350" swimtime="00:19:08.65" />
                    <SPLIT distance="1400" swimtime="00:19:52.31" />
                    <SPLIT distance="1450" swimtime="00:20:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="4978" heatid="9029" lane="2" entrytime="00:02:44.00" entrycourse="SCM" />
                <RESULT eventid="1578" points="267" reactiontime="+90" swimtime="00:06:05.71" resultid="4979" heatid="9121" lane="9" entrytime="00:05:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="150" swimtime="00:02:09.35" />
                    <SPLIT distance="200" swimtime="00:02:59.34" />
                    <SPLIT distance="250" swimtime="00:03:51.82" />
                    <SPLIT distance="300" swimtime="00:04:43.93" />
                    <SPLIT distance="350" swimtime="00:05:24.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="282" reactiontime="+93" swimtime="00:01:13.85" resultid="4980" heatid="9134" lane="9" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="4981" heatid="9190" lane="8" entrytime="00:04:59.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SLO" clubid="3400" name="Športový plavecký klub Kúpele Piešťany - KUPI" shortname="Športový plavecký klub Kúpele ">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1986-01-15" firstname="Lucia" gender="F" lastname="Vachanová" nation="SLO" athleteid="3414">
              <RESULTS>
                <RESULT eventid="1187" points="389" reactiontime="+75" swimtime="00:00:35.16" resultid="3415" heatid="8952" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1256" points="469" reactiontime="+90" swimtime="00:01:05.64" resultid="3416" heatid="8983" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="406" reactiontime="+83" swimtime="00:01:14.28" resultid="3417" heatid="9077" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="442" reactiontime="+88" swimtime="00:02:25.40" resultid="3418" heatid="9093" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:10.89" />
                    <SPLIT distance="150" swimtime="00:01:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="401" reactiontime="+76" swimtime="00:02:41.58" resultid="3419" heatid="9141" lane="9" entrytime="00:02:49.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:20.00" />
                    <SPLIT distance="150" swimtime="00:02:01.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="422" reactiontime="+98" swimtime="00:05:12.63" resultid="3420" heatid="9181" lane="0" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:13.90" />
                    <SPLIT distance="150" swimtime="00:01:53.40" />
                    <SPLIT distance="200" swimtime="00:02:33.29" />
                    <SPLIT distance="250" swimtime="00:03:13.28" />
                    <SPLIT distance="300" swimtime="00:03:54.00" />
                    <SPLIT distance="350" swimtime="00:04:34.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-04-20" firstname="Anna" gender="F" lastname="Kičínová" nation="SLO" athleteid="3401">
              <RESULTS>
                <RESULT eventid="1222" points="283" reactiontime="+100" swimtime="00:03:24.94" resultid="3402" heatid="8969" lane="3" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                    <SPLIT distance="100" swimtime="00:01:38.39" />
                    <SPLIT distance="150" swimtime="00:02:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="229" reactiontime="+104" swimtime="00:03:15.32" resultid="3403" heatid="9024" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:30.53" />
                    <SPLIT distance="150" swimtime="00:02:21.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="274" reactiontime="+98" swimtime="00:01:36.01" resultid="3404" heatid="9040" lane="1" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="237" reactiontime="+85" swimtime="00:00:39.38" resultid="3405" heatid="9056" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1595" points="247" reactiontime="+93" swimtime="00:01:27.03" resultid="3406" heatid="9125" lane="4" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="274" reactiontime="+96" swimtime="00:00:44.34" resultid="3407" heatid="9155" lane="5" entrytime="00:00:44.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-04-03" firstname="Juraj" gender="M" lastname="Horil" nation="SLO" athleteid="3421">
              <RESULTS>
                <RESULT eventid="1239" points="276" reactiontime="+88" swimtime="00:03:04.86" resultid="3422" heatid="8976" lane="9" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:01:24.87" />
                    <SPLIT distance="150" swimtime="00:02:14.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="269" reactiontime="+82" swimtime="00:01:18.46" resultid="3423" heatid="9013" lane="4" entrytime="00:01:19.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="316" reactiontime="+88" swimtime="00:01:21.58" resultid="3424" heatid="9050" lane="1" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="206" reactiontime="+93" swimtime="00:00:36.89" resultid="3425" heatid="9064" lane="1" entrytime="00:00:35.20" />
                <RESULT eventid="1681" points="328" reactiontime="+82" swimtime="00:00:36.58" resultid="3426" heatid="9168" lane="3" entrytime="00:00:36.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-10-27" firstname="Pavol" gender="M" lastname="Škodný" nation="SLO" athleteid="3408">
              <RESULTS>
                <RESULT eventid="1341" points="273" reactiontime="+108" swimtime="00:02:47.18" resultid="3409" heatid="9029" lane="0" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:18.29" />
                    <SPLIT distance="150" swimtime="00:02:02.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="331" reactiontime="+64" swimtime="00:01:10.72" resultid="3410" heatid="9084" lane="5" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="337" reactiontime="+100" swimtime="00:05:38.30" resultid="3411" heatid="9121" lane="2" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:02:00.01" />
                    <SPLIT distance="200" swimtime="00:02:42.84" />
                    <SPLIT distance="250" swimtime="00:03:33.44" />
                    <SPLIT distance="300" swimtime="00:04:23.74" />
                    <SPLIT distance="350" swimtime="00:05:03.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="319" reactiontime="+97" swimtime="00:01:10.84" resultid="3412" heatid="9133" lane="3" entrytime="00:01:13.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="310" reactiontime="+75" swimtime="00:02:36.70" resultid="3413" heatid="9148" lane="5" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:15.35" />
                    <SPLIT distance="150" swimtime="00:01:56.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1698" points="280" reactiontime="+88" swimtime="00:02:18.19" resultid="3427" heatid="9175" lane="0" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:11.45" />
                    <SPLIT distance="150" swimtime="00:01:51.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3414" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3421" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="3401" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3408" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

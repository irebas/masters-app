<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="KS Warszawianka" version="11.69132">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Łódź" name="Otwarte Letnie Mistrzostwa Okręgu Łódzkiego 2021 oraz Letnie Mistrzostwa Masters" course="LCM" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2021-05-30" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Łódź" nation="POL" />
      <POINTTABLE pointtableid="3014" name="FINA Point Scoring" version="2021" />
      <QUALIFY from="2020-01-01" until="2021-05-28" />
      <SESSIONS>
        <SESSION date="2021-05-29" daytime="13:45" endtime="17:55" name="I Blok" number="1" warmupfrom="13:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="13:45" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3864" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3865" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2260" />
                    <RANKING order="2" place="2" resultid="3112" />
                    <RANKING order="3" place="3" resultid="3486" />
                    <RANKING order="4" place="4" resultid="3119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3866" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3106" />
                    <RANKING order="2" place="2" resultid="3589" />
                    <RANKING order="3" place="3" resultid="3592" />
                    <RANKING order="4" place="4" resultid="3480" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4011" daytime="13:45" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1065" daytime="13:52" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3861" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3138" />
                    <RANKING order="2" place="2" resultid="3597" />
                    <RANKING order="3" place="3" resultid="3145" />
                    <RANKING order="4" place="4" resultid="3152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3862" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2268" />
                    <RANKING order="2" place="2" resultid="3126" />
                    <RANKING order="3" place="3" resultid="2277" />
                    <RANKING order="4" place="4" resultid="2284" />
                    <RANKING order="5" place="5" resultid="3326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3863" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3320" />
                    <RANKING order="2" place="2" resultid="3133" />
                    <RANKING order="3" place="3" resultid="2419" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4012" daytime="13:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4013" daytime="13:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1070" daytime="14:04" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1071" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3607" />
                    <RANKING order="2" place="2" resultid="2038" />
                    <RANKING order="3" place="3" resultid="2888" />
                    <RANKING order="4" place="4" resultid="2127" />
                    <RANKING order="5" place="5" resultid="2223" />
                    <RANKING order="6" place="6" resultid="3614" />
                    <RANKING order="7" place="7" resultid="3492" />
                    <RANKING order="8" place="8" resultid="3497" />
                    <RANKING order="9" place="9" resultid="2046" />
                    <RANKING order="10" place="10" resultid="2905" />
                    <RANKING order="11" place="11" resultid="2900" />
                    <RANKING order="12" place="12" resultid="2440" />
                    <RANKING order="13" place="13" resultid="3158" />
                    <RANKING order="14" place="14" resultid="2229" />
                    <RANKING order="15" place="15" resultid="3503" />
                    <RANKING order="16" place="16" resultid="2675" />
                    <RANKING order="17" place="-1" resultid="2445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3388" />
                    <RANKING order="2" place="2" resultid="3508" />
                    <RANKING order="3" place="3" resultid="2117" />
                    <RANKING order="4" place="4" resultid="2829" />
                    <RANKING order="5" place="5" resultid="2122" />
                    <RANKING order="6" place="6" resultid="3350" />
                    <RANKING order="7" place="7" resultid="3602" />
                    <RANKING order="8" place="8" resultid="2431" />
                    <RANKING order="9" place="9" resultid="3382" />
                    <RANKING order="10" place="10" resultid="2051" />
                    <RANKING order="11" place="11" resultid="2218" />
                    <RANKING order="12" place="12" resultid="3356" />
                    <RANKING order="13" place="13" resultid="2057" />
                    <RANKING order="14" place="14" resultid="2848" />
                    <RANKING order="15" place="15" resultid="2234" />
                    <RANKING order="16" place="16" resultid="2133" />
                    <RANKING order="17" place="17" resultid="2042" />
                    <RANKING order="18" place="18" resultid="2664" />
                    <RANKING order="19" place="19" resultid="3376" />
                    <RANKING order="20" place="20" resultid="3365" />
                    <RANKING order="21" place="21" resultid="3534" />
                    <RANKING order="22" place="22" resultid="2645" />
                    <RANKING order="23" place="23" resultid="2237" />
                    <RANKING order="24" place="24" resultid="2661" />
                    <RANKING order="25" place="25" resultid="2894" />
                    <RANKING order="26" place="26" resultid="2651" />
                    <RANKING order="27" place="27" resultid="2656" />
                    <RANKING order="28" place="28" resultid="3371" />
                    <RANKING order="29" place="29" resultid="2307" />
                    <RANKING order="30" place="-1" resultid="2436" />
                    <RANKING order="31" place="-1" resultid="3519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2835" />
                    <RANKING order="2" place="2" resultid="3332" />
                    <RANKING order="3" place="3" resultid="3514" />
                    <RANKING order="4" place="4" resultid="3338" />
                    <RANKING order="5" place="5" resultid="2297" />
                    <RANKING order="6" place="6" resultid="2878" />
                    <RANKING order="7" place="7" resultid="3163" />
                    <RANKING order="8" place="8" resultid="3056" />
                    <RANKING order="9" place="9" resultid="3344" />
                    <RANKING order="10" place="10" resultid="3171" />
                    <RANKING order="11" place="11" resultid="3524" />
                    <RANKING order="12" place="12" resultid="2842" />
                    <RANKING order="13" place="13" resultid="3529" />
                    <RANKING order="14" place="14" resultid="2304" />
                    <RANKING order="15" place="15" resultid="2883" />
                    <RANKING order="16" place="-1" resultid="3062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3362" />
                    <RANKING order="2" place="2" resultid="2424" />
                    <RANKING order="3" place="3" resultid="2032" />
                    <RANKING order="4" place="4" resultid="2019" />
                    <RANKING order="5" place="5" resultid="2291" />
                    <RANKING order="6" place="6" resultid="2669" />
                    <RANKING order="7" place="7" resultid="3035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2763" />
                    <RANKING order="2" place="2" resultid="2768" />
                    <RANKING order="3" place="3" resultid="2759" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4014" daytime="14:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4015" daytime="14:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4016" daytime="14:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4017" daytime="14:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4018" daytime="14:09" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4019" daytime="14:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4020" daytime="14:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4021" daytime="14:13" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4022" daytime="14:14" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1120" daytime="14:15" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3867" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2472" />
                    <RANKING order="2" place="2" resultid="3213" />
                    <RANKING order="3" place="3" resultid="2146" />
                    <RANKING order="4" place="4" resultid="2867" />
                    <RANKING order="5" place="5" resultid="2932" />
                    <RANKING order="6" place="6" resultid="3189" />
                    <RANKING order="7" place="7" resultid="3553" />
                    <RANKING order="8" place="8" resultid="2353" />
                    <RANKING order="9" place="9" resultid="2329" />
                    <RANKING order="10" place="10" resultid="2854" />
                    <RANKING order="11" place="11" resultid="2686" />
                    <RANKING order="12" place="12" resultid="2719" />
                    <RANKING order="13" place="13" resultid="3178" />
                    <RANKING order="14" place="14" resultid="2478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3868" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2949" />
                    <RANKING order="2" place="2" resultid="2346" />
                    <RANKING order="3" place="3" resultid="3220" />
                    <RANKING order="4" place="4" resultid="2465" />
                    <RANKING order="5" place="5" resultid="2702" />
                    <RANKING order="6" place="6" resultid="2240" />
                    <RANKING order="7" place="7" resultid="2460" />
                    <RANKING order="8" place="8" resultid="2152" />
                    <RANKING order="9" place="9" resultid="3429" />
                    <RANKING order="10" place="10" resultid="3558" />
                    <RANKING order="11" place="11" resultid="2926" />
                    <RANKING order="12" place="12" resultid="2713" />
                    <RANKING order="13" place="13" resultid="2696" />
                    <RANKING order="14" place="14" resultid="3563" />
                    <RANKING order="15" place="15" resultid="3424" />
                    <RANKING order="16" place="16" resultid="2251" />
                    <RANKING order="17" place="17" resultid="2335" />
                    <RANKING order="18" place="18" resultid="2364" />
                    <RANKING order="19" place="19" resultid="3227" />
                    <RANKING order="20" place="20" resultid="2691" />
                    <RANKING order="21" place="21" resultid="2943" />
                    <RANKING order="22" place="22" resultid="2341" />
                    <RANKING order="23" place="23" resultid="2921" />
                    <RANKING order="24" place="24" resultid="2938" />
                    <RANKING order="25" place="25" resultid="2860" />
                    <RANKING order="26" place="26" resultid="2139" />
                    <RANKING order="27" place="27" resultid="2488" />
                    <RANKING order="28" place="28" resultid="3620" />
                    <RANKING order="29" place="29" resultid="2956" />
                    <RANKING order="30" place="30" resultid="3183" />
                    <RANKING order="31" place="31" resultid="2681" />
                    <RANKING order="32" place="32" resultid="2494" />
                    <RANKING order="33" place="33" resultid="2510" />
                    <RANKING order="34" place="34" resultid="2505" />
                    <RANKING order="35" place="35" resultid="2917" />
                    <RANKING order="36" place="36" resultid="2246" />
                    <RANKING order="37" place="37" resultid="2500" />
                    <RANKING order="38" place="38" resultid="2312" />
                    <RANKING order="39" place="-1" resultid="2483" />
                    <RANKING order="40" place="-1" resultid="2063" />
                    <RANKING order="41" place="-1" resultid="2911" />
                    <RANKING order="42" place="-1" resultid="2961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3869" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2377" />
                    <RANKING order="2" place="2" resultid="2369" />
                    <RANKING order="3" place="3" resultid="2450" />
                    <RANKING order="4" place="4" resultid="2360" />
                    <RANKING order="5" place="5" resultid="3394" />
                    <RANKING order="6" place="6" resultid="3406" />
                    <RANKING order="7" place="7" resultid="3418" />
                    <RANKING order="8" place="8" resultid="3856" />
                    <RANKING order="9" place="9" resultid="3400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3870" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3545" />
                    <RANKING order="2" place="2" resultid="3201" />
                    <RANKING order="3" place="3" resultid="2323" />
                    <RANKING order="4" place="4" resultid="3195" />
                    <RANKING order="5" place="5" resultid="3207" />
                    <RANKING order="6" place="6" resultid="2025" />
                    <RANKING order="7" place="7" resultid="3301" />
                    <RANKING order="8" place="8" resultid="2455" />
                    <RANKING order="9" place="9" resultid="3305" />
                    <RANKING order="10" place="10" resultid="3412" />
                    <RANKING order="11" place="11" resultid="2318" />
                    <RANKING order="12" place="12" resultid="3540" />
                    <RANKING order="13" place="12" resultid="3550" />
                    <RANKING order="14" place="14" resultid="2708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3871" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2179" />
                    <RANKING order="2" place="2" resultid="3042" />
                    <RANKING order="3" place="3" resultid="2788" />
                    <RANKING order="4" place="4" resultid="2784" />
                    <RANKING order="5" place="5" resultid="2772" />
                    <RANKING order="6" place="6" resultid="2777" />
                    <RANKING order="7" place="7" resultid="2793" />
                    <RANKING order="8" place="8" resultid="2780" />
                    <RANKING order="9" place="-1" resultid="2005" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4023" daytime="14:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4024" daytime="14:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4025" daytime="14:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4026" daytime="14:19" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4027" daytime="14:21" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4028" daytime="14:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4029" daytime="14:23" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4030" daytime="14:24" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4031" daytime="14:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4032" daytime="14:26" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1143" daytime="14:28" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3872" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2984" />
                    <RANKING order="2" place="2" resultid="2989" />
                    <RANKING order="3" place="3" resultid="2224" />
                    <RANKING order="4" place="4" resultid="2128" />
                    <RANKING order="5" place="5" resultid="3626" />
                    <RANKING order="6" place="6" resultid="2441" />
                    <RANKING order="7" place="7" resultid="3159" />
                    <RANKING order="8" place="8" resultid="2733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3873" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3068" />
                    <RANKING order="2" place="2" resultid="3357" />
                    <RANKING order="3" place="3" resultid="3383" />
                    <RANKING order="4" place="4" resultid="3509" />
                    <RANKING order="5" place="5" resultid="2123" />
                    <RANKING order="6" place="6" resultid="3435" />
                    <RANKING order="7" place="7" resultid="3234" />
                    <RANKING order="8" place="8" resultid="3366" />
                    <RANKING order="9" place="9" resultid="2972" />
                    <RANKING order="10" place="10" resultid="2967" />
                    <RANKING order="11" place="11" resultid="2978" />
                    <RANKING order="12" place="12" resultid="2527" />
                    <RANKING order="13" place="13" resultid="2849" />
                    <RANKING order="14" place="14" resultid="2652" />
                    <RANKING order="15" place="15" resultid="2895" />
                    <RANKING order="16" place="16" resultid="2523" />
                    <RANKING order="17" place="17" resultid="3372" />
                    <RANKING order="18" place="-1" resultid="2437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3874" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3572" />
                    <RANKING order="2" place="2" resultid="2729" />
                    <RANKING order="3" place="3" resultid="3345" />
                    <RANKING order="4" place="4" resultid="2515" />
                    <RANKING order="5" place="5" resultid="2519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3875" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2723" />
                    <RANKING order="2" place="2" resultid="2425" />
                    <RANKING order="3" place="3" resultid="3075" />
                    <RANKING order="4" place="4" resultid="3481" />
                    <RANKING order="5" place="5" resultid="3036" />
                    <RANKING order="6" place="6" resultid="3240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3876" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2796" />
                    <RANKING order="2" place="2" resultid="2769" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4033" daytime="14:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4034" daytime="14:29" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4035" daytime="14:31" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4036" daytime="14:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4037" daytime="14:34" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1166" daytime="14:35" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3877" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2387" />
                    <RANKING order="2" place="2" resultid="3004" />
                    <RANKING order="3" place="3" resultid="2147" />
                    <RANKING order="4" place="4" resultid="2394" />
                    <RANKING order="5" place="5" resultid="2555" />
                    <RANKING order="6" place="6" resultid="3010" />
                    <RANKING order="7" place="7" resultid="2560" />
                    <RANKING order="8" place="8" resultid="2330" />
                    <RANKING order="9" place="9" resultid="2568" />
                    <RANKING order="10" place="10" resultid="2742" />
                    <RANKING order="11" place="11" resultid="2687" />
                    <RANKING order="12" place="12" resultid="2855" />
                    <RANKING order="13" place="-1" resultid="2564" />
                    <RANKING order="14" place="-1" resultid="2720" />
                    <RANKING order="15" place="-1" resultid="3190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3878" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3266" />
                    <RANKING order="2" place="2" resultid="3139" />
                    <RANKING order="3" place="3" resultid="3441" />
                    <RANKING order="4" place="3" resultid="3633" />
                    <RANKING order="5" place="5" resultid="2543" />
                    <RANKING order="6" place="6" resultid="3447" />
                    <RANKING order="7" place="7" resultid="2998" />
                    <RANKING order="8" place="8" resultid="2697" />
                    <RANKING order="9" place="9" resultid="3245" />
                    <RANKING order="10" place="10" resultid="2714" />
                    <RANKING order="11" place="11" resultid="2140" />
                    <RANKING order="12" place="12" resultid="2342" />
                    <RANKING order="13" place="13" resultid="2552" />
                    <RANKING order="14" place="14" resultid="2692" />
                    <RANKING order="15" place="15" resultid="2484" />
                    <RANKING order="16" place="16" resultid="4161" />
                    <RANKING order="17" place="17" resultid="2336" />
                    <RANKING order="18" place="18" resultid="2944" />
                    <RANKING order="19" place="19" resultid="2994" />
                    <RANKING order="20" place="20" resultid="2506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3879" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3251" />
                    <RANKING order="2" place="2" resultid="2537" />
                    <RANKING order="3" place="3" resultid="3407" />
                    <RANKING order="4" place="4" resultid="3079" />
                    <RANKING order="5" place="5" resultid="2285" />
                    <RANKING order="6" place="6" resultid="2547" />
                    <RANKING order="7" place="7" resultid="3261" />
                    <RANKING order="8" place="8" resultid="3858" />
                    <RANKING order="9" place="9" resultid="3419" />
                    <RANKING order="10" place="10" resultid="3327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3880" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3578" />
                    <RANKING order="2" place="2" resultid="2738" />
                    <RANKING order="3" place="3" resultid="2319" />
                    <RANKING order="4" place="4" resultid="3256" />
                    <RANKING order="5" place="5" resultid="2709" />
                    <RANKING order="6" place="6" resultid="2533" />
                    <RANKING order="7" place="-1" resultid="3853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3881" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2010" />
                    <RANKING order="2" place="2" resultid="2800" />
                    <RANKING order="3" place="3" resultid="2781" />
                    <RANKING order="4" place="4" resultid="2111" />
                    <RANKING order="5" place="5" resultid="2069" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4038" daytime="14:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4039" daytime="14:37" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4040" daytime="14:39" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4041" daytime="14:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4042" daytime="14:41" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4043" daytime="14:43" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1189" daytime="14:44" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3882" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3608" />
                    <RANKING order="2" place="2" resultid="3013" />
                    <RANKING order="3" place="3" resultid="2585" />
                    <RANKING order="4" place="4" resultid="3639" />
                    <RANKING order="5" place="5" resultid="3493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3883" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3389" />
                    <RANKING order="2" place="2" resultid="2830" />
                    <RANKING order="3" place="3" resultid="3069" />
                    <RANKING order="4" place="4" resultid="3315" />
                    <RANKING order="5" place="5" resultid="3465" />
                    <RANKING order="6" place="6" resultid="3084" />
                    <RANKING order="7" place="7" resultid="2528" />
                    <RANKING order="8" place="8" resultid="2058" />
                    <RANKING order="9" place="9" resultid="3377" />
                    <RANKING order="10" place="10" resultid="2256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3884" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2261" />
                    <RANKING order="2" place="2" resultid="3453" />
                    <RANKING order="3" place="3" resultid="3113" />
                    <RANKING order="4" place="4" resultid="2879" />
                    <RANKING order="5" place="5" resultid="3459" />
                    <RANKING order="6" place="6" resultid="3057" />
                    <RANKING order="7" place="7" resultid="2579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3885" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2020" />
                    <RANKING order="2" place="2" resultid="2573" />
                    <RANKING order="3" place="3" resultid="2426" />
                    <RANKING order="4" place="4" resultid="2747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3886" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2803" />
                    <RANKING order="2" place="2" resultid="2807" />
                    <RANKING order="3" place="3" resultid="2184" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4044" daytime="14:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4045" daytime="14:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4046" daytime="14:48" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1212" daytime="14:51" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3887" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2868" />
                    <RANKING order="2" place="2" resultid="3658" />
                    <RANKING order="3" place="3" resultid="3276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3888" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2347" />
                    <RANKING order="2" place="2" resultid="2950" />
                    <RANKING order="3" place="3" resultid="3153" />
                    <RANKING order="4" place="4" resultid="2466" />
                    <RANKING order="5" place="5" resultid="2600" />
                    <RANKING order="6" place="6" resultid="2590" />
                    <RANKING order="7" place="7" resultid="3221" />
                    <RANKING order="8" place="8" resultid="3430" />
                    <RANKING order="9" place="9" resultid="2153" />
                    <RANKING order="10" place="10" resultid="3645" />
                    <RANKING order="11" place="11" resultid="3425" />
                    <RANKING order="12" place="12" resultid="3271" />
                    <RANKING order="13" place="13" resultid="3621" />
                    <RANKING order="14" place="14" resultid="3651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3889" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2378" />
                    <RANKING order="2" place="2" resultid="2398" />
                    <RANKING order="3" place="3" resultid="3281" />
                    <RANKING order="4" place="4" resultid="2538" />
                    <RANKING order="5" place="5" resultid="2361" />
                    <RANKING order="6" place="6" resultid="3127" />
                    <RANKING order="7" place="7" resultid="2370" />
                    <RANKING order="8" place="8" resultid="3408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3890" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3090" />
                    <RANKING order="2" place="2" resultid="3413" />
                    <RANKING order="3" place="3" resultid="2456" />
                    <RANKING order="4" place="4" resultid="2595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3891" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2013" />
                    <RANKING order="2" place="2" resultid="2180" />
                    <RANKING order="3" place="-1" resultid="2006" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4047" daytime="14:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4048" daytime="14:53" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4049" daytime="14:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4050" daytime="14:57" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1235" daytime="14:59" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3892" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2039" />
                    <RANKING order="2" place="2" resultid="2612" />
                    <RANKING order="3" place="3" resultid="2889" />
                    <RANKING order="4" place="4" resultid="3615" />
                    <RANKING order="5" place="5" resultid="3014" />
                    <RANKING order="6" place="6" resultid="2047" />
                    <RANKING order="7" place="7" resultid="2906" />
                    <RANKING order="8" place="8" resultid="3627" />
                    <RANKING order="9" place="9" resultid="3680" />
                    <RANKING order="10" place="10" resultid="2230" />
                    <RANKING order="11" place="11" resultid="2676" />
                    <RANKING order="12" place="-1" resultid="2446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3893" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3390" />
                    <RANKING order="2" place="2" resultid="3466" />
                    <RANKING order="3" place="3" resultid="3351" />
                    <RANKING order="4" place="4" resultid="3664" />
                    <RANKING order="5" place="5" resultid="2973" />
                    <RANKING order="6" place="6" resultid="3670" />
                    <RANKING order="7" place="7" resultid="2134" />
                    <RANKING order="8" place="8" resultid="2043" />
                    <RANKING order="9" place="9" resultid="2646" />
                    <RANKING order="10" place="10" resultid="3535" />
                    <RANKING order="11" place="11" resultid="2657" />
                    <RANKING order="12" place="12" resultid="3378" />
                    <RANKING order="13" place="13" resultid="2665" />
                    <RANKING order="14" place="14" resultid="2524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3894" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3333" />
                    <RANKING order="2" place="2" resultid="2298" />
                    <RANKING order="3" place="3" resultid="2836" />
                    <RANKING order="4" place="4" resultid="3473" />
                    <RANKING order="5" place="5" resultid="2606" />
                    <RANKING order="6" place="6" resultid="2843" />
                    <RANKING order="7" place="7" resultid="3063" />
                    <RANKING order="8" place="8" resultid="3675" />
                    <RANKING order="9" place="9" resultid="2884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3895" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3471" />
                    <RANKING order="2" place="2" resultid="2292" />
                    <RANKING order="3" place="3" resultid="2574" />
                    <RANKING order="4" place="4" resultid="3363" />
                    <RANKING order="5" place="5" resultid="2033" />
                    <RANKING order="6" place="6" resultid="2670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3896" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2189" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4051" daytime="14:59" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4052" daytime="15:01" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4053" daytime="15:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4054" daytime="15:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4055" daytime="15:05" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1258" daytime="15:07" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3897" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3214" />
                    <RANKING order="2" place="2" resultid="2388" />
                    <RANKING order="3" place="3" resultid="3005" />
                    <RANKING order="4" place="4" resultid="2933" />
                    <RANKING order="5" place="5" resultid="3019" />
                    <RANKING order="6" place="6" resultid="3659" />
                    <RANKING order="7" place="7" resultid="2354" />
                    <RANKING order="8" place="8" resultid="2856" />
                    <RANKING order="9" place="9" resultid="2721" />
                    <RANKING order="10" place="-1" resultid="2331" />
                    <RANKING order="11" place="-1" resultid="2565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3898" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2467" />
                    <RANKING order="2" place="2" resultid="3431" />
                    <RANKING order="3" place="3" resultid="2591" />
                    <RANKING order="4" place="4" resultid="2241" />
                    <RANKING order="5" place="5" resultid="2703" />
                    <RANKING order="6" place="6" resultid="3564" />
                    <RANKING order="7" place="7" resultid="2927" />
                    <RANKING order="8" place="8" resultid="3228" />
                    <RANKING order="9" place="9" resultid="2999" />
                    <RANKING order="10" place="10" resultid="2252" />
                    <RANKING order="11" place="11" resultid="2365" />
                    <RANKING order="12" place="12" resultid="3652" />
                    <RANKING order="13" place="13" resultid="2489" />
                    <RANKING order="14" place="14" resultid="3184" />
                    <RANKING order="15" place="15" resultid="2957" />
                    <RANKING order="16" place="16" resultid="3685" />
                    <RANKING order="17" place="17" resultid="2501" />
                    <RANKING order="18" place="18" resultid="2313" />
                    <RANKING order="19" place="19" resultid="2247" />
                    <RANKING order="20" place="-1" resultid="2912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3899" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3287" />
                    <RANKING order="2" place="2" resultid="2269" />
                    <RANKING order="3" place="3" resultid="2617" />
                    <RANKING order="4" place="4" resultid="3395" />
                    <RANKING order="5" place="5" resultid="2371" />
                    <RANKING order="6" place="6" resultid="3328" />
                    <RANKING order="7" place="-1" resultid="3583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3900" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3541" />
                    <RANKING order="2" place="2" resultid="2324" />
                    <RANKING order="3" place="3" resultid="2026" />
                    <RANKING order="4" place="4" resultid="2406" />
                    <RANKING order="5" place="5" resultid="3306" />
                    <RANKING order="6" place="6" resultid="2710" />
                    <RANKING order="7" place="-1" resultid="3302" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3901" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2789" />
                    <RANKING order="2" place="2" resultid="2812" />
                    <RANKING order="3" place="3" resultid="2070" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4056" daytime="15:07" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4057" daytime="15:09" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4058" daytime="15:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4059" daytime="15:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4060" daytime="15:13" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1281" daytime="15:15" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3902" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3609" />
                    <RANKING order="2" place="2" resultid="2586" />
                    <RANKING order="3" place="3" resultid="3640" />
                    <RANKING order="4" place="4" resultid="3498" />
                    <RANKING order="5" place="5" resultid="2907" />
                    <RANKING order="6" place="6" resultid="3681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3903" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2432" />
                    <RANKING order="2" place="2" resultid="3391" />
                    <RANKING order="3" place="3" resultid="3085" />
                    <RANKING order="4" place="4" resultid="3316" />
                    <RANKING order="5" place="5" resultid="3467" />
                    <RANKING order="6" place="6" resultid="3603" />
                    <RANKING order="7" place="7" resultid="3384" />
                    <RANKING order="8" place="8" resultid="2052" />
                    <RANKING order="9" place="9" resultid="3436" />
                    <RANKING order="10" place="10" resultid="2979" />
                    <RANKING order="11" place="11" resultid="3665" />
                    <RANKING order="12" place="12" resultid="3671" />
                    <RANKING order="13" place="13" resultid="3379" />
                    <RANKING order="14" place="14" resultid="2647" />
                    <RANKING order="15" place="15" resultid="3536" />
                    <RANKING order="16" place="16" resultid="3367" />
                    <RANKING order="17" place="-1" resultid="3520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3904" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2262" />
                    <RANKING order="2" place="2" resultid="3164" />
                    <RANKING order="3" place="3" resultid="3339" />
                    <RANKING order="4" place="4" resultid="3120" />
                    <RANKING order="5" place="5" resultid="3487" />
                    <RANKING order="6" place="6" resultid="2837" />
                    <RANKING order="7" place="7" resultid="3058" />
                    <RANKING order="8" place="8" resultid="3172" />
                    <RANKING order="9" place="9" resultid="3064" />
                    <RANKING order="10" place="10" resultid="3474" />
                    <RANKING order="11" place="11" resultid="3460" />
                    <RANKING order="12" place="12" resultid="2607" />
                    <RANKING order="13" place="13" resultid="3525" />
                    <RANKING order="14" place="14" resultid="3346" />
                    <RANKING order="15" place="15" resultid="2520" />
                    <RANKING order="16" place="16" resultid="3530" />
                    <RANKING order="17" place="17" resultid="2580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3905" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2427" />
                    <RANKING order="2" place="2" resultid="2623" />
                    <RANKING order="3" place="3" resultid="2671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3906" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2185" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4061" daytime="15:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4062" daytime="15:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4063" daytime="15:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4064" daytime="15:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4065" daytime="15:28" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1304" daytime="15:32" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3907" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3277" />
                    <RANKING order="2" place="2" resultid="2473" />
                    <RANKING order="3" place="3" resultid="3215" />
                    <RANKING order="4" place="4" resultid="3554" />
                    <RANKING order="5" place="5" resultid="2355" />
                    <RANKING order="6" place="6" resultid="3179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3908" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2348" />
                    <RANKING order="2" place="2" resultid="3222" />
                    <RANKING order="3" place="3" resultid="2951" />
                    <RANKING order="4" place="4" resultid="3146" />
                    <RANKING order="5" place="5" resultid="2461" />
                    <RANKING order="6" place="6" resultid="3559" />
                    <RANKING order="7" place="7" resultid="2601" />
                    <RANKING order="8" place="8" resultid="3442" />
                    <RANKING order="9" place="9" resultid="3154" />
                    <RANKING order="10" place="10" resultid="3432" />
                    <RANKING order="11" place="11" resultid="3229" />
                    <RANKING order="12" place="12" resultid="3565" />
                    <RANKING order="13" place="13" resultid="2628" />
                    <RANKING order="14" place="14" resultid="2366" />
                    <RANKING order="15" place="15" resultid="3426" />
                    <RANKING order="16" place="16" resultid="3448" />
                    <RANKING order="17" place="17" resultid="3622" />
                    <RANKING order="18" place="18" resultid="2861" />
                    <RANKING order="19" place="19" resultid="2939" />
                    <RANKING order="20" place="20" resultid="3686" />
                    <RANKING order="21" place="21" resultid="2495" />
                    <RANKING order="22" place="22" resultid="3185" />
                    <RANKING order="23" place="-1" resultid="2064" />
                    <RANKING order="24" place="-1" resultid="2913" />
                    <RANKING order="25" place="-1" resultid="2962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3909" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2379" />
                    <RANKING order="2" place="2" resultid="2399" />
                    <RANKING order="3" place="3" resultid="2451" />
                    <RANKING order="4" place="4" resultid="3288" />
                    <RANKING order="5" place="5" resultid="2278" />
                    <RANKING order="6" place="6" resultid="2548" />
                    <RANKING order="7" place="7" resultid="2372" />
                    <RANKING order="8" place="8" resultid="3329" />
                    <RANKING order="9" place="9" resultid="2618" />
                    <RANKING order="10" place="10" resultid="3420" />
                    <RANKING order="11" place="11" resultid="3401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3910" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3202" />
                    <RANKING order="2" place="2" resultid="3208" />
                    <RANKING order="3" place="3" resultid="2420" />
                    <RANKING order="4" place="4" resultid="3321" />
                    <RANKING order="5" place="5" resultid="3093" />
                    <RANKING order="6" place="6" resultid="2410" />
                    <RANKING order="7" place="7" resultid="2633" />
                    <RANKING order="8" place="8" resultid="3551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3911" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3043" />
                    <RANKING order="2" place="2" resultid="3697" />
                    <RANKING order="3" place="3" resultid="2825" />
                    <RANKING order="4" place="4" resultid="2813" />
                    <RANKING order="5" place="5" resultid="2773" />
                    <RANKING order="6" place="6" resultid="2820" />
                    <RANKING order="7" place="7" resultid="2817" />
                    <RANKING order="8" place="-1" resultid="2794" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4066" daytime="15:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4067" daytime="15:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4068" daytime="15:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4069" daytime="15:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4070" daytime="15:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4071" daytime="15:51" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4072" daytime="15:54" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1327" daytime="15:57" gender="F" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3912" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2985" />
                    <RANKING order="2" place="2" resultid="2990" />
                    <RANKING order="3" place="3" resultid="2129" />
                    <RANKING order="4" place="4" resultid="3628" />
                    <RANKING order="5" place="5" resultid="2901" />
                    <RANKING order="6" place="6" resultid="2734" />
                    <RANKING order="7" place="7" resultid="3504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3913" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3070" />
                    <RANKING order="2" place="2" resultid="3358" />
                    <RANKING order="3" place="3" resultid="3385" />
                    <RANKING order="4" place="4" resultid="3510" />
                    <RANKING order="5" place="5" resultid="2118" />
                    <RANKING order="6" place="6" resultid="3437" />
                    <RANKING order="7" place="7" resultid="2968" />
                    <RANKING order="8" place="8" resultid="2974" />
                    <RANKING order="9" place="9" resultid="3235" />
                    <RANKING order="10" place="10" resultid="2980" />
                    <RANKING order="11" place="11" resultid="3368" />
                    <RANKING order="12" place="12" resultid="2235" />
                    <RANKING order="13" place="13" resultid="2896" />
                    <RANKING order="14" place="14" resultid="2238" />
                    <RANKING order="15" place="15" resultid="3373" />
                    <RANKING order="16" place="16" resultid="2308" />
                    <RANKING order="17" place="17" resultid="2525" />
                    <RANKING order="18" place="-1" resultid="2438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3914" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2263" />
                    <RANKING order="2" place="2" resultid="3573" />
                    <RANKING order="3" place="3" resultid="2730" />
                    <RANKING order="4" place="4" resultid="3454" />
                    <RANKING order="5" place="5" resultid="2516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3915" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2724" />
                    <RANKING order="2" place="2" resultid="3076" />
                    <RANKING order="3" place="3" resultid="3482" />
                    <RANKING order="4" place="4" resultid="3241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3916" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2797" />
                    <RANKING order="2" place="2" resultid="2760" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4073" daytime="15:57" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4074" daytime="16:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4075" daytime="16:03" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4076" daytime="16:05" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1350" daytime="16:07" gender="M" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3917" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2389" />
                    <RANKING order="2" place="2" resultid="3006" />
                    <RANKING order="3" place="3" resultid="3660" />
                    <RANKING order="4" place="4" resultid="2556" />
                    <RANKING order="5" place="5" resultid="2395" />
                    <RANKING order="6" place="6" resultid="2332" />
                    <RANKING order="7" place="7" resultid="2561" />
                    <RANKING order="8" place="8" resultid="2569" />
                    <RANKING order="9" place="9" resultid="2743" />
                    <RANKING order="10" place="-1" resultid="3011" />
                    <RANKING order="11" place="-1" resultid="2566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3918" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3140" />
                    <RANKING order="2" place="2" resultid="3267" />
                    <RANKING order="3" place="3" resultid="3443" />
                    <RANKING order="4" place="4" resultid="3634" />
                    <RANKING order="5" place="5" resultid="3246" />
                    <RANKING order="6" place="6" resultid="3449" />
                    <RANKING order="7" place="7" resultid="2544" />
                    <RANKING order="8" place="8" resultid="3000" />
                    <RANKING order="9" place="9" resultid="2715" />
                    <RANKING order="10" place="10" resultid="3646" />
                    <RANKING order="11" place="11" resultid="2343" />
                    <RANKING order="12" place="12" resultid="2922" />
                    <RANKING order="13" place="13" resultid="2553" />
                    <RANKING order="14" place="14" resultid="3272" />
                    <RANKING order="15" place="15" resultid="2485" />
                    <RANKING order="16" place="16" resultid="2337" />
                    <RANKING order="17" place="17" resultid="2995" />
                    <RANKING order="18" place="18" resultid="2918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3919" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3252" />
                    <RANKING order="2" place="2" resultid="2270" />
                    <RANKING order="3" place="3" resultid="2539" />
                    <RANKING order="4" place="4" resultid="3080" />
                    <RANKING order="5" place="5" resultid="3409" />
                    <RANKING order="6" place="6" resultid="2286" />
                    <RANKING order="7" place="7" resultid="3262" />
                    <RANKING order="8" place="8" resultid="3421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3920" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3579" />
                    <RANKING order="2" place="2" resultid="3307" />
                    <RANKING order="3" place="3" resultid="2739" />
                    <RANKING order="4" place="4" resultid="3257" />
                    <RANKING order="5" place="5" resultid="2534" />
                    <RANKING order="6" place="-1" resultid="3854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3921" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2011" />
                    <RANKING order="2" place="2" resultid="2785" />
                    <RANKING order="3" place="3" resultid="2801" />
                    <RANKING order="4" place="4" resultid="2782" />
                    <RANKING order="5" place="5" resultid="2112" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4077" daytime="16:07" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4078" daytime="16:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4079" daytime="16:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4080" daytime="16:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4081" daytime="16:17" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1373" daytime="16:19" gender="F" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3922" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2040" />
                    <RANKING order="2" place="2" resultid="3610" />
                    <RANKING order="3" place="3" resultid="2890" />
                    <RANKING order="4" place="4" resultid="2130" />
                    <RANKING order="5" place="5" resultid="3015" />
                    <RANKING order="6" place="6" resultid="3616" />
                    <RANKING order="7" place="7" resultid="2613" />
                    <RANKING order="8" place="8" resultid="3494" />
                    <RANKING order="9" place="9" resultid="2225" />
                    <RANKING order="10" place="10" resultid="3499" />
                    <RANKING order="11" place="11" resultid="3641" />
                    <RANKING order="12" place="12" resultid="2048" />
                    <RANKING order="13" place="-1" resultid="2677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3923" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3392" />
                    <RANKING order="2" place="2" resultid="2831" />
                    <RANKING order="3" place="3" resultid="3071" />
                    <RANKING order="4" place="4" resultid="3086" />
                    <RANKING order="5" place="5" resultid="3386" />
                    <RANKING order="6" place="6" resultid="2969" />
                    <RANKING order="7" place="7" resultid="2850" />
                    <RANKING order="8" place="8" resultid="2529" />
                    <RANKING order="9" place="9" resultid="2059" />
                    <RANKING order="10" place="10" resultid="3236" />
                    <RANKING order="11" place="11" resultid="2053" />
                    <RANKING order="12" place="12" resultid="3666" />
                    <RANKING order="13" place="13" resultid="2135" />
                    <RANKING order="14" place="14" resultid="2219" />
                    <RANKING order="15" place="15" resultid="2044" />
                    <RANKING order="16" place="16" resultid="3369" />
                    <RANKING order="17" place="17" resultid="3380" />
                    <RANKING order="18" place="18" resultid="2666" />
                    <RANKING order="19" place="19" resultid="2662" />
                    <RANKING order="20" place="20" resultid="2257" />
                    <RANKING order="21" place="21" resultid="3374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3924" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3515" />
                    <RANKING order="2" place="2" resultid="3455" />
                    <RANKING order="3" place="3" resultid="3114" />
                    <RANKING order="4" place="4" resultid="2880" />
                    <RANKING order="5" place="5" resultid="3121" />
                    <RANKING order="6" place="6" resultid="2299" />
                    <RANKING order="7" place="7" resultid="3475" />
                    <RANKING order="8" place="8" resultid="2844" />
                    <RANKING order="9" place="9" resultid="2608" />
                    <RANKING order="10" place="10" resultid="3676" />
                    <RANKING order="11" place="11" resultid="3347" />
                    <RANKING order="12" place="12" resultid="2581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3925" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2021" />
                    <RANKING order="2" place="2" resultid="2293" />
                    <RANKING order="3" place="3" resultid="3077" />
                    <RANKING order="4" place="4" resultid="2725" />
                    <RANKING order="5" place="5" resultid="2748" />
                    <RANKING order="6" place="6" resultid="2034" />
                    <RANKING order="7" place="7" resultid="2575" />
                    <RANKING order="8" place="8" resultid="3483" />
                    <RANKING order="9" place="9" resultid="2624" />
                    <RANKING order="10" place="10" resultid="3037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3926" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2804" />
                    <RANKING order="2" place="2" resultid="2764" />
                    <RANKING order="3" place="3" resultid="2808" />
                    <RANKING order="4" place="4" resultid="2190" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4082" daytime="16:19" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4083" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4084" daytime="16:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4085" daytime="16:23" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4086" daytime="16:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4087" daytime="16:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4088" daytime="16:27" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1396" daytime="16:29" gender="M" number="16" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3927" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2474" />
                    <RANKING order="2" place="2" resultid="2869" />
                    <RANKING order="3" place="3" resultid="3661" />
                    <RANKING order="4" place="4" resultid="3191" />
                    <RANKING order="5" place="5" resultid="2148" />
                    <RANKING order="6" place="6" resultid="3020" />
                    <RANKING order="7" place="-1" resultid="2479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3928" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2349" />
                    <RANKING order="2" place="2" resultid="2952" />
                    <RANKING order="3" place="3" resultid="2602" />
                    <RANKING order="4" place="4" resultid="2704" />
                    <RANKING order="5" place="5" resultid="3433" />
                    <RANKING order="6" place="6" resultid="2154" />
                    <RANKING order="7" place="7" resultid="3635" />
                    <RANKING order="8" place="8" resultid="3223" />
                    <RANKING order="9" place="9" resultid="3427" />
                    <RANKING order="10" place="10" resultid="2698" />
                    <RANKING order="11" place="11" resultid="2928" />
                    <RANKING order="12" place="12" resultid="3647" />
                    <RANKING order="13" place="13" resultid="2693" />
                    <RANKING order="14" place="14" resultid="2338" />
                    <RANKING order="15" place="15" resultid="2141" />
                    <RANKING order="16" place="16" resultid="2496" />
                    <RANKING order="17" place="17" resultid="2945" />
                    <RANKING order="18" place="18" resultid="2511" />
                    <RANKING order="19" place="19" resultid="2862" />
                    <RANKING order="20" place="20" resultid="2490" />
                    <RANKING order="21" place="21" resultid="3653" />
                    <RANKING order="22" place="22" resultid="2682" />
                    <RANKING order="23" place="23" resultid="3687" />
                    <RANKING order="24" place="24" resultid="2314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3929" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2380" />
                    <RANKING order="2" place="2" resultid="2362" />
                    <RANKING order="3" place="3" resultid="3289" />
                    <RANKING order="4" place="4" resultid="2400" />
                    <RANKING order="5" place="5" resultid="2373" />
                    <RANKING order="6" place="6" resultid="3282" />
                    <RANKING order="7" place="7" resultid="3396" />
                    <RANKING order="8" place="8" resultid="2619" />
                    <RANKING order="9" place="9" resultid="3857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3930" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2325" />
                    <RANKING order="2" place="2" resultid="3414" />
                    <RANKING order="3" place="3" resultid="3580" />
                    <RANKING order="4" place="4" resultid="3196" />
                    <RANKING order="5" place="5" resultid="3546" />
                    <RANKING order="6" place="6" resultid="2634" />
                    <RANKING order="7" place="7" resultid="2027" />
                    <RANKING order="8" place="8" resultid="2407" />
                    <RANKING order="9" place="9" resultid="3303" />
                    <RANKING order="10" place="10" resultid="2320" />
                    <RANKING order="11" place="11" resultid="2711" />
                    <RANKING order="12" place="-1" resultid="3091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3931" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2007" />
                    <RANKING order="2" place="2" resultid="2014" />
                    <RANKING order="3" place="-1" resultid="2778" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4089" daytime="16:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4090" daytime="16:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4091" daytime="16:31" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4092" daytime="16:33" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4093" daytime="16:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4094" daytime="16:35" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1419" daytime="16:37" gender="F" number="17" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3932" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="3933" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3165" />
                    <RANKING order="2" place="2" resultid="3173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3934" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3107" />
                    <RANKING order="2" place="2" resultid="3593" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4095" daytime="16:37" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1446" daytime="16:57" gender="M" number="18" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3935" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3147" />
                    <RANKING order="2" place="2" resultid="2629" />
                    <RANKING order="3" place="3" resultid="3598" />
                    <RANKING order="4" place="-1" resultid="2963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3936" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2381" />
                    <RANKING order="2" place="2" resultid="2401" />
                    <RANKING order="3" place="3" resultid="2279" />
                    <RANKING order="4" place="4" resultid="3128" />
                    <RANKING order="5" place="5" resultid="3330" />
                    <RANKING order="6" place="6" resultid="3402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3937" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3134" />
                    <RANKING order="2" place="2" resultid="3203" />
                    <RANKING order="3" place="3" resultid="3209" />
                    <RANKING order="4" place="4" resultid="2411" />
                    <RANKING order="5" place="5" resultid="2596" />
                    <RANKING order="6" place="-1" resultid="3197" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4096" daytime="16:57" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4097" daytime="17:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-05-30" daytime="08:45" endtime="13:18" name="II Blok" number="2" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1451" daytime="08:45" gender="F" number="19" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3938" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3611" />
                    <RANKING order="2" place="2" resultid="2587" />
                    <RANKING order="3" place="3" resultid="2131" />
                    <RANKING order="4" place="4" resultid="2226" />
                    <RANKING order="5" place="5" resultid="3617" />
                    <RANKING order="6" place="6" resultid="3500" />
                    <RANKING order="7" place="7" resultid="3495" />
                    <RANKING order="8" place="8" resultid="2442" />
                    <RANKING order="9" place="9" resultid="2902" />
                    <RANKING order="10" place="10" resultid="3160" />
                    <RANKING order="11" place="11" resultid="2752" />
                    <RANKING order="12" place="12" resultid="3682" />
                    <RANKING order="13" place="13" resultid="3629" />
                    <RANKING order="14" place="14" resultid="2638" />
                    <RANKING order="15" place="15" resultid="2231" />
                    <RANKING order="16" place="16" resultid="3505" />
                    <RANKING order="17" place="17" resultid="2678" />
                    <RANKING order="18" place="-1" resultid="2447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3939" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3604" />
                    <RANKING order="2" place="2" resultid="2832" />
                    <RANKING order="3" place="3" resultid="2119" />
                    <RANKING order="4" place="4" resultid="3352" />
                    <RANKING order="5" place="5" resultid="3511" />
                    <RANKING order="6" place="6" resultid="3087" />
                    <RANKING order="7" place="7" resultid="2054" />
                    <RANKING order="8" place="8" resultid="2124" />
                    <RANKING order="9" place="9" resultid="2220" />
                    <RANKING order="10" place="10" resultid="2060" />
                    <RANKING order="11" place="11" resultid="2530" />
                    <RANKING order="12" place="12" resultid="2136" />
                    <RANKING order="13" place="13" resultid="2648" />
                    <RANKING order="14" place="14" resultid="2851" />
                    <RANKING order="15" place="15" resultid="2667" />
                    <RANKING order="16" place="16" resultid="2653" />
                    <RANKING order="17" place="17" resultid="3024" />
                    <RANKING order="18" place="18" resultid="2658" />
                    <RANKING order="19" place="-1" resultid="3521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3940" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2838" />
                    <RANKING order="2" place="2" resultid="3516" />
                    <RANKING order="3" place="3" resultid="3340" />
                    <RANKING order="4" place="4" resultid="3166" />
                    <RANKING order="5" place="5" resultid="3488" />
                    <RANKING order="6" place="6" resultid="2300" />
                    <RANKING order="7" place="7" resultid="3059" />
                    <RANKING order="8" place="8" resultid="2881" />
                    <RANKING order="9" place="9" resultid="2609" />
                    <RANKING order="10" place="10" resultid="3348" />
                    <RANKING order="11" place="11" resultid="3526" />
                    <RANKING order="12" place="12" resultid="3174" />
                    <RANKING order="13" place="13" resultid="3531" />
                    <RANKING order="14" place="14" resultid="3065" />
                    <RANKING order="15" place="15" resultid="2521" />
                    <RANKING order="16" place="16" resultid="2582" />
                    <RANKING order="17" place="17" resultid="2305" />
                    <RANKING order="18" place="18" resultid="2885" />
                    <RANKING order="19" place="-1" resultid="3096" />
                    <RANKING order="20" place="-1" resultid="3334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3941" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2428" />
                    <RANKING order="2" place="2" resultid="2022" />
                    <RANKING order="3" place="3" resultid="3293" />
                    <RANKING order="4" place="4" resultid="2576" />
                    <RANKING order="5" place="5" resultid="2035" />
                    <RANKING order="6" place="6" resultid="2625" />
                    <RANKING order="7" place="7" resultid="2672" />
                    <RANKING order="8" place="8" resultid="2415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3942" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2765" />
                    <RANKING order="2" place="2" resultid="2770" />
                    <RANKING order="3" place="3" resultid="2761" />
                    <RANKING order="4" place="-1" resultid="2191" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4098" daytime="08:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4099" daytime="08:47" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4100" daytime="08:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4101" daytime="08:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4102" daytime="08:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4103" daytime="08:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4104" daytime="08:58" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4105" daytime="08:59" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1475" daytime="09:01" gender="M" number="20" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3943" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3216" />
                    <RANKING order="2" place="2" resultid="2475" />
                    <RANKING order="3" place="3" resultid="2870" />
                    <RANKING order="4" place="4" resultid="2149" />
                    <RANKING order="5" place="5" resultid="2934" />
                    <RANKING order="6" place="6" resultid="3192" />
                    <RANKING order="7" place="7" resultid="3555" />
                    <RANKING order="8" place="8" resultid="2356" />
                    <RANKING order="9" place="9" resultid="2333" />
                    <RANKING order="10" place="10" resultid="2857" />
                    <RANKING order="11" place="11" resultid="2688" />
                    <RANKING order="12" place="12" resultid="2570" />
                    <RANKING order="13" place="13" resultid="2562" />
                    <RANKING order="14" place="14" resultid="3180" />
                    <RANKING order="15" place="15" resultid="2480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3944" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2953" />
                    <RANKING order="2" place="2" resultid="2350" />
                    <RANKING order="3" place="3" resultid="3224" />
                    <RANKING order="4" place="4" resultid="2705" />
                    <RANKING order="5" place="5" resultid="2462" />
                    <RANKING order="6" place="6" resultid="2242" />
                    <RANKING order="7" place="7" resultid="3560" />
                    <RANKING order="8" place="8" resultid="2716" />
                    <RANKING order="9" place="9" resultid="2155" />
                    <RANKING order="10" place="10" resultid="2699" />
                    <RANKING order="11" place="11" resultid="2545" />
                    <RANKING order="12" place="12" resultid="3450" />
                    <RANKING order="13" place="13" resultid="2253" />
                    <RANKING order="14" place="14" resultid="3230" />
                    <RANKING order="15" place="15" resultid="2367" />
                    <RANKING order="16" place="16" resultid="2486" />
                    <RANKING order="17" place="17" resultid="2339" />
                    <RANKING order="18" place="18" resultid="2694" />
                    <RANKING order="19" place="19" resultid="2641" />
                    <RANKING order="20" place="20" resultid="2946" />
                    <RANKING order="21" place="21" resultid="2940" />
                    <RANKING order="22" place="22" resultid="2142" />
                    <RANKING order="23" place="23" resultid="2863" />
                    <RANKING order="24" place="24" resultid="2958" />
                    <RANKING order="25" place="25" resultid="2491" />
                    <RANKING order="26" place="26" resultid="2497" />
                    <RANKING order="27" place="27" resultid="2923" />
                    <RANKING order="28" place="28" resultid="3186" />
                    <RANKING order="29" place="29" resultid="2512" />
                    <RANKING order="30" place="30" resultid="2507" />
                    <RANKING order="31" place="31" resultid="2248" />
                    <RANKING order="32" place="32" resultid="2683" />
                    <RANKING order="33" place="33" resultid="2502" />
                    <RANKING order="34" place="34" resultid="2315" />
                    <RANKING order="35" place="-1" resultid="2065" />
                    <RANKING order="36" place="-1" resultid="2914" />
                    <RANKING order="37" place="-1" resultid="2964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3945" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2382" />
                    <RANKING order="2" place="2" resultid="2540" />
                    <RANKING order="3" place="3" resultid="2452" />
                    <RANKING order="4" place="4" resultid="2374" />
                    <RANKING order="5" place="5" resultid="3410" />
                    <RANKING order="6" place="6" resultid="3859" />
                    <RANKING order="7" place="7" resultid="3422" />
                    <RANKING order="8" place="7" resultid="3584" />
                    <RANKING order="9" place="9" resultid="3081" />
                    <RANKING order="10" place="10" resultid="2620" />
                    <RANKING order="11" place="11" resultid="3403" />
                    <RANKING order="12" place="12" resultid="2755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3946" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3547" />
                    <RANKING order="2" place="2" resultid="3198" />
                    <RANKING order="3" place="3" resultid="3204" />
                    <RANKING order="4" place="4" resultid="2326" />
                    <RANKING order="5" place="5" resultid="2457" />
                    <RANKING order="6" place="6" resultid="3210" />
                    <RANKING order="7" place="7" resultid="3099" />
                    <RANKING order="8" place="8" resultid="2028" />
                    <RANKING order="9" place="9" resultid="2740" />
                    <RANKING order="10" place="10" resultid="3094" />
                    <RANKING order="11" place="11" resultid="2321" />
                    <RANKING order="12" place="12" resultid="3542" />
                    <RANKING order="13" place="13" resultid="2597" />
                    <RANKING order="14" place="14" resultid="2412" />
                    <RANKING order="15" place="15" resultid="2635" />
                    <RANKING order="16" place="16" resultid="3322" />
                    <RANKING order="17" place="17" resultid="2535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3947" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2181" />
                    <RANKING order="2" place="2" resultid="2814" />
                    <RANKING order="3" place="3" resultid="2790" />
                    <RANKING order="4" place="4" resultid="2774" />
                    <RANKING order="5" place="5" resultid="2786" />
                    <RANKING order="6" place="6" resultid="3102" />
                    <RANKING order="7" place="7" resultid="4226" />
                    <RANKING order="8" place="8" resultid="2113" />
                    <RANKING order="9" place="-1" resultid="2008" />
                    <RANKING order="10" place="-1" resultid="2015" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4106" daytime="09:01" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4107" daytime="09:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4108" daytime="09:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4109" daytime="09:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4110" daytime="09:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4111" daytime="09:13" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4112" daytime="09:14" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4113" daytime="09:16" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4114" daytime="09:18" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4115" daytime="09:19" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1498" daytime="09:21" gender="F" number="21" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3948" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2991" />
                    <RANKING order="2" place="2" resultid="2986" />
                    <RANKING order="3" place="3" resultid="3630" />
                    <RANKING order="4" place="4" resultid="3027" />
                    <RANKING order="5" place="5" resultid="2443" />
                    <RANKING order="6" place="6" resultid="2903" />
                    <RANKING order="7" place="7" resultid="3161" />
                    <RANKING order="8" place="8" resultid="2639" />
                    <RANKING order="9" place="9" resultid="2735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3949" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3072" />
                    <RANKING order="2" place="2" resultid="3359" />
                    <RANKING order="3" place="3" resultid="3438" />
                    <RANKING order="4" place="4" resultid="2970" />
                    <RANKING order="5" place="5" resultid="2981" />
                    <RANKING order="6" place="6" resultid="2654" />
                    <RANKING order="7" place="7" resultid="2897" />
                    <RANKING order="8" place="8" resultid="2309" />
                    <RANKING order="9" place="-1" resultid="2975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3950" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2264" />
                    <RANKING order="2" place="2" resultid="3122" />
                    <RANKING order="3" place="3" resultid="2731" />
                    <RANKING order="4" place="4" resultid="3574" />
                    <RANKING order="5" place="5" resultid="2517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3951" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2726" />
                    <RANKING order="2" place="2" resultid="3108" />
                    <RANKING order="3" place="3" resultid="3242" />
                    <RANKING order="4" place="4" resultid="3484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3952" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2798" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4116" daytime="09:21" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4117" daytime="09:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4118" daytime="09:31" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1521" daytime="09:35" gender="M" number="22" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3953" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2390" />
                    <RANKING order="2" place="2" resultid="4009" />
                    <RANKING order="3" place="3" resultid="3007" />
                    <RANKING order="4" place="4" resultid="2557" />
                    <RANKING order="5" place="5" resultid="2396" />
                    <RANKING order="6" place="6" resultid="2744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3954" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3141" />
                    <RANKING order="2" place="2" resultid="3444" />
                    <RANKING order="3" place="3" resultid="3268" />
                    <RANKING order="4" place="4" resultid="3599" />
                    <RANKING order="5" place="5" resultid="3247" />
                    <RANKING order="6" place="6" resultid="3451" />
                    <RANKING order="7" place="7" resultid="2463" />
                    <RANKING order="8" place="8" resultid="3648" />
                    <RANKING order="9" place="9" resultid="2700" />
                    <RANKING order="10" place="10" resultid="3273" />
                    <RANKING order="11" place="11" resultid="3001" />
                    <RANKING order="12" place="12" resultid="2924" />
                    <RANKING order="13" place="13" resultid="2344" />
                    <RANKING order="14" place="14" resultid="2143" />
                    <RANKING order="15" place="15" resultid="2919" />
                    <RANKING order="16" place="16" resultid="2996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3955" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3253" />
                    <RANKING order="2" place="2" resultid="2271" />
                    <RANKING order="3" place="3" resultid="3082" />
                    <RANKING order="4" place="4" resultid="2287" />
                    <RANKING order="5" place="5" resultid="3263" />
                    <RANKING order="6" place="6" resultid="2549" />
                    <RANKING order="7" place="7" resultid="2756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3956" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3581" />
                    <RANKING order="2" place="2" resultid="3258" />
                    <RANKING order="3" place="3" resultid="3323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3957" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2071" />
                    <RANKING order="2" place="2" resultid="2821" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4119" daytime="09:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4120" daytime="09:39" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4121" daytime="09:43" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4122" daytime="09:47" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1544" daytime="09:51" gender="F" number="23" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1936" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1937" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3115" />
                    <RANKING order="2" place="2" resultid="3456" />
                    <RANKING order="3" place="3" resultid="3461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1938" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3594" />
                    <RANKING order="2" place="2" resultid="3590" />
                    <RANKING order="3" place="3" resultid="2749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1939" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2805" />
                    <RANKING order="2" place="2" resultid="2809" />
                    <RANKING order="3" place="3" resultid="2186" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4123" daytime="09:51" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1567" daytime="09:55" gender="M" number="24" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3958" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2954" />
                    <RANKING order="2" place="2" resultid="3155" />
                    <RANKING order="3" place="3" resultid="2603" />
                    <RANKING order="4" place="4" resultid="3148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3959" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2383" />
                    <RANKING order="2" place="2" resultid="2402" />
                    <RANKING order="3" place="3" resultid="3129" />
                    <RANKING order="4" place="4" resultid="3283" />
                    <RANKING order="5" place="5" resultid="2288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3960" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3135" />
                    <RANKING order="2" place="2" resultid="2421" />
                    <RANKING order="3" place="3" resultid="3415" />
                    <RANKING order="4" place="4" resultid="2598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3961" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2182" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4124" daytime="09:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4125" daytime="09:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1590" daytime="10:02" gender="F" number="25" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3962" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2614" />
                    <RANKING order="2" place="2" resultid="2891" />
                    <RANKING order="3" place="3" resultid="2227" />
                    <RANKING order="4" place="4" resultid="3642" />
                    <RANKING order="5" place="5" resultid="3016" />
                    <RANKING order="6" place="6" resultid="3618" />
                    <RANKING order="7" place="7" resultid="2908" />
                    <RANKING order="8" place="8" resultid="3501" />
                    <RANKING order="9" place="9" resultid="2753" />
                    <RANKING order="10" place="10" resultid="3028" />
                    <RANKING order="11" place="11" resultid="2448" />
                    <RANKING order="12" place="12" resultid="2232" />
                    <RANKING order="13" place="13" resultid="2679" />
                    <RANKING order="14" place="14" resultid="3506" />
                    <RANKING order="15" place="15" resultid="2736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3963" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3468" />
                    <RANKING order="2" place="2" resultid="3353" />
                    <RANKING order="3" place="3" resultid="2833" />
                    <RANKING order="4" place="4" resultid="3667" />
                    <RANKING order="5" place="5" resultid="3237" />
                    <RANKING order="6" place="6" resultid="2055" />
                    <RANKING order="7" place="7" resultid="2221" />
                    <RANKING order="8" place="8" resultid="2137" />
                    <RANKING order="9" place="9" resultid="3537" />
                    <RANKING order="10" place="10" resultid="2649" />
                    <RANKING order="11" place="11" resultid="2659" />
                    <RANKING order="12" place="-1" resultid="3522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3964" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2265" />
                    <RANKING order="2" place="2" resultid="2301" />
                    <RANKING order="3" place="3" resultid="2839" />
                    <RANKING order="4" place="4" resultid="3476" />
                    <RANKING order="5" place="5" resultid="2845" />
                    <RANKING order="6" place="6" resultid="2610" />
                    <RANKING order="7" place="7" resultid="2583" />
                    <RANKING order="8" place="8" resultid="3532" />
                    <RANKING order="9" place="9" resultid="3527" />
                    <RANKING order="10" place="10" resultid="2886" />
                    <RANKING order="11" place="-1" resultid="3335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3965" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2294" />
                    <RANKING order="2" place="2" resultid="3294" />
                    <RANKING order="3" place="3" resultid="2673" />
                    <RANKING order="4" place="4" resultid="2036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3966" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2766" />
                    <RANKING order="2" place="-1" resultid="2192" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4126" daytime="10:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4127" daytime="10:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4128" daytime="10:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4129" daytime="10:09" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4130" daytime="10:11" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1613" daytime="10:13" gender="M" number="26" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3967" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3217" />
                    <RANKING order="2" place="2" resultid="3193" />
                    <RANKING order="3" place="3" resultid="2935" />
                    <RANKING order="4" place="4" resultid="3021" />
                    <RANKING order="5" place="5" resultid="3662" />
                    <RANKING order="6" place="6" resultid="2357" />
                    <RANKING order="7" place="7" resultid="3556" />
                    <RANKING order="8" place="8" resultid="2858" />
                    <RANKING order="9" place="9" resultid="2689" />
                    <RANKING order="10" place="10" resultid="2571" />
                    <RANKING order="11" place="11" resultid="3181" />
                    <RANKING order="12" place="12" resultid="2745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3968" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2468" />
                    <RANKING order="2" place="2" resultid="2243" />
                    <RANKING order="3" place="3" resultid="2706" />
                    <RANKING order="4" place="4" resultid="2929" />
                    <RANKING order="5" place="5" resultid="2254" />
                    <RANKING order="6" place="6" resultid="2717" />
                    <RANKING order="7" place="7" resultid="3002" />
                    <RANKING order="8" place="8" resultid="2642" />
                    <RANKING order="9" place="9" resultid="3654" />
                    <RANKING order="10" place="10" resultid="3623" />
                    <RANKING order="11" place="11" resultid="3187" />
                    <RANKING order="12" place="12" resultid="2941" />
                    <RANKING order="13" place="13" resultid="2508" />
                    <RANKING order="14" place="14" resultid="2503" />
                    <RANKING order="15" place="15" resultid="2684" />
                    <RANKING order="16" place="16" resultid="2249" />
                    <RANKING order="17" place="-1" resultid="2066" />
                    <RANKING order="18" place="-1" resultid="2915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3969" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2874" />
                    <RANKING order="2" place="2" resultid="3290" />
                    <RANKING order="3" place="3" resultid="2272" />
                    <RANKING order="4" place="4" resultid="3397" />
                    <RANKING order="5" place="5" resultid="2621" />
                    <RANKING order="6" place="6" resultid="3585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3970" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3297" />
                    <RANKING order="2" place="2" resultid="2458" />
                    <RANKING order="3" place="3" resultid="2327" />
                    <RANKING order="4" place="4" resultid="2408" />
                    <RANKING order="5" place="5" resultid="3324" />
                    <RANKING order="6" place="6" resultid="2029" />
                    <RANKING order="7" place="-1" resultid="3543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3971" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2791" />
                    <RANKING order="2" place="2" resultid="2815" />
                    <RANKING order="3" place="3" resultid="2072" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4131" daytime="10:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4132" daytime="10:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4133" daytime="10:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4134" daytime="10:21" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4135" daytime="10:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4136" daytime="10:26" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1636" daytime="10:28" gender="F" number="27" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3972" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3973" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3317" />
                    <RANKING order="2" place="2" resultid="3073" />
                    <RANKING order="3" place="3" resultid="3512" />
                    <RANKING order="4" place="4" resultid="3439" />
                    <RANKING order="5" place="5" resultid="2061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3974" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2266" />
                    <RANKING order="2" place="2" resultid="3116" />
                    <RANKING order="3" place="3" resultid="3123" />
                    <RANKING order="4" place="4" resultid="3489" />
                    <RANKING order="5" place="5" resultid="3167" />
                    <RANKING order="6" place="6" resultid="3060" />
                    <RANKING order="7" place="7" resultid="3457" />
                    <RANKING order="8" place="8" resultid="3677" />
                    <RANKING order="9" place="-1" resultid="3575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3975" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2727" />
                    <RANKING order="2" place="2" resultid="2750" />
                    <RANKING order="3" place="3" resultid="2626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3976" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2810" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4137" daytime="10:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4138" daytime="10:32" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1659" daytime="10:36" gender="M" number="28" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3977" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2391" />
                    <RANKING order="2" place="2" resultid="3008" />
                    <RANKING order="3" place="3" resultid="2871" />
                    <RANKING order="4" place="-1" resultid="2481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3978" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2592" />
                    <RANKING order="2" place="2" resultid="2469" />
                    <RANKING order="3" place="3" resultid="3142" />
                    <RANKING order="4" place="4" resultid="3149" />
                    <RANKING order="5" place="5" resultid="3636" />
                    <RANKING order="6" place="6" resultid="3248" />
                    <RANKING order="7" place="7" resultid="3269" />
                    <RANKING order="8" place="8" resultid="3274" />
                    <RANKING order="9" place="9" resultid="3231" />
                    <RANKING order="10" place="10" resultid="2144" />
                    <RANKING order="11" place="11" resultid="3624" />
                    <RANKING order="12" place="12" resultid="2947" />
                    <RANKING order="13" place="13" resultid="2498" />
                    <RANKING order="14" place="14" resultid="2492" />
                    <RANKING order="15" place="15" resultid="3655" />
                    <RANKING order="16" place="-1" resultid="2513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3979" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2273" />
                    <RANKING order="2" place="2" resultid="2280" />
                    <RANKING order="3" place="3" resultid="3130" />
                    <RANKING order="4" place="4" resultid="2541" />
                    <RANKING order="5" place="5" resultid="2375" />
                    <RANKING order="6" place="6" resultid="3254" />
                    <RANKING order="7" place="7" resultid="3284" />
                    <RANKING order="8" place="8" resultid="3264" />
                    <RANKING order="9" place="9" resultid="2289" />
                    <RANKING order="10" place="10" resultid="3860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3980" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3199" />
                    <RANKING order="2" place="2" resultid="3259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3981" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2822" />
                    <RANKING order="2" place="-1" resultid="2016" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4139" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4140" daytime="10:39" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4141" daytime="10:43" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4142" daytime="10:47" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1682" daytime="10:50" gender="F" number="29" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3982" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3612" />
                    <RANKING order="2" place="2" resultid="2588" />
                    <RANKING order="3" place="3" resultid="2987" />
                    <RANKING order="4" place="4" resultid="2909" />
                    <RANKING order="5" place="5" resultid="3017" />
                    <RANKING order="6" place="6" resultid="3683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3983" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2433" />
                    <RANKING order="2" place="2" resultid="3605" />
                    <RANKING order="3" place="3" resultid="3360" />
                    <RANKING order="4" place="4" resultid="2982" />
                    <RANKING order="5" place="5" resultid="2531" />
                    <RANKING order="6" place="6" resultid="3025" />
                    <RANKING order="7" place="7" resultid="2310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3984" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3168" />
                    <RANKING order="2" place="2" resultid="3117" />
                    <RANKING order="3" place="3" resultid="3517" />
                    <RANKING order="4" place="4" resultid="3341" />
                    <RANKING order="5" place="5" resultid="3175" />
                    <RANKING order="6" place="6" resultid="3462" />
                    <RANKING order="7" place="-1" resultid="3097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3985" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3109" />
                    <RANKING order="2" place="2" resultid="2429" />
                    <RANKING order="3" place="3" resultid="3595" />
                    <RANKING order="4" place="4" resultid="2416" />
                    <RANKING order="5" place="5" resultid="3243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3986" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2187" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4143" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4144" daytime="10:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4145" daytime="11:03" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1705" daytime="11:09" gender="M" number="30" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3987" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3278" />
                    <RANKING order="2" place="2" resultid="2476" />
                    <RANKING order="3" place="3" resultid="2150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3988" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2351" />
                    <RANKING order="2" place="2" resultid="3225" />
                    <RANKING order="3" place="3" resultid="3445" />
                    <RANKING order="4" place="4" resultid="2244" />
                    <RANKING order="5" place="5" resultid="2630" />
                    <RANKING order="6" place="6" resultid="3649" />
                    <RANKING order="7" place="7" resultid="4227" />
                    <RANKING order="8" place="8" resultid="3688" />
                    <RANKING order="9" place="9" resultid="2864" />
                    <RANKING order="10" place="10" resultid="2959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3989" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2384" />
                    <RANKING order="2" place="2" resultid="2403" />
                    <RANKING order="3" place="3" resultid="3131" />
                    <RANKING order="4" place="4" resultid="2281" />
                    <RANKING order="5" place="5" resultid="2453" />
                    <RANKING order="6" place="6" resultid="3285" />
                    <RANKING order="7" place="7" resultid="2550" />
                    <RANKING order="8" place="8" resultid="3404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3990" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3205" />
                    <RANKING order="2" place="2" resultid="2422" />
                    <RANKING order="3" place="3" resultid="3211" />
                    <RANKING order="4" place="4" resultid="2413" />
                    <RANKING order="5" place="5" resultid="3416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3991" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3698" />
                    <RANKING order="2" place="2" resultid="2826" />
                    <RANKING order="3" place="3" resultid="2775" />
                    <RANKING order="4" place="4" resultid="3103" />
                    <RANKING order="5" place="5" resultid="2114" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4146" daytime="11:09" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4147" daytime="11:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4148" daytime="11:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4149" daytime="11:29" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1728" daytime="11:34" gender="F" number="31" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3992" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2615" />
                    <RANKING order="2" place="2" resultid="2892" />
                    <RANKING order="3" place="3" resultid="2992" />
                    <RANKING order="4" place="4" resultid="3643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3993" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3318" />
                    <RANKING order="2" place="2" resultid="3469" />
                    <RANKING order="3" place="3" resultid="3668" />
                    <RANKING order="4" place="4" resultid="3354" />
                    <RANKING order="5" place="5" resultid="2120" />
                    <RANKING order="6" place="6" resultid="3672" />
                    <RANKING order="7" place="7" resultid="3238" />
                    <RANKING order="8" place="8" resultid="3538" />
                    <RANKING order="9" place="9" resultid="2898" />
                    <RANKING order="10" place="-1" resultid="2976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3994" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3124" />
                    <RANKING order="2" place="2" resultid="2302" />
                    <RANKING order="3" place="3" resultid="2840" />
                    <RANKING order="4" place="4" resultid="3477" />
                    <RANKING order="5" place="5" resultid="3576" />
                    <RANKING order="6" place="6" resultid="2846" />
                    <RANKING order="7" place="7" resultid="3678" />
                    <RANKING order="8" place="-1" resultid="3336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3995" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2295" />
                    <RANKING order="2" place="2" resultid="2577" />
                    <RANKING order="3" place="3" resultid="3295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3996" agemax="-1" agemin="25" name="Open Masters" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4150" daytime="11:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4151" daytime="11:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4152" daytime="11:42" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1751" daytime="11:45" gender="M" number="32" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3997" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3218" />
                    <RANKING order="2" place="2" resultid="2392" />
                    <RANKING order="3" place="3" resultid="4010" />
                    <RANKING order="4" place="4" resultid="2936" />
                    <RANKING order="5" place="5" resultid="3279" />
                    <RANKING order="6" place="6" resultid="2558" />
                    <RANKING order="7" place="7" resultid="3022" />
                    <RANKING order="8" place="8" resultid="2358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3998" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2470" />
                    <RANKING order="2" place="2" resultid="2604" />
                    <RANKING order="3" place="3" resultid="2593" />
                    <RANKING order="4" place="4" resultid="2930" />
                    <RANKING order="5" place="5" resultid="3249" />
                    <RANKING order="6" place="6" resultid="3232" />
                    <RANKING order="7" place="7" resultid="2865" />
                    <RANKING order="8" place="8" resultid="3656" />
                    <RANKING order="9" place="9" resultid="2316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3999" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2875" />
                    <RANKING order="2" place="2" resultid="2274" />
                    <RANKING order="3" place="3" resultid="3291" />
                    <RANKING order="4" place="4" resultid="3398" />
                    <RANKING order="5" place="5" resultid="3586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4000" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3298" />
                    <RANKING order="2" place="2" resultid="2636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4001" agemax="-1" agemin="25" name="Open Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2823" />
                    <RANKING order="2" place="-1" resultid="2818" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4153" daytime="11:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4154" daytime="11:49" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4155" daytime="11:53" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1774" daytime="11:57" gender="F" number="33" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4002" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2434" />
                    <RANKING order="2" place="2" resultid="3088" />
                    <RANKING order="3" place="3" resultid="2125" />
                    <RANKING order="4" place="4" resultid="3673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4003" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3169" />
                    <RANKING order="2" place="2" resultid="3490" />
                    <RANKING order="3" place="3" resultid="3066" />
                    <RANKING order="4" place="4" resultid="3342" />
                    <RANKING order="5" place="5" resultid="3176" />
                    <RANKING order="6" place="6" resultid="3463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4004" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3110" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4156" daytime="11:57" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4157" daytime="12:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1797" daytime="12:19" gender="M" number="34" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4005" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3150" />
                    <RANKING order="2" place="2" resultid="3143" />
                    <RANKING order="3" place="3" resultid="3156" />
                    <RANKING order="4" place="4" resultid="3637" />
                    <RANKING order="5" place="5" resultid="2631" />
                    <RANKING order="6" place="6" resultid="3600" />
                    <RANKING order="7" place="7" resultid="3561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4006" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2385" />
                    <RANKING order="2" place="2" resultid="2404" />
                    <RANKING order="3" place="3" resultid="2282" />
                    <RANKING order="4" place="4" resultid="2275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4007" agemax="24" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3136" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4158" daytime="12:19" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4159" daytime="12:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="00905" nation="POL" region="05" clubid="2417" name="MKS Trójka Łódź">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Sekściński" birthdate="2009-10-03" gender="M" nation="POL" license="100905700404" swrid="5260899" athleteid="2471">
              <RESULTS>
                <RESULT eventid="1120" points="350" reactiontime="+64" swimtime="00:00:29.67" resultid="2472" heatid="4029" lane="8" entrytime="00:00:30.72" entrycourse="LCM" />
                <RESULT eventid="1304" points="330" reactiontime="+55" swimtime="00:02:27.52" resultid="2473" heatid="4070" lane="9" entrytime="00:02:26.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                    <SPLIT distance="150" swimtime="00:01:52.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="327" reactiontime="+67" swimtime="00:00:32.30" resultid="2474" heatid="4092" lane="9" entrytime="00:00:33.08" entrycourse="LCM" />
                <RESULT eventid="1475" points="346" reactiontime="+72" swimtime="00:01:06.79" resultid="2475" heatid="4112" lane="0" entrytime="00:01:06.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="314" reactiontime="+54" swimtime="00:05:23.59" resultid="2476" heatid="4147" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:18.97" />
                    <SPLIT distance="150" swimtime="00:02:01.00" />
                    <SPLIT distance="200" swimtime="00:02:42.88" />
                    <SPLIT distance="250" swimtime="00:03:24.86" />
                    <SPLIT distance="300" swimtime="00:04:06.69" />
                    <SPLIT distance="350" swimtime="00:04:47.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Franciszek" lastname="Janiszewski" birthdate="2009-01-14" gender="M" nation="POL" license="100905700413" swrid="5260890" athleteid="2563">
              <RESULTS>
                <RESULT eventid="1166" status="DNS" swimtime="00:00:00.00" resultid="2564" heatid="4039" lane="3" entrytime="00:00:49.30" entrycourse="LCM" />
                <RESULT eventid="1258" status="DNS" swimtime="00:00:00.00" resultid="2565" heatid="4057" lane="4" entrytime="00:00:43.08" entrycourse="LCM" />
                <RESULT eventid="1350" status="DNS" swimtime="00:00:00.00" resultid="2566" heatid="4078" lane="3" entrytime="00:01:43.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Dziśnieńska" birthdate="2007-03-27" gender="F" nation="POL" license="100905600346" swrid="5225034" athleteid="2522">
              <RESULTS>
                <RESULT eventid="1143" points="257" reactiontime="+93" swimtime="00:00:46.23" resultid="2523" heatid="4035" lane="0" entrytime="00:00:45.82" entrycourse="LCM" />
                <RESULT eventid="1235" points="168" reactiontime="+86" swimtime="00:00:48.83" resultid="2524" heatid="4051" lane="2" />
                <RESULT eventid="1327" points="213" swimtime="00:01:47.25" resultid="2525" heatid="4074" lane="8" entrytime="00:01:38.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Feliks" lastname="Rubin" birthdate="2008-01-31" gender="M" nation="POL" license="100905700428" swrid="5197994" athleteid="2459">
              <RESULTS>
                <RESULT eventid="1120" points="416" reactiontime="+84" swimtime="00:00:27.99" resultid="2460" heatid="4030" lane="1" entrytime="00:00:28.38" entrycourse="LCM" />
                <RESULT eventid="1304" points="449" reactiontime="+77" swimtime="00:02:13.14" resultid="2461" heatid="4071" lane="9" entrytime="00:02:13.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:05.12" />
                    <SPLIT distance="150" swimtime="00:01:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="462" reactiontime="+79" swimtime="00:01:00.65" resultid="2462" heatid="4113" lane="0" entrytime="00:01:01.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="342" reactiontime="+66" swimtime="00:03:00.33" resultid="2463" heatid="4120" lane="5" entrytime="00:03:12.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:26.96" />
                    <SPLIT distance="150" swimtime="00:02:13.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymoteusz" lastname="Kaczmarek" birthdate="2008-01-22" gender="M" nation="POL" license="100905700387" swrid="5093347" athleteid="2551">
              <RESULTS>
                <RESULT eventid="1166" points="269" reactiontime="+58" swimtime="00:00:40.16" resultid="2552" heatid="4040" lane="2" entrytime="00:00:43.66" entrycourse="LCM" />
                <RESULT eventid="1350" points="249" swimtime="00:01:30.38" resultid="2553" heatid="4079" lane="0" entrytime="00:01:34.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Dziśnieński" birthdate="2009-08-17" gender="M" nation="POL" license="100905700419" swrid="5331235" athleteid="2559">
              <RESULTS>
                <RESULT eventid="1166" points="166" reactiontime="+56" swimtime="00:00:47.18" resultid="2560" heatid="4040" lane="9" entrytime="00:00:47.41" entrycourse="LCM" />
                <RESULT eventid="1350" points="136" reactiontime="+70" swimtime="00:01:50.35" resultid="2561" heatid="4078" lane="7" entrytime="00:01:46.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="120" reactiontime="+72" swimtime="00:01:34.97" resultid="2562" heatid="4109" lane="6" entrytime="00:01:32.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Jędrzejak" birthdate="2009-08-26" gender="F" nation="POL" license="100905600423" swrid="4977215" athleteid="2439">
              <RESULTS>
                <RESULT eventid="1070" points="268" reactiontime="+89" swimtime="00:00:36.67" resultid="2440" heatid="4017" lane="2" entrytime="00:00:35.72" entrycourse="LCM" />
                <RESULT eventid="1143" points="244" reactiontime="+82" swimtime="00:00:47.03" resultid="2441" heatid="4034" lane="4" entrytime="00:00:46.63" entrycourse="LCM" />
                <RESULT eventid="1451" points="272" reactiontime="+78" swimtime="00:01:19.74" resultid="2442" heatid="4101" lane="8" entrytime="00:01:19.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="264" reactiontime="+96" swimtime="00:03:36.82" resultid="2443" heatid="4117" lane="0" entrytime="00:03:30.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.13" />
                    <SPLIT distance="100" swimtime="00:01:44.87" />
                    <SPLIT distance="150" swimtime="00:02:40.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Milczarczyk" birthdate="2008-12-08" gender="M" nation="POL" license="100905700390" swrid="5094215" athleteid="2504">
              <RESULTS>
                <RESULT eventid="1120" points="220" reactiontime="+71" swimtime="00:00:34.63" resultid="2505" heatid="4027" lane="0" entrytime="00:00:35.51" entrycourse="LCM" />
                <RESULT eventid="1166" points="197" swimtime="00:00:44.58" resultid="2506" heatid="4040" lane="0" entrytime="00:00:47.19" entrycourse="LCM" />
                <RESULT eventid="1475" points="217" reactiontime="+75" swimtime="00:01:18.04" resultid="2507" heatid="4108" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="177" reactiontime="+74" swimtime="00:01:32.19" resultid="2508" heatid="4134" lane="1" entrytime="00:01:35.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kazimierz" lastname="Janeczek" birthdate="2008-07-16" gender="M" nation="POL" license="100905700389" swrid="5096066" athleteid="2493">
              <RESULTS>
                <RESULT eventid="1120" points="230" reactiontime="+85" swimtime="00:00:34.12" resultid="2494" heatid="4024" lane="5" />
                <RESULT eventid="1304" points="223" reactiontime="+92" swimtime="00:02:47.96" resultid="2495" heatid="4069" lane="0" entrytime="00:02:46.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:22.15" />
                    <SPLIT distance="150" swimtime="00:02:06.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="202" reactiontime="+90" swimtime="00:00:37.95" resultid="2496" heatid="4091" lane="1" entrytime="00:00:37.77" entrycourse="LCM" />
                <RESULT eventid="1475" points="247" reactiontime="+87" swimtime="00:01:14.71" resultid="2497" heatid="4110" lane="8" entrytime="00:01:16.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="236" reactiontime="+69" swimtime="00:03:04.22" resultid="2498" heatid="4141" lane="9" entrytime="00:03:02.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:28.84" />
                    <SPLIT distance="150" swimtime="00:02:25.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystian" lastname="Selder" birthdate="2007-06-18" gender="M" nation="POL" license="100905700353" swrid="5197962" athleteid="2627">
              <RESULTS>
                <RESULT eventid="1304" points="329" reactiontime="+81" swimtime="00:02:27.69" resultid="2628" heatid="4070" lane="5" entrytime="00:02:14.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:10.30" />
                    <SPLIT distance="150" swimtime="00:01:49.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="492" reactiontime="+76" swimtime="00:09:32.47" resultid="2629" heatid="4097" lane="8" entrytime="00:09:43.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="150" swimtime="00:01:44.80" />
                    <SPLIT distance="200" swimtime="00:02:20.35" />
                    <SPLIT distance="250" swimtime="00:02:56.03" />
                    <SPLIT distance="300" swimtime="00:03:31.96" />
                    <SPLIT distance="350" swimtime="00:04:08.33" />
                    <SPLIT distance="400" swimtime="00:04:44.75" />
                    <SPLIT distance="450" swimtime="00:05:21.09" />
                    <SPLIT distance="500" swimtime="00:05:57.26" />
                    <SPLIT distance="550" swimtime="00:06:33.48" />
                    <SPLIT distance="600" swimtime="00:07:09.98" />
                    <SPLIT distance="650" swimtime="00:07:46.36" />
                    <SPLIT distance="700" swimtime="00:08:22.31" />
                    <SPLIT distance="750" swimtime="00:08:57.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="370" reactiontime="+73" swimtime="00:05:06.49" resultid="2630" heatid="4149" lane="9" entrytime="00:04:34.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:51.18" />
                    <SPLIT distance="200" swimtime="00:02:30.52" />
                    <SPLIT distance="250" swimtime="00:03:09.64" />
                    <SPLIT distance="300" swimtime="00:03:49.41" />
                    <SPLIT distance="350" swimtime="00:04:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="504" reactiontime="+80" swimtime="00:18:14.16" resultid="2631" heatid="4159" lane="7" entrytime="00:18:24.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:45.08" />
                    <SPLIT distance="200" swimtime="00:02:20.90" />
                    <SPLIT distance="250" swimtime="00:02:56.66" />
                    <SPLIT distance="300" swimtime="00:03:32.83" />
                    <SPLIT distance="350" swimtime="00:04:08.52" />
                    <SPLIT distance="400" swimtime="00:04:44.29" />
                    <SPLIT distance="450" swimtime="00:05:19.95" />
                    <SPLIT distance="500" swimtime="00:05:56.04" />
                    <SPLIT distance="550" swimtime="00:06:32.73" />
                    <SPLIT distance="600" swimtime="00:07:09.20" />
                    <SPLIT distance="650" swimtime="00:07:45.67" />
                    <SPLIT distance="700" swimtime="00:08:22.07" />
                    <SPLIT distance="750" swimtime="00:08:58.62" />
                    <SPLIT distance="800" swimtime="00:09:35.07" />
                    <SPLIT distance="850" swimtime="00:10:12.08" />
                    <SPLIT distance="900" swimtime="00:10:49.07" />
                    <SPLIT distance="950" swimtime="00:11:25.56" />
                    <SPLIT distance="1000" swimtime="00:12:02.96" />
                    <SPLIT distance="1050" swimtime="00:12:40.12" />
                    <SPLIT distance="1100" swimtime="00:13:17.62" />
                    <SPLIT distance="1150" swimtime="00:13:55.05" />
                    <SPLIT distance="1200" swimtime="00:14:32.49" />
                    <SPLIT distance="1250" swimtime="00:15:09.95" />
                    <SPLIT distance="1300" swimtime="00:15:47.49" />
                    <SPLIT distance="1350" swimtime="00:16:25.02" />
                    <SPLIT distance="1400" swimtime="00:17:02.30" />
                    <SPLIT distance="1450" swimtime="00:17:39.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julian" lastname="Świderski" birthdate="2006-02-19" gender="M" nation="POL" license="100905700340" swrid="5170220" athleteid="2449">
              <RESULTS>
                <RESULT eventid="1120" points="519" reactiontime="+65" swimtime="00:00:26.01" resultid="2450" heatid="4031" lane="4" entrytime="00:00:25.72" entrycourse="LCM" />
                <RESULT eventid="1304" points="508" reactiontime="+68" swimtime="00:02:07.83" resultid="2451" heatid="4072" lane="1" entrytime="00:02:04.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                    <SPLIT distance="100" swimtime="00:01:00.54" />
                    <SPLIT distance="150" swimtime="00:01:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="573" reactiontime="+66" swimtime="00:00:56.45" resultid="2452" heatid="4114" lane="4" entrytime="00:00:56.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="512" reactiontime="+66" swimtime="00:04:35.02" resultid="2453" heatid="4148" lane="4" entrytime="00:04:35.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.82" />
                    <SPLIT distance="150" swimtime="00:01:44.43" />
                    <SPLIT distance="200" swimtime="00:02:20.59" />
                    <SPLIT distance="250" swimtime="00:02:56.20" />
                    <SPLIT distance="300" swimtime="00:03:31.19" />
                    <SPLIT distance="350" swimtime="00:04:05.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Ledzion" birthdate="2006-10-31" gender="M" nation="POL" license="100905700599" swrid="5025339" athleteid="2546">
              <RESULTS>
                <RESULT eventid="1166" points="420" reactiontime="+78" swimtime="00:00:34.64" resultid="2547" heatid="4042" lane="1" entrytime="00:00:35.84" entrycourse="LCM" />
                <RESULT eventid="1304" points="436" reactiontime="+77" swimtime="00:02:14.46" resultid="2548" heatid="4068" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                    <SPLIT distance="100" swimtime="00:01:05.12" />
                    <SPLIT distance="150" swimtime="00:01:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="416" reactiontime="+75" swimtime="00:02:48.93" resultid="2549" heatid="4122" lane="8" entrytime="00:02:44.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:20.01" />
                    <SPLIT distance="150" swimtime="00:02:04.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="475" reactiontime="+79" swimtime="00:04:41.97" resultid="2550" heatid="4147" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="100" swimtime="00:01:07.12" />
                    <SPLIT distance="150" swimtime="00:01:43.46" />
                    <SPLIT distance="200" swimtime="00:02:19.41" />
                    <SPLIT distance="250" swimtime="00:02:55.98" />
                    <SPLIT distance="300" swimtime="00:03:32.37" />
                    <SPLIT distance="350" swimtime="00:04:08.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nikodem" lastname="Jędryka" birthdate="2004-09-14" gender="M" nation="POL" license="100905700429" swrid="5034796" athleteid="2418">
              <RESULTS>
                <RESULT eventid="1065" points="534" reactiontime="+69" swimtime="00:05:00.44" resultid="2419" heatid="4013" lane="6" entrytime="00:04:58.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:01:05.29" />
                    <SPLIT distance="150" swimtime="00:01:43.84" />
                    <SPLIT distance="200" swimtime="00:02:23.47" />
                    <SPLIT distance="250" swimtime="00:03:08.68" />
                    <SPLIT distance="300" swimtime="00:03:52.45" />
                    <SPLIT distance="350" swimtime="00:04:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="602" reactiontime="+69" swimtime="00:02:00.76" resultid="2420" heatid="4072" lane="6" entrytime="00:02:00.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                    <SPLIT distance="100" swimtime="00:00:58.47" />
                    <SPLIT distance="150" swimtime="00:01:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="570" reactiontime="+69" swimtime="00:02:13.54" resultid="2421" heatid="4125" lane="2" entrytime="00:02:12.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="100" swimtime="00:01:02.85" />
                    <SPLIT distance="150" swimtime="00:01:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="640" reactiontime="+67" swimtime="00:04:15.34" resultid="2422" heatid="4149" lane="2" entrytime="00:04:18.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:01:00.71" />
                    <SPLIT distance="150" swimtime="00:01:33.07" />
                    <SPLIT distance="200" swimtime="00:02:06.19" />
                    <SPLIT distance="250" swimtime="00:02:38.95" />
                    <SPLIT distance="300" swimtime="00:03:12.11" />
                    <SPLIT distance="350" swimtime="00:03:45.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Węgrzycka" birthdate="2007-01-04" gender="F" nation="POL" license="100905600363" swrid="5197964" athleteid="2430">
              <RESULTS>
                <RESULT eventid="1070" points="497" reactiontime="+77" swimtime="00:00:29.88" resultid="2431" heatid="4020" lane="5" entrytime="00:00:29.90" entrycourse="LCM" />
                <RESULT eventid="1281" points="536" reactiontime="+74" swimtime="00:02:19.07" resultid="2432" heatid="4064" lane="7" entrytime="00:02:21.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:07.05" />
                    <SPLIT distance="150" swimtime="00:01:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="461" reactiontime="+74" swimtime="00:05:05.92" resultid="2433" heatid="4145" lane="9" entrytime="00:04:58.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:51.01" />
                    <SPLIT distance="200" swimtime="00:02:29.40" />
                    <SPLIT distance="250" swimtime="00:03:08.79" />
                    <SPLIT distance="300" swimtime="00:03:49.02" />
                    <SPLIT distance="350" swimtime="00:04:28.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="510" reactiontime="+74" swimtime="00:10:06.53" resultid="2434" heatid="4156" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:10.02" />
                    <SPLIT distance="150" swimtime="00:01:47.97" />
                    <SPLIT distance="200" swimtime="00:02:25.98" />
                    <SPLIT distance="250" swimtime="00:03:03.91" />
                    <SPLIT distance="300" swimtime="00:03:42.63" />
                    <SPLIT distance="350" swimtime="00:04:20.65" />
                    <SPLIT distance="400" swimtime="00:04:58.93" />
                    <SPLIT distance="450" swimtime="00:05:37.93" />
                    <SPLIT distance="500" swimtime="00:06:16.68" />
                    <SPLIT distance="550" swimtime="00:06:55.27" />
                    <SPLIT distance="600" swimtime="00:07:33.92" />
                    <SPLIT distance="650" swimtime="00:08:12.97" />
                    <SPLIT distance="700" swimtime="00:08:51.43" />
                    <SPLIT distance="750" swimtime="00:09:29.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Jakubowski" birthdate="2008-06-17" gender="M" nation="POL" license="100905700385" swrid="5096063" athleteid="2487">
              <RESULTS>
                <RESULT eventid="1120" points="255" reactiontime="+82" swimtime="00:00:32.96" resultid="2488" heatid="4026" lane="5" entrytime="00:00:36.65" entrycourse="LCM" />
                <RESULT eventid="1258" points="227" reactiontime="+91" swimtime="00:00:39.29" resultid="2489" heatid="4058" lane="0" entrytime="00:00:42.87" entrycourse="LCM" />
                <RESULT eventid="1396" points="160" reactiontime="+77" swimtime="00:00:40.97" resultid="2490" heatid="4089" lane="4" />
                <RESULT eventid="1475" points="255" reactiontime="+92" swimtime="00:01:13.91" resultid="2491" heatid="4108" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="215" reactiontime="+85" swimtime="00:03:10.08" resultid="2492" heatid="4140" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:32.98" />
                    <SPLIT distance="150" swimtime="00:02:30.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Piątkiewicz" birthdate="2007-04-11" gender="M" nation="POL" license="100905700351" swrid="5197967" athleteid="2599">
              <RESULTS>
                <RESULT eventid="1212" points="426" reactiontime="+64" swimtime="00:01:05.74" resultid="2600" heatid="4049" lane="0" entrytime="00:01:07.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="430" reactiontime="+66" swimtime="00:02:15.11" resultid="2601" heatid="4067" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:06.50" />
                    <SPLIT distance="150" swimtime="00:01:41.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="449" reactiontime="+66" swimtime="00:00:29.08" resultid="2602" heatid="4092" lane="4" entrytime="00:00:29.27" entrycourse="LCM" />
                <RESULT eventid="1567" points="448" reactiontime="+69" swimtime="00:02:24.66" resultid="2603" heatid="4125" lane="0" entrytime="00:02:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:07.79" />
                    <SPLIT distance="150" swimtime="00:01:46.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="448" reactiontime="+69" swimtime="00:02:26.21" resultid="2604" heatid="4155" lane="9" entrytime="00:02:26.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="150" swimtime="00:01:50.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Walas" birthdate="2004-01-17" gender="M" nation="POL" license="100905700437" swrid="5034877" athleteid="2532">
              <RESULTS>
                <RESULT eventid="1166" points="412" reactiontime="+71" swimtime="00:00:34.85" resultid="2533" heatid="4042" lane="3" entrytime="00:00:34.37" entrycourse="LCM" />
                <RESULT eventid="1350" points="397" reactiontime="+72" swimtime="00:01:17.36" resultid="2534" heatid="4080" lane="5" entrytime="00:01:16.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="435" reactiontime="+73" swimtime="00:01:01.87" resultid="2535" heatid="4113" lane="9" entrytime="00:01:01.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Świderski" birthdate="2008-03-04" gender="M" nation="POL" license="100905700384" swrid="5170219" athleteid="2589">
              <RESULTS>
                <RESULT eventid="1212" points="415" reactiontime="+80" swimtime="00:01:06.33" resultid="2590" heatid="4049" lane="1" entrytime="00:01:06.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="404" reactiontime="+80" swimtime="00:00:32.45" resultid="2591" heatid="4059" lane="0" entrytime="00:00:35.83" entrycourse="LCM" />
                <RESULT eventid="1659" points="482" reactiontime="+76" swimtime="00:02:25.30" resultid="2592" heatid="4142" lane="9" entrytime="00:02:29.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:52.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="422" reactiontime="+84" swimtime="00:02:29.12" resultid="2593" heatid="4154" lane="4" entrytime="00:02:28.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="100" swimtime="00:01:11.79" />
                    <SPLIT distance="150" swimtime="00:01:51.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Padyk" birthdate="2008-03-17" gender="M" nation="POL" license="100905700391" swrid="4976662" athleteid="2509">
              <RESULTS>
                <RESULT eventid="1120" points="229" reactiontime="+83" swimtime="00:00:34.17" resultid="2510" heatid="4027" lane="7" entrytime="00:00:33.99" entrycourse="LCM" />
                <RESULT eventid="1396" points="178" reactiontime="+87" swimtime="00:00:39.53" resultid="2511" heatid="4091" lane="0" entrytime="00:00:39.58" entrycourse="LCM" />
                <RESULT eventid="1475" points="228" reactiontime="+94" swimtime="00:01:16.72" resultid="2512" heatid="4110" lane="0" entrytime="00:01:19.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu." eventid="1659" reactiontime="+88" status="DSQ" swimtime="00:03:23.11" resultid="2513" heatid="4139" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="100" swimtime="00:01:34.35" />
                    <SPLIT distance="150" swimtime="00:02:38.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Lewenhaupt" birthdate="2006-01-09" gender="M" nation="POL" license="100905700338" swrid="4686775" athleteid="2536">
              <RESULTS>
                <RESULT eventid="1166" points="561" reactiontime="+76" swimtime="00:00:31.45" resultid="2537" heatid="4043" lane="6" entrytime="00:00:31.77" entrycourse="LCM" />
                <RESULT eventid="1212" points="515" reactiontime="+82" swimtime="00:01:01.72" resultid="2538" heatid="4050" lane="0" entrytime="00:01:01.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="498" reactiontime="+75" swimtime="00:01:11.74" resultid="2539" heatid="4081" lane="3" entrytime="00:01:08.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="595" reactiontime="+73" swimtime="00:00:55.75" resultid="2540" heatid="4114" lane="6" entrytime="00:00:56.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="524" reactiontime="+76" swimtime="00:02:21.37" resultid="2541" heatid="4142" lane="3" entrytime="00:02:18.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                    <SPLIT distance="100" swimtime="00:01:07.28" />
                    <SPLIT distance="150" swimtime="00:01:48.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Pawłowska" birthdate="2006-06-10" gender="F" nation="POL" license="100905600598" swrid="5170217" athleteid="2578">
              <RESULTS>
                <RESULT eventid="1189" points="357" reactiontime="+77" swimtime="00:01:18.15" resultid="2579" heatid="4044" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="370" reactiontime="+77" swimtime="00:02:37.25" resultid="2580" heatid="4061" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:01:56.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="334" reactiontime="+76" swimtime="00:00:35.20" resultid="2581" heatid="4086" lane="6" entrytime="00:00:35.24" entrycourse="LCM" />
                <RESULT eventid="1451" points="361" reactiontime="+82" swimtime="00:01:12.61" resultid="2582" heatid="4099" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="387" reactiontime="+64" swimtime="00:01:18.95" resultid="2583" heatid="4129" lane="7" entrytime="00:01:18.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Kowalczyk" birthdate="2004-12-01" gender="F" nation="POL" license="100905600241" swrid="4941665" athleteid="2423">
              <RESULTS>
                <RESULT eventid="1070" points="544" reactiontime="+69" swimtime="00:00:28.98" resultid="2424" heatid="4020" lane="4" entrytime="00:00:29.86" entrycourse="LCM" />
                <RESULT eventid="1143" points="606" reactiontime="+67" swimtime="00:00:34.73" resultid="2425" heatid="4037" lane="6" entrytime="00:00:35.04" entrycourse="LCM" />
                <RESULT eventid="1189" points="532" reactiontime="+65" swimtime="00:01:08.44" resultid="2426" heatid="4046" lane="9" entrytime="00:01:09.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="599" reactiontime="+67" swimtime="00:02:13.97" resultid="2427" heatid="4065" lane="7" entrytime="00:02:17.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:05.57" />
                    <SPLIT distance="150" swimtime="00:01:40.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="573" reactiontime="+69" swimtime="00:01:02.24" resultid="2428" heatid="4104" lane="4" entrytime="00:01:03.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="586" reactiontime="+67" swimtime="00:04:42.41" resultid="2429" heatid="4143" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:07.43" />
                    <SPLIT distance="150" swimtime="00:01:43.56" />
                    <SPLIT distance="200" swimtime="00:02:19.44" />
                    <SPLIT distance="250" swimtime="00:02:55.16" />
                    <SPLIT distance="300" swimtime="00:03:31.32" />
                    <SPLIT distance="350" swimtime="00:04:07.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Koch" birthdate="2006-07-07" gender="M" nation="POL" license="100905700329" swrid="5195505" athleteid="2616">
              <RESULTS>
                <RESULT eventid="1258" points="500" reactiontime="+62" swimtime="00:00:30.23" resultid="2617" heatid="4059" lane="4" entrytime="00:00:30.26" entrycourse="LCM" />
                <RESULT eventid="1304" points="405" reactiontime="+75" swimtime="00:02:17.75" resultid="2618" heatid="4070" lane="4" entrytime="00:02:14.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="450" reactiontime="+82" swimtime="00:00:29.04" resultid="2619" heatid="4093" lane="0" entrytime="00:00:28.39" entrycourse="LCM" />
                <RESULT eventid="1475" points="436" reactiontime="+79" swimtime="00:01:01.84" resultid="2620" heatid="4114" lane="1" entrytime="00:00:57.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="448" reactiontime="+73" swimtime="00:01:07.76" resultid="2621" heatid="4136" lane="0" entrytime="00:01:04.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Piątkiewicz" birthdate="2009-01-09" gender="F" nation="POL" license="100905600403" swrid="5260908" athleteid="2611">
              <RESULTS>
                <RESULT eventid="1235" points="421" reactiontime="+69" swimtime="00:00:35.99" resultid="2612" heatid="4051" lane="3" />
                <RESULT eventid="1373" points="288" reactiontime="+76" swimtime="00:00:36.98" resultid="2613" heatid="4083" lane="9" />
                <RESULT eventid="1590" points="381" reactiontime="+69" swimtime="00:01:19.40" resultid="2614" heatid="4126" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="382" reactiontime="+71" swimtime="00:02:49.98" resultid="2615" heatid="4150" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                    <SPLIT distance="100" swimtime="00:01:25.75" />
                    <SPLIT distance="150" swimtime="00:02:10.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonina" lastname="Zys" birthdate="2007-06-18" gender="F" nation="POL" license="100905600359" swrid="5093449" athleteid="2435">
              <RESULTS>
                <RESULT eventid="1070" status="DNS" swimtime="00:00:00.00" resultid="2436" heatid="4015" lane="4" />
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="2437" heatid="4033" lane="4" />
                <RESULT eventid="1327" status="DNS" swimtime="00:00:00.00" resultid="2438" heatid="4073" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Żelaskowska" birthdate="2009-01-27" gender="F" nation="POL" license="100905600439" swrid="5254125" athleteid="2584">
              <RESULTS>
                <RESULT eventid="1189" points="283" reactiontime="+73" swimtime="00:01:24.45" resultid="2585" heatid="4044" lane="4" entrytime="00:01:26.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="418" reactiontime="+72" swimtime="00:02:31.08" resultid="2586" heatid="4063" lane="1" entrytime="00:02:33.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:54.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="427" reactiontime="+83" swimtime="00:01:08.63" resultid="2587" heatid="4102" lane="6" entrytime="00:01:08.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="436" reactiontime="+56" swimtime="00:05:11.67" resultid="2588" heatid="4144" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:52.27" />
                    <SPLIT distance="200" swimtime="00:02:32.44" />
                    <SPLIT distance="250" swimtime="00:03:13.90" />
                    <SPLIT distance="300" swimtime="00:03:54.04" />
                    <SPLIT distance="350" swimtime="00:04:34.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Olczak" birthdate="2004-09-15" gender="M" nation="POL" license="100905700250" swrid="4971376" athleteid="2454">
              <RESULTS>
                <RESULT eventid="1120" points="574" reactiontime="+69" swimtime="00:00:25.15" resultid="2455" heatid="4032" lane="0" entrytime="00:00:25.39" entrycourse="LCM" />
                <RESULT eventid="1212" points="539" reactiontime="+69" swimtime="00:01:00.79" resultid="2456" heatid="4050" lane="1" entrytime="00:01:00.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="666" reactiontime="+64" swimtime="00:00:53.71" resultid="2457" heatid="4115" lane="7" entrytime="00:00:53.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="601" reactiontime="+88" swimtime="00:01:01.43" resultid="2458" heatid="4136" lane="1" entrytime="00:01:03.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Sieroń" birthdate="2007-07-14" gender="M" nation="POL" license="100905700354" swrid="5225027" athleteid="2482">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1120" status="DSQ" swimtime="00:00:30.95" resultid="2483" heatid="4028" lane="7" entrytime="00:00:31.64" entrycourse="LCM" />
                <RESULT eventid="1166" points="245" reactiontime="+71" swimtime="00:00:41.45" resultid="2484" heatid="4041" lane="8" entrytime="00:00:40.89" entrycourse="LCM" />
                <RESULT eventid="1350" points="243" reactiontime="+76" swimtime="00:01:31.03" resultid="2485" heatid="4078" lane="2" entrytime="00:01:44.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="306" reactiontime="+75" swimtime="00:01:09.57" resultid="2486" heatid="4111" lane="1" entrytime="00:01:09.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ziemowit" lastname="Walasiak" birthdate="2007-01-26" gender="M" nation="POL" license="100905700399" swrid="5225098" athleteid="2640">
              <RESULTS>
                <RESULT eventid="1475" points="295" reactiontime="+85" swimtime="00:01:10.43" resultid="2641" heatid="4111" lane="8" entrytime="00:01:09.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="237" reactiontime="+89" swimtime="00:01:23.74" resultid="2642" heatid="4135" lane="9" entrytime="00:01:21.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roksana" lastname="Kałczak" birthdate="2009-04-04" gender="F" nation="POL" license="100905600414" swrid="4976976" athleteid="2637">
              <RESULTS>
                <RESULT eventid="1451" points="213" swimtime="00:01:26.54" resultid="2638" heatid="4100" lane="7" entrytime="00:01:26.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="187" reactiontime="+93" swimtime="00:04:03.02" resultid="2639" heatid="4116" lane="4" entrytime="00:04:05.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.63" />
                    <SPLIT distance="100" swimtime="00:01:58.48" />
                    <SPLIT distance="150" swimtime="00:03:00.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Krysiak" birthdate="2004-12-25" gender="M" nation="POL" license="100905700242" swrid="4971377" athleteid="2594">
              <RESULTS>
                <RESULT eventid="1212" points="507" reactiontime="+81" swimtime="00:01:02.06" resultid="2595" heatid="4049" lane="3" entrytime="00:01:04.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="533" reactiontime="+76" swimtime="00:09:17.48" resultid="2596" heatid="4097" lane="1" entrytime="00:09:42.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="100" swimtime="00:01:02.96" />
                    <SPLIT distance="150" swimtime="00:01:36.51" />
                    <SPLIT distance="200" swimtime="00:02:10.95" />
                    <SPLIT distance="250" swimtime="00:02:45.98" />
                    <SPLIT distance="300" swimtime="00:03:21.43" />
                    <SPLIT distance="350" swimtime="00:03:57.16" />
                    <SPLIT distance="400" swimtime="00:04:33.14" />
                    <SPLIT distance="450" swimtime="00:05:09.05" />
                    <SPLIT distance="500" swimtime="00:05:45.12" />
                    <SPLIT distance="550" swimtime="00:06:20.85" />
                    <SPLIT distance="600" swimtime="00:06:56.80" />
                    <SPLIT distance="650" swimtime="00:07:32.41" />
                    <SPLIT distance="700" swimtime="00:08:07.94" />
                    <SPLIT distance="750" swimtime="00:08:43.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="527" reactiontime="+73" swimtime="00:00:58.04" resultid="2597" heatid="4113" lane="3" entrytime="00:01:00.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="474" reactiontime="+83" swimtime="00:02:21.94" resultid="2598" heatid="4125" lane="9" entrytime="00:02:24.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="100" swimtime="00:01:06.95" />
                    <SPLIT distance="150" swimtime="00:01:44.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Barański" birthdate="2007-09-12" gender="M" nation="POL" license="100905700377" swrid="5225103" athleteid="2542">
              <RESULTS>
                <RESULT eventid="1166" points="353" reactiontime="+73" swimtime="00:00:36.71" resultid="2543" heatid="4042" lane="0" entrytime="00:00:35.92" entrycourse="LCM" />
                <RESULT eventid="1350" points="324" reactiontime="+69" swimtime="00:01:22.74" resultid="2544" heatid="4080" lane="8" entrytime="00:01:20.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="346" reactiontime="+69" swimtime="00:01:06.80" resultid="2545" heatid="4111" lane="4" entrytime="00:01:07.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Furmaniak" birthdate="2006-04-04" gender="F" nation="POL" license="100905600490" swrid="5190496" athleteid="2605">
              <RESULTS>
                <RESULT eventid="1235" points="520" reactiontime="+66" swimtime="00:00:33.54" resultid="2606" heatid="4055" lane="0" entrytime="00:00:33.16" entrycourse="LCM" />
                <RESULT eventid="1281" points="483" reactiontime="+80" swimtime="00:02:23.99" resultid="2607" heatid="4061" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:09.76" />
                    <SPLIT distance="150" swimtime="00:01:47.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="386" reactiontime="+76" swimtime="00:00:33.55" resultid="2608" heatid="4087" lane="2" entrytime="00:00:32.67" entrycourse="LCM" />
                <RESULT eventid="1451" points="505" reactiontime="+83" swimtime="00:01:04.91" resultid="2609" heatid="4103" lane="0" entrytime="00:01:06.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="457" reactiontime="+60" swimtime="00:01:14.73" resultid="2610" heatid="4130" lane="8" entrytime="00:01:12.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sandra" lastname="Jawor" birthdate="2005-06-05" gender="F" nation="POL" license="100905600294" swrid="5190449" athleteid="2518">
              <RESULTS>
                <RESULT eventid="1143" points="364" reactiontime="+78" swimtime="00:00:41.14" resultid="2519" heatid="4036" lane="9" entrytime="00:00:41.93" entrycourse="LCM" />
                <RESULT eventid="1281" points="462" reactiontime="+79" swimtime="00:02:26.10" resultid="2520" heatid="4063" lane="5" entrytime="00:02:28.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="150" swimtime="00:01:49.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="425" reactiontime="+82" swimtime="00:01:08.75" resultid="2521" heatid="4102" lane="5" entrytime="00:01:07.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Kowacka" birthdate="2004-10-03" gender="F" nation="POL" license="100905600434" swrid="5088808" athleteid="2622">
              <RESULTS>
                <RESULT eventid="1281" points="531" reactiontime="+72" swimtime="00:02:19.45" resultid="2623" heatid="4065" lane="8" entrytime="00:02:18.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:06.90" />
                    <SPLIT distance="150" swimtime="00:01:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="409" reactiontime="+67" swimtime="00:00:32.90" resultid="2624" heatid="4087" lane="7" entrytime="00:00:32.68" entrycourse="LCM" />
                <RESULT eventid="1451" points="506" reactiontime="+76" swimtime="00:01:04.87" resultid="2625" heatid="4104" lane="1" entrytime="00:01:04.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="484" reactiontime="+73" swimtime="00:02:40.56" resultid="2626" heatid="4137" lane="3" entrytime="00:02:40.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:02:04.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matylda" lastname="Barańska" birthdate="2006-02-10" gender="F" nation="POL" license="100905600376" swrid="5195529" athleteid="2514">
              <RESULTS>
                <RESULT eventid="1143" points="397" reactiontime="+86" swimtime="00:00:39.97" resultid="2515" heatid="4036" lane="6" entrytime="00:00:39.11" entrycourse="LCM" />
                <RESULT eventid="1327" points="360" reactiontime="+82" swimtime="00:01:30.11" resultid="2516" heatid="4075" lane="9" entrytime="00:01:29.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="359" reactiontime="+84" swimtime="00:03:15.70" resultid="2517" heatid="4117" lane="5" entrytime="00:03:09.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                    <SPLIT distance="100" swimtime="00:01:35.14" />
                    <SPLIT distance="150" swimtime="00:02:26.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Stanisławski" birthdate="2004-06-12" gender="M" nation="POL" license="100905700425" swrid="4980419" athleteid="2632">
              <RESULTS>
                <RESULT eventid="1304" points="528" reactiontime="+74" swimtime="00:02:06.15" resultid="2633" heatid="4071" lane="6" entrytime="00:02:10.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:01:00.18" />
                    <SPLIT distance="150" swimtime="00:01:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="564" reactiontime="+71" swimtime="00:00:26.95" resultid="2634" heatid="4093" lane="5" entrytime="00:00:27.42" entrycourse="LCM" />
                <RESULT eventid="1475" points="520" reactiontime="+81" swimtime="00:00:58.30" resultid="2635" heatid="4114" lane="0" entrytime="00:00:58.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="474" reactiontime="+71" swimtime="00:02:23.45" resultid="2636" heatid="4155" lane="1" entrytime="00:02:19.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:07.49" />
                    <SPLIT distance="150" swimtime="00:01:45.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Czyżak" birthdate="2009-09-23" gender="M" nation="POL" license="100905700438" swrid="5398856" athleteid="2554">
              <RESULTS>
                <RESULT eventid="1166" points="215" reactiontime="+62" swimtime="00:00:43.26" resultid="2555" heatid="4040" lane="1" entrytime="00:00:44.84" entrycourse="LCM" />
                <RESULT eventid="1350" points="228" reactiontime="+72" swimtime="00:01:33.09" resultid="2556" heatid="4078" lane="4" entrytime="00:01:37.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="258" reactiontime="+64" swimtime="00:03:17.88" resultid="2557" heatid="4120" lane="6" entrytime="00:03:24.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                    <SPLIT distance="100" swimtime="00:01:35.02" />
                    <SPLIT distance="150" swimtime="00:02:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="237" reactiontime="+69" swimtime="00:03:00.79" resultid="2558" heatid="4153" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:29.39" />
                    <SPLIT distance="150" swimtime="00:02:15.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Zajączkowska" birthdate="2004-08-25" gender="F" nation="POL" license="100905600372" swrid="5034878" athleteid="2572">
              <RESULTS>
                <RESULT eventid="1189" points="550" reactiontime="+75" swimtime="00:01:07.70" resultid="2573" heatid="4046" lane="8" entrytime="00:01:08.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="563" reactiontime="+65" swimtime="00:00:32.66" resultid="2574" heatid="4055" lane="7" entrytime="00:00:32.61" entrycourse="LCM" />
                <RESULT eventid="1373" points="464" reactiontime="+78" swimtime="00:00:31.55" resultid="2575" heatid="4083" lane="6" />
                <RESULT eventid="1451" points="536" reactiontime="+78" swimtime="00:01:03.65" resultid="2576" heatid="4104" lane="7" entrytime="00:01:04.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="557" reactiontime="+62" swimtime="00:02:29.89" resultid="2577" heatid="4152" lane="2" entrytime="00:02:29.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                    <SPLIT distance="150" swimtime="00:01:51.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Węgrzycka" birthdate="2008-08-20" gender="F" nation="POL" license="100905600383" swrid="5096198" athleteid="2526">
              <RESULTS>
                <RESULT eventid="1143" points="335" reactiontime="+96" swimtime="00:00:42.31" resultid="2527" heatid="4035" lane="6" entrytime="00:00:43.07" entrycourse="LCM" />
                <RESULT eventid="1189" points="310" swimtime="00:01:21.90" resultid="2528" heatid="4045" lane="0" entrytime="00:01:22.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="318" reactiontime="+98" swimtime="00:00:35.77" resultid="2529" heatid="4085" lane="4" entrytime="00:00:36.31" entrycourse="LCM" />
                <RESULT eventid="1451" points="360" reactiontime="+97" swimtime="00:01:12.65" resultid="2530" heatid="4101" lane="1" entrytime="00:01:19.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="318" reactiontime="+89" swimtime="00:05:46.29" resultid="2531" heatid="4144" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:19.97" />
                    <SPLIT distance="150" swimtime="00:02:05.27" />
                    <SPLIT distance="200" swimtime="00:02:50.22" />
                    <SPLIT distance="250" swimtime="00:03:35.71" />
                    <SPLIT distance="300" swimtime="00:04:20.42" />
                    <SPLIT distance="350" swimtime="00:05:04.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Królewski" birthdate="2008-09-20" gender="M" nation="POL" license="100905700381" swrid="5096077" athleteid="2499">
              <RESULTS>
                <RESULT eventid="1120" points="163" reactiontime="+68" swimtime="00:00:38.22" resultid="2500" heatid="4026" lane="2" entrytime="00:00:37.86" entrycourse="LCM" />
                <RESULT eventid="1258" points="153" reactiontime="+69" swimtime="00:00:44.85" resultid="2501" heatid="4057" lane="6" entrytime="00:00:45.20" entrycourse="LCM" />
                <RESULT eventid="1475" points="178" swimtime="00:01:23.39" resultid="2502" heatid="4109" lane="5" entrytime="00:01:24.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="161" reactiontime="+76" swimtime="00:01:35.25" resultid="2503" heatid="4134" lane="0" entrytime="00:01:37.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Cichacz" birthdate="2009-02-09" gender="M" nation="POL" license="100905700407" swrid="4976851" athleteid="2477">
              <RESULTS>
                <RESULT eventid="1120" points="114" reactiontime="+65" swimtime="00:00:43.01" resultid="2478" heatid="4026" lane="7" entrytime="00:00:41.59" entrycourse="LCM" />
                <RESULT comment="M4 - Pływak wykonał nierównoczesne ruchy ramion." eventid="1396" reactiontime="+76" status="DSQ" swimtime="00:00:57.87" resultid="2479" heatid="4090" lane="7" />
                <RESULT eventid="1475" points="110" reactiontime="+89" swimtime="00:01:37.74" resultid="2480" heatid="4109" lane="1" entrytime="00:01:41.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M4 - Pływak wykonał nierównoczesne ruchy ramion." eventid="1659" status="DSQ" swimtime="00:04:19.80" resultid="2481" heatid="4139" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:02.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Samulczyk" birthdate="2009-03-29" gender="F" nation="POL" license="100905600416" swrid="4976893" athleteid="2444">
              <RESULTS>
                <RESULT eventid="1070" status="DNS" swimtime="00:00:00.00" resultid="2445" heatid="4014" lane="3" />
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="2446" heatid="4052" lane="0" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1451" reactiontime="+62" status="DSQ" swimtime="00:01:23.37" resultid="2447" heatid="4099" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="200" swimtime="00:01:38.41" resultid="2448" heatid="4126" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivier" lastname="Urbaniak" birthdate="2007-06-01" gender="M" nation="POL" license="100905700356" swrid="5197965" athleteid="2464">
              <RESULTS>
                <RESULT eventid="1120" points="427" reactiontime="+81" swimtime="00:00:27.75" resultid="2465" heatid="4030" lane="0" entrytime="00:00:28.88" entrycourse="LCM" />
                <RESULT eventid="1212" points="429" reactiontime="+75" swimtime="00:01:05.63" resultid="2466" heatid="4049" lane="7" entrytime="00:01:06.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="499" reactiontime="+71" swimtime="00:00:30.25" resultid="2467" heatid="4060" lane="8" entrytime="00:00:29.53" entrycourse="LCM" />
                <RESULT eventid="1613" points="534" reactiontime="+66" swimtime="00:01:03.89" resultid="2468" heatid="4136" lane="4" entrytime="00:01:01.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="481" reactiontime="+73" swimtime="00:02:25.45" resultid="2469" heatid="4142" lane="7" entrytime="00:02:23.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:09.17" />
                    <SPLIT distance="150" swimtime="00:01:53.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="525" reactiontime="+68" swimtime="00:02:18.71" resultid="2470" heatid="4155" lane="3" entrytime="00:02:14.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:08.58" />
                    <SPLIT distance="150" swimtime="00:01:45.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Mikołajewski" birthdate="2009-03-06" gender="M" nation="POL" license="100905700418" swrid="5260894" athleteid="2567">
              <RESULTS>
                <RESULT eventid="1166" points="136" swimtime="00:00:50.43" resultid="2568" heatid="4039" lane="5" entrytime="00:00:48.80" entrycourse="LCM" />
                <RESULT eventid="1350" points="129" swimtime="00:01:52.45" resultid="2569" heatid="4078" lane="6" entrytime="00:01:44.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="124" swimtime="00:01:33.90" resultid="2570" heatid="4109" lane="2" entrytime="00:01:34.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="104" reactiontime="+87" swimtime="00:01:49.94" resultid="2571" heatid="4133" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01610" nation="POL" region="10" clubid="2067" name="Grupa Pływacka Gdynia Masters">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Skwarło" birthdate="1939-05-03" gender="M" nation="POL" license="501610700017" swrid="4302086" athleteid="2068">
              <RESULTS>
                <RESULT eventid="1166" points="102" swimtime="00:00:55.42" resultid="2069" heatid="4038" lane="4" />
                <RESULT eventid="1258" points="54" reactiontime="+94" swimtime="00:01:03.30" resultid="2070" heatid="4057" lane="9" />
                <RESULT eventid="1521" points="80" swimtime="00:04:52.26" resultid="2071" heatid="4120" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.08" />
                    <SPLIT distance="100" swimtime="00:02:20.69" />
                    <SPLIT distance="150" swimtime="00:03:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="42" reactiontime="+95" swimtime="00:02:28.07" resultid="2072" heatid="4132" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="3695" name="Warsaw Masters Team">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Grochowski" birthdate="1991-08-29" gender="M" nation="POL" license="504214700106" athleteid="3696">
              <RESULTS>
                <RESULT eventid="1304" points="302" reactiontime="+79" swimtime="00:02:32.02" resultid="3697" heatid="4067" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="307" reactiontime="+78" swimtime="00:05:26.16" resultid="3698" heatid="4146" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:16.26" />
                    <SPLIT distance="150" swimtime="00:01:57.40" />
                    <SPLIT distance="200" swimtime="00:02:38.80" />
                    <SPLIT distance="250" swimtime="00:03:20.41" />
                    <SPLIT distance="300" swimtime="00:04:02.88" />
                    <SPLIT distance="350" swimtime="00:04:45.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04115" nation="POL" region="15" clubid="2193" name="KTP Iskra Konin">
          <ATHLETES>
            <ATHLETE firstname="Alan" lastname="Bidziński" birthdate="2006-06-28" gender="M" nation="POL" license="104115700040" swrid="5190174" athleteid="2211">
              <RESULTS>
                <RESULT eventid="1120" points="511" reactiontime="+71" swimtime="00:00:26.14" resultid="2212" heatid="4024" lane="7" />
                <RESULT eventid="1258" points="425" reactiontime="+77" swimtime="00:00:31.91" resultid="2213" heatid="4056" lane="1" />
                <RESULT eventid="1304" points="415" reactiontime="+77" swimtime="00:02:16.64" resultid="2214" heatid="4068" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:05.28" />
                    <SPLIT distance="150" swimtime="00:01:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="538" reactiontime="+75" swimtime="00:00:57.66" resultid="2215" heatid="4108" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Janiak" birthdate="2006-02-26" gender="F" nation="POL" license="104115600068" swrid="5197714" athleteid="2205">
              <RESULTS>
                <RESULT eventid="1070" points="488" reactiontime="+75" swimtime="00:00:30.05" resultid="2206" heatid="4015" lane="2" />
                <RESULT eventid="1143" points="407" reactiontime="+72" swimtime="00:00:39.66" resultid="2207" heatid="4033" lane="3" />
                <RESULT eventid="1327" points="412" reactiontime="+73" swimtime="00:01:26.14" resultid="2208" heatid="4073" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="354" reactiontime="+75" swimtime="00:00:34.53" resultid="2209" heatid="4084" lane="2" />
                <RESULT eventid="1451" points="458" reactiontime="+75" swimtime="00:01:07.08" resultid="2210" heatid="4098" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Chestkowska" birthdate="2006-10-01" gender="F" nation="POL" license="104115600047" swrid="5249565" athleteid="2200">
              <RESULTS>
                <RESULT eventid="1070" points="286" reactiontime="+85" swimtime="00:00:35.91" resultid="2201" heatid="4016" lane="0" />
                <RESULT eventid="1143" points="299" reactiontime="+77" swimtime="00:00:43.94" resultid="2202" heatid="4034" lane="2" />
                <RESULT eventid="1327" points="302" reactiontime="+78" swimtime="00:01:35.49" resultid="2203" heatid="4073" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="257" reactiontime="+68" swimtime="00:01:21.32" resultid="2204" heatid="4098" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Klaudia" lastname="Borkiewicz" birthdate="2006-07-21" gender="F" nation="POL" license="104115600034" swrid="5009625" athleteid="2194">
              <RESULTS>
                <RESULT eventid="1070" points="580" reactiontime="+70" swimtime="00:00:28.38" resultid="2195" heatid="4014" lane="5" />
                <RESULT eventid="1235" points="602" reactiontime="+65" swimtime="00:00:31.94" resultid="2196" heatid="4051" lane="7" />
                <RESULT eventid="1373" points="537" reactiontime="+75" swimtime="00:00:30.04" resultid="2197" heatid="4082" lane="3" />
                <RESULT eventid="1451" points="508" reactiontime="+68" swimtime="00:01:04.77" resultid="2198" heatid="4099" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="502" reactiontime="+66" swimtime="00:01:12.43" resultid="2199" heatid="4127" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00414" nation="POL" region="14" clubid="2023" name="Buks">
          <ATHLETES>
            <ATHLETE firstname="Szymon" lastname="Berner" birthdate="2004-06-09" gender="M" nation="POL" license="100414700261" swrid="4011653" athleteid="2024">
              <RESULTS>
                <RESULT eventid="1120" points="592" reactiontime="+72" swimtime="00:00:24.90" resultid="2025" heatid="4032" lane="7" entrytime="00:00:24.89" entrycourse="LCM" />
                <RESULT eventid="1258" points="572" reactiontime="+63" swimtime="00:00:28.91" resultid="2026" heatid="4060" lane="9" entrytime="00:00:29.73" entrycourse="LCM" />
                <RESULT eventid="1396" points="557" reactiontime="+65" swimtime="00:00:27.06" resultid="2027" heatid="4094" lane="9" entrytime="00:00:27.36" entrycourse="LCM" />
                <RESULT eventid="1475" points="606" reactiontime="+75" swimtime="00:00:55.42" resultid="2028" heatid="4115" lane="0" entrytime="00:00:54.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="519" reactiontime="+61" swimtime="00:01:04.51" resultid="2029" heatid="4133" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02305" nation="POL" region="05" clubid="2017" name="AZS Łódź">
          <ATHLETES>
            <ATHLETE firstname="Wiktoria" lastname="Raczyńska" birthdate="2004-04-16" gender="F" nation="POL" license="102305600064" swrid="5034876" athleteid="2018">
              <RESULTS>
                <RESULT eventid="1070" points="503" reactiontime="+66" swimtime="00:00:29.76" resultid="2019" heatid="4016" lane="9" />
                <RESULT eventid="1189" points="552" reactiontime="+71" swimtime="00:01:07.61" resultid="2020" heatid="4046" lane="2" entrytime="00:01:07.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="540" reactiontime="+67" swimtime="00:00:30.00" resultid="2021" heatid="4088" lane="6" entrytime="00:00:29.82" entrycourse="LCM" />
                <RESULT eventid="1451" points="568" reactiontime="+67" swimtime="00:01:02.42" resultid="2022" heatid="4105" lane="3" entrytime="00:01:02.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01605" nation="POL" region="05" clubid="3104" name="UKS 190 Łódź">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Nieckarz" birthdate="2006-04-06" gender="M" nation="POL" license="101605700184" swrid="5195522" athleteid="3260">
              <RESULTS>
                <RESULT eventid="1166" points="377" reactiontime="+70" swimtime="00:00:35.91" resultid="3261" heatid="4042" lane="6" entrytime="00:00:34.80" entrycourse="LCM" />
                <RESULT eventid="1350" points="401" reactiontime="+78" swimtime="00:01:17.11" resultid="3262" heatid="4080" lane="4" entrytime="00:01:16.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="450" reactiontime="+84" swimtime="00:02:44.51" resultid="3263" heatid="4122" lane="1" entrytime="00:02:43.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:18.57" />
                    <SPLIT distance="150" swimtime="00:02:01.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="429" reactiontime="+76" swimtime="00:02:31.14" resultid="3264" heatid="4139" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="100" swimtime="00:01:13.09" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Janiszewski" birthdate="2006-05-17" gender="M" nation="POL" license="101605700331" swrid="5025340" athleteid="3280">
              <RESULTS>
                <RESULT eventid="1212" points="537" reactiontime="+66" swimtime="00:01:00.89" resultid="3281" heatid="4050" lane="7" entrytime="00:01:00.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="523" reactiontime="+59" swimtime="00:00:27.64" resultid="3282" heatid="4093" lane="4" entrytime="00:00:27.37" entrycourse="LCM" />
                <RESULT eventid="1567" points="509" reactiontime="+67" swimtime="00:02:18.67" resultid="3283" heatid="4125" lane="7" entrytime="00:02:16.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:43.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="483" reactiontime="+63" swimtime="00:02:25.21" resultid="3284" heatid="4139" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                    <SPLIT distance="100" swimtime="00:01:09.14" />
                    <SPLIT distance="150" swimtime="00:01:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="508" reactiontime="+71" swimtime="00:04:35.72" resultid="3285" heatid="4148" lane="3" entrytime="00:04:48.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:46.43" />
                    <SPLIT distance="200" swimtime="00:02:23.25" />
                    <SPLIT distance="250" swimtime="00:02:58.81" />
                    <SPLIT distance="300" swimtime="00:03:34.91" />
                    <SPLIT distance="350" swimtime="00:04:06.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Pawlak" birthdate="2008-08-20" gender="M" nation="POL" license="101605700228" swrid="5249645" athleteid="3270">
              <RESULTS>
                <RESULT eventid="1212" points="257" reactiontime="+90" swimtime="00:01:17.76" resultid="3271" heatid="4048" lane="2" entrytime="00:01:17.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="245" swimtime="00:01:30.81" resultid="3272" heatid="4079" lane="2" entrytime="00:01:30.09" entrycourse="LCM" />
                <RESULT eventid="1521" points="292" reactiontime="+78" swimtime="00:03:09.95" resultid="3273" heatid="4120" lane="3" entrytime="00:03:13.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.34" />
                    <SPLIT distance="100" swimtime="00:01:34.40" />
                    <SPLIT distance="150" swimtime="00:02:22.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="320" reactiontime="+91" swimtime="00:02:46.59" resultid="3274" heatid="4141" lane="1" entrytime="00:02:49.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:01:22.83" />
                    <SPLIT distance="150" swimtime="00:02:10.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roksana" lastname="Wodecka" birthdate="2003-02-20" gender="F" nation="POL" license="101605600249" swrid="4896414" athleteid="3292">
              <RESULTS>
                <RESULT eventid="1451" points="542" reactiontime="+68" swimtime="00:01:03.41" resultid="3293" heatid="4105" lane="7" entrytime="00:01:02.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="529" reactiontime="+61" swimtime="00:01:11.17" resultid="3294" heatid="4130" lane="2" entrytime="00:01:09.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="494" reactiontime="+62" swimtime="00:02:35.94" resultid="3295" heatid="4152" lane="6" entrytime="00:02:29.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="150" swimtime="00:01:57.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Kobus" birthdate="2005-02-01" gender="M" nation="POL" license="101605700268" swrid="5113373" athleteid="3250">
              <RESULTS>
                <RESULT eventid="1166" points="579" reactiontime="+62" swimtime="00:00:31.13" resultid="3251" heatid="4043" lane="3" entrytime="00:00:31.34" entrycourse="LCM" />
                <RESULT eventid="1350" points="585" reactiontime="+61" swimtime="00:01:08.00" resultid="3252" heatid="4081" lane="5" entrytime="00:01:07.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="628" reactiontime="+62" swimtime="00:02:27.27" resultid="3253" heatid="4122" lane="4" entrytime="00:02:24.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:10.31" />
                    <SPLIT distance="150" swimtime="00:01:49.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="502" reactiontime="+66" swimtime="00:02:23.35" resultid="3254" heatid="4142" lane="1" entrytime="00:02:24.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:49.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ignacy" lastname="Trudnos" birthdate="2008-02-13" gender="M" nation="POL" license="101605700221" swrid="5269112" athleteid="3244">
              <RESULTS>
                <RESULT eventid="1166" points="333" reactiontime="+74" swimtime="00:00:37.41" resultid="3245" heatid="4041" lane="9" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1350" points="339" reactiontime="+79" swimtime="00:01:21.53" resultid="3246" heatid="4080" lane="1" entrytime="00:01:20.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="382" reactiontime="+65" swimtime="00:02:53.78" resultid="3247" heatid="4121" lane="5" entrytime="00:02:52.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                    <SPLIT distance="100" swimtime="00:01:24.35" />
                    <SPLIT distance="150" swimtime="00:02:09.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="371" reactiontime="+70" swimtime="00:02:38.55" resultid="3248" heatid="4141" lane="5" entrytime="00:02:38.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:02:01.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="356" reactiontime="+74" swimtime="00:02:37.78" resultid="3249" heatid="4154" lane="5" entrytime="00:02:38.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="150" swimtime="00:01:58.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Gomułka" birthdate="2006-05-17" gender="F" nation="POL" license="101605600182" swrid="5170204" athleteid="3118">
              <RESULTS>
                <RESULT eventid="1060" points="581" reactiontime="+77" swimtime="00:05:19.15" resultid="3119" heatid="4011" lane="5" entrytime="00:05:14.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:54.36" />
                    <SPLIT distance="200" swimtime="00:02:34.40" />
                    <SPLIT distance="250" swimtime="00:03:19.86" />
                    <SPLIT distance="300" swimtime="00:04:05.95" />
                    <SPLIT distance="350" swimtime="00:04:42.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="578" reactiontime="+79" swimtime="00:02:15.61" resultid="3120" heatid="4065" lane="6" entrytime="00:02:15.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:06.71" />
                    <SPLIT distance="150" swimtime="00:01:41.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="497" reactiontime="+75" swimtime="00:00:30.84" resultid="3121" heatid="4083" lane="5" />
                <RESULT eventid="1498" points="495" reactiontime="+76" swimtime="00:02:55.81" resultid="3122" heatid="4118" lane="6" entrytime="00:02:55.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:24.90" />
                    <SPLIT distance="150" swimtime="00:02:10.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="609" reactiontime="+77" swimtime="00:02:28.76" resultid="3123" heatid="4138" lane="3" entrytime="00:02:29.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:01:54.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="612" reactiontime="+77" swimtime="00:02:25.28" resultid="3124" heatid="4152" lane="5" entrytime="00:02:26.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:48.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabian" lastname="Janiszewski" birthdate="2009-01-24" gender="M" nation="POL" license="101605700234" swrid="4976858" athleteid="3188">
              <RESULTS>
                <RESULT eventid="1120" points="260" reactiontime="+87" swimtime="00:00:32.75" resultid="3189" heatid="4028" lane="9" entrytime="00:00:32.45" entrycourse="LCM" />
                <RESULT eventid="1166" status="DNS" swimtime="00:00:00.00" resultid="3190" heatid="4038" lane="1" />
                <RESULT eventid="1396" points="211" reactiontime="+96" swimtime="00:00:37.35" resultid="3191" heatid="4091" lane="6" entrytime="00:00:36.86" entrycourse="LCM" />
                <RESULT eventid="1475" points="289" swimtime="00:01:10.89" resultid="3192" heatid="4111" lane="0" entrytime="00:01:10.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="286" reactiontime="+76" swimtime="00:01:18.61" resultid="3193" heatid="4134" lane="6" entrytime="00:01:23.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Walkowski" birthdate="2007-12-11" gender="M" nation="POL" license="101605700215" swrid="5254768" athleteid="3144">
              <RESULTS>
                <RESULT eventid="1065" points="489" reactiontime="+68" swimtime="00:05:09.49" resultid="3145" heatid="4013" lane="1" entrytime="00:05:06.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:09.12" />
                    <SPLIT distance="150" swimtime="00:01:50.39" />
                    <SPLIT distance="200" swimtime="00:02:29.60" />
                    <SPLIT distance="250" swimtime="00:03:14.48" />
                    <SPLIT distance="300" swimtime="00:04:00.53" />
                    <SPLIT distance="350" swimtime="00:04:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="453" reactiontime="+61" swimtime="00:02:12.72" resultid="3146" heatid="4071" lane="7" entrytime="00:02:11.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:05.90" />
                    <SPLIT distance="150" swimtime="00:01:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="532" reactiontime="+69" swimtime="00:09:17.94" resultid="3147" heatid="4097" lane="7" entrytime="00:09:19.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:07.45" />
                    <SPLIT distance="150" swimtime="00:01:42.58" />
                    <SPLIT distance="200" swimtime="00:02:18.18" />
                    <SPLIT distance="250" swimtime="00:02:53.56" />
                    <SPLIT distance="300" swimtime="00:03:28.59" />
                    <SPLIT distance="350" swimtime="00:04:03.83" />
                    <SPLIT distance="400" swimtime="00:04:39.12" />
                    <SPLIT distance="450" swimtime="00:05:14.17" />
                    <SPLIT distance="500" swimtime="00:05:49.86" />
                    <SPLIT distance="550" swimtime="00:06:25.03" />
                    <SPLIT distance="600" swimtime="00:07:00.35" />
                    <SPLIT distance="650" swimtime="00:07:35.18" />
                    <SPLIT distance="700" swimtime="00:08:10.53" />
                    <SPLIT distance="750" swimtime="00:08:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="429" reactiontime="+69" swimtime="00:02:26.71" resultid="3148" heatid="4124" lane="5" entrytime="00:02:25.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:11.04" />
                    <SPLIT distance="150" swimtime="00:01:49.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="461" reactiontime="+70" swimtime="00:02:27.56" resultid="3149" heatid="4142" lane="0" entrytime="00:02:26.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:12.22" />
                    <SPLIT distance="150" swimtime="00:01:54.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="566" reactiontime="+76" swimtime="00:17:32.71" resultid="3150" heatid="4159" lane="2" entrytime="00:17:49.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.03" />
                    <SPLIT distance="150" swimtime="00:01:42.27" />
                    <SPLIT distance="200" swimtime="00:02:17.73" />
                    <SPLIT distance="250" swimtime="00:02:52.81" />
                    <SPLIT distance="300" swimtime="00:03:27.86" />
                    <SPLIT distance="350" swimtime="00:04:03.14" />
                    <SPLIT distance="400" swimtime="00:04:38.25" />
                    <SPLIT distance="450" swimtime="00:05:13.34" />
                    <SPLIT distance="500" swimtime="00:05:48.16" />
                    <SPLIT distance="550" swimtime="00:06:23.22" />
                    <SPLIT distance="600" swimtime="00:06:58.29" />
                    <SPLIT distance="650" swimtime="00:07:33.47" />
                    <SPLIT distance="700" swimtime="00:08:08.96" />
                    <SPLIT distance="750" swimtime="00:08:44.29" />
                    <SPLIT distance="800" swimtime="00:09:19.56" />
                    <SPLIT distance="850" swimtime="00:09:55.07" />
                    <SPLIT distance="900" swimtime="00:10:30.62" />
                    <SPLIT distance="950" swimtime="00:11:06.25" />
                    <SPLIT distance="1000" swimtime="00:11:41.92" />
                    <SPLIT distance="1050" swimtime="00:12:17.46" />
                    <SPLIT distance="1100" swimtime="00:12:52.98" />
                    <SPLIT distance="1150" swimtime="00:13:28.62" />
                    <SPLIT distance="1200" swimtime="00:14:04.12" />
                    <SPLIT distance="1250" swimtime="00:14:39.42" />
                    <SPLIT distance="1300" swimtime="00:15:14.94" />
                    <SPLIT distance="1350" swimtime="00:15:49.94" />
                    <SPLIT distance="1400" swimtime="00:16:25.31" />
                    <SPLIT distance="1450" swimtime="00:16:59.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Cierpiał" birthdate="2004-12-08" gender="M" nation="POL" license="101605700247" swrid="5038593" athleteid="3255">
              <RESULTS>
                <RESULT eventid="1166" points="422" reactiontime="+67" swimtime="00:00:34.57" resultid="3256" heatid="4043" lane="8" entrytime="00:00:33.36" entrycourse="LCM" />
                <RESULT eventid="1350" points="447" reactiontime="+70" swimtime="00:01:14.37" resultid="3257" heatid="4081" lane="1" entrytime="00:01:13.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="502" reactiontime="+72" swimtime="00:02:38.60" resultid="3258" heatid="4122" lane="2" entrytime="00:02:34.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                    <SPLIT distance="100" swimtime="00:01:18.91" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="433" reactiontime="+67" swimtime="00:02:30.67" resultid="3259" heatid="4142" lane="8" entrytime="00:02:25.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:54.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ignacy" lastname="Czajka" birthdate="2009-12-23" gender="M" nation="POL" license="101605700250" swrid="5398851" athleteid="3177">
              <RESULTS>
                <RESULT eventid="1120" points="119" swimtime="00:00:42.45" resultid="3178" heatid="4026" lane="8" entrytime="00:00:43.08" entrycourse="LCM" />
                <RESULT eventid="1304" points="127" reactiontime="+85" swimtime="00:03:22.78" resultid="3179" heatid="4068" lane="6" entrytime="00:03:47.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.14" />
                    <SPLIT distance="100" swimtime="00:01:36.85" />
                    <SPLIT distance="150" swimtime="00:02:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="115" reactiontime="+99" swimtime="00:01:36.37" resultid="3180" heatid="4109" lane="7" entrytime="00:01:35.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="97" swimtime="00:01:52.48" resultid="3181" heatid="4133" lane="4" entrytime="00:01:51.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Skrobisz" birthdate="2007-06-15" gender="M" nation="POL" license="101605700212" swrid="5198004" athleteid="3265">
              <RESULTS>
                <RESULT eventid="1166" points="435" reactiontime="+85" swimtime="00:00:34.23" resultid="3266" heatid="4042" lane="4" entrytime="00:00:34.10" entrycourse="LCM" />
                <RESULT eventid="1350" points="428" reactiontime="+86" swimtime="00:01:15.45" resultid="3267" heatid="4081" lane="0" entrytime="00:01:14.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="436" reactiontime="+82" swimtime="00:02:46.32" resultid="3268" heatid="4121" lane="4" entrytime="00:02:45.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:21.15" />
                    <SPLIT distance="150" swimtime="00:02:04.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="340" reactiontime="+91" swimtime="00:02:43.29" resultid="3269" heatid="4141" lane="2" entrytime="00:02:48.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="150" swimtime="00:02:04.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Zieliński" birthdate="2003-04-13" gender="M" nation="POL" license="101605700161" swrid="4933033" athleteid="3200">
              <RESULTS>
                <RESULT eventid="1120" points="643" reactiontime="+63" swimtime="00:00:24.22" resultid="3201" heatid="4032" lane="6" entrytime="00:00:24.52" entrycourse="LCM" />
                <RESULT eventid="1304" points="621" reactiontime="+64" swimtime="00:01:59.52" resultid="3202" heatid="4072" lane="5" entrytime="00:01:55.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.07" />
                    <SPLIT distance="100" swimtime="00:00:56.63" />
                    <SPLIT distance="150" swimtime="00:01:27.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="652" reactiontime="+68" swimtime="00:08:41.22" resultid="3203" heatid="4096" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="100" swimtime="00:01:03.77" />
                    <SPLIT distance="150" swimtime="00:01:37.10" />
                    <SPLIT distance="200" swimtime="00:02:10.30" />
                    <SPLIT distance="250" swimtime="00:02:43.54" />
                    <SPLIT distance="300" swimtime="00:03:16.94" />
                    <SPLIT distance="350" swimtime="00:03:50.13" />
                    <SPLIT distance="400" swimtime="00:04:23.39" />
                    <SPLIT distance="450" swimtime="00:04:56.27" />
                    <SPLIT distance="500" swimtime="00:05:29.27" />
                    <SPLIT distance="550" swimtime="00:06:02.18" />
                    <SPLIT distance="600" swimtime="00:06:35.27" />
                    <SPLIT distance="650" swimtime="00:07:07.84" />
                    <SPLIT distance="700" swimtime="00:07:40.15" />
                    <SPLIT distance="750" swimtime="00:08:11.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="679" reactiontime="+68" swimtime="00:00:53.35" resultid="3204" heatid="4115" lane="1" entrytime="00:00:53.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="652" reactiontime="+65" swimtime="00:04:13.75" resultid="3205" heatid="4149" lane="5" entrytime="00:04:09.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                    <SPLIT distance="100" swimtime="00:00:59.42" />
                    <SPLIT distance="150" swimtime="00:01:31.08" />
                    <SPLIT distance="200" swimtime="00:02:03.45" />
                    <SPLIT distance="250" swimtime="00:02:36.57" />
                    <SPLIT distance="300" swimtime="00:03:09.06" />
                    <SPLIT distance="350" swimtime="00:03:41.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Tarczyński" birthdate="2007-04-15" gender="M" nation="POL" license="101605700214" swrid="5198007" athleteid="3137">
              <RESULTS>
                <RESULT eventid="1065" points="517" reactiontime="+83" swimtime="00:05:03.71" resultid="3138" heatid="4013" lane="7" entrytime="00:05:05.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:11.89" />
                    <SPLIT distance="150" swimtime="00:01:53.97" />
                    <SPLIT distance="200" swimtime="00:02:33.20" />
                    <SPLIT distance="250" swimtime="00:03:13.77" />
                    <SPLIT distance="300" swimtime="00:03:55.06" />
                    <SPLIT distance="350" swimtime="00:04:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="430" reactiontime="+82" swimtime="00:00:34.36" resultid="3139" heatid="4043" lane="0" entrytime="00:00:33.56" entrycourse="LCM" />
                <RESULT eventid="1350" points="449" reactiontime="+82" swimtime="00:01:14.25" resultid="3140" heatid="4081" lane="7" entrytime="00:01:12.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="492" reactiontime="+82" swimtime="00:02:39.73" resultid="3141" heatid="4122" lane="6" entrytime="00:02:34.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:18.20" />
                    <SPLIT distance="150" swimtime="00:02:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="477" reactiontime="+80" swimtime="00:02:25.86" resultid="3142" heatid="4142" lane="2" entrytime="00:02:22.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="150" swimtime="00:01:53.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="546" reactiontime="+80" swimtime="00:17:45.47" resultid="3143" heatid="4159" lane="6" entrytime="00:17:42.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:08.48" />
                    <SPLIT distance="150" swimtime="00:01:44.16" />
                    <SPLIT distance="200" swimtime="00:02:19.73" />
                    <SPLIT distance="250" swimtime="00:02:54.81" />
                    <SPLIT distance="300" swimtime="00:03:30.53" />
                    <SPLIT distance="350" swimtime="00:04:06.01" />
                    <SPLIT distance="400" swimtime="00:04:41.51" />
                    <SPLIT distance="450" swimtime="00:05:16.76" />
                    <SPLIT distance="500" swimtime="00:05:52.66" />
                    <SPLIT distance="550" swimtime="00:06:28.09" />
                    <SPLIT distance="600" swimtime="00:07:03.65" />
                    <SPLIT distance="650" swimtime="00:07:39.19" />
                    <SPLIT distance="700" swimtime="00:08:15.09" />
                    <SPLIT distance="750" swimtime="00:08:50.32" />
                    <SPLIT distance="800" swimtime="00:09:26.41" />
                    <SPLIT distance="850" swimtime="00:10:02.00" />
                    <SPLIT distance="900" swimtime="00:10:37.85" />
                    <SPLIT distance="950" swimtime="00:11:13.20" />
                    <SPLIT distance="1000" swimtime="00:11:49.42" />
                    <SPLIT distance="1050" swimtime="00:12:25.37" />
                    <SPLIT distance="1100" swimtime="00:13:01.61" />
                    <SPLIT distance="1150" swimtime="00:13:37.26" />
                    <SPLIT distance="1200" swimtime="00:14:14.05" />
                    <SPLIT distance="1250" swimtime="00:14:49.51" />
                    <SPLIT distance="1300" swimtime="00:15:25.84" />
                    <SPLIT distance="1350" swimtime="00:16:01.37" />
                    <SPLIT distance="1400" swimtime="00:16:37.17" />
                    <SPLIT distance="1450" swimtime="00:17:12.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sergiusz" lastname="Gołacki" birthdate="2004-09-02" gender="M" nation="POL" license="101605700173" swrid="5034812" athleteid="3132">
              <RESULTS>
                <RESULT eventid="1065" points="599" reactiontime="+66" swimtime="00:04:49.15" resultid="3133" heatid="4013" lane="2" entrytime="00:04:59.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                    <SPLIT distance="100" swimtime="00:01:02.11" />
                    <SPLIT distance="150" swimtime="00:01:41.50" />
                    <SPLIT distance="200" swimtime="00:02:19.35" />
                    <SPLIT distance="250" swimtime="00:03:02.31" />
                    <SPLIT distance="300" swimtime="00:03:45.32" />
                    <SPLIT distance="350" swimtime="00:04:17.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="662" reactiontime="+64" swimtime="00:08:38.73" resultid="3134" heatid="4097" lane="4" entrytime="00:08:33.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:01:02.46" />
                    <SPLIT distance="150" swimtime="00:01:34.88" />
                    <SPLIT distance="200" swimtime="00:02:07.58" />
                    <SPLIT distance="250" swimtime="00:04:51.56" />
                    <SPLIT distance="300" swimtime="00:03:13.32" />
                    <SPLIT distance="350" swimtime="00:05:57.43" />
                    <SPLIT distance="400" swimtime="00:04:18.73" />
                    <SPLIT distance="450" swimtime="00:07:02.80" />
                    <SPLIT distance="500" swimtime="00:05:24.66" />
                    <SPLIT distance="550" swimtime="00:08:07.86" />
                    <SPLIT distance="600" swimtime="00:06:30.32" />
                    <SPLIT distance="700" swimtime="00:07:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="645" reactiontime="+60" swimtime="00:02:08.10" resultid="3135" heatid="4125" lane="5" entrytime="00:02:06.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:01.72" />
                    <SPLIT distance="150" swimtime="00:01:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="678" reactiontime="+64" swimtime="00:16:31.46" resultid="3136" heatid="4159" lane="4" entrytime="00:16:12.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.92" />
                    <SPLIT distance="100" swimtime="00:01:02.21" />
                    <SPLIT distance="150" swimtime="00:08:14.32" />
                    <SPLIT distance="200" swimtime="00:02:07.88" />
                    <SPLIT distance="250" swimtime="00:11:34.37" />
                    <SPLIT distance="300" swimtime="00:03:14.34" />
                    <SPLIT distance="350" swimtime="00:12:40.97" />
                    <SPLIT distance="400" swimtime="00:04:20.86" />
                    <SPLIT distance="450" swimtime="00:13:47.47" />
                    <SPLIT distance="500" swimtime="00:05:27.50" />
                    <SPLIT distance="550" swimtime="00:14:54.42" />
                    <SPLIT distance="600" swimtime="00:06:34.15" />
                    <SPLIT distance="650" swimtime="00:15:59.61" />
                    <SPLIT distance="700" swimtime="00:07:40.79" />
                    <SPLIT distance="800" swimtime="00:08:47.85" />
                    <SPLIT distance="900" swimtime="00:09:54.67" />
                    <SPLIT distance="1000" swimtime="00:11:01.13" />
                    <SPLIT distance="1100" swimtime="00:12:07.65" />
                    <SPLIT distance="1200" swimtime="00:13:14.36" />
                    <SPLIT distance="1300" swimtime="00:14:20.95" />
                    <SPLIT distance="1400" swimtime="00:15:27.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Olszyca" birthdate="2009-02-01" gender="M" nation="POL" license="101605700236" swrid="4976741" athleteid="3275">
              <RESULTS>
                <RESULT eventid="1212" points="210" reactiontime="+86" swimtime="00:01:23.24" resultid="3276" heatid="4048" lane="1" entrytime="00:01:21.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="331" reactiontime="+78" swimtime="00:02:27.31" resultid="3277" heatid="4069" lane="4" entrytime="00:02:27.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="150" swimtime="00:01:50.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="365" reactiontime="+70" swimtime="00:05:07.81" resultid="3278" heatid="4147" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="150" swimtime="00:01:54.81" />
                    <SPLIT distance="200" swimtime="00:02:34.05" />
                    <SPLIT distance="250" swimtime="00:03:13.40" />
                    <SPLIT distance="300" swimtime="00:03:52.73" />
                    <SPLIT distance="350" swimtime="00:04:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="263" reactiontime="+79" swimtime="00:02:54.49" resultid="3279" heatid="4154" lane="1" entrytime="00:02:50.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:26.50" />
                    <SPLIT distance="150" swimtime="00:02:11.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Walkowski" birthdate="2007-12-11" gender="M" nation="POL" license="101605700216" swrid="5254775" athleteid="3151">
              <RESULTS>
                <RESULT eventid="1065" points="448" reactiontime="+76" swimtime="00:05:18.66" resultid="3152" heatid="4012" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:10.78" />
                    <SPLIT distance="150" swimtime="00:01:53.36" />
                    <SPLIT distance="200" swimtime="00:02:35.00" />
                    <SPLIT distance="250" swimtime="00:03:21.98" />
                    <SPLIT distance="300" swimtime="00:04:08.79" />
                    <SPLIT distance="350" swimtime="00:04:44.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="431" reactiontime="+75" swimtime="00:01:05.50" resultid="3153" heatid="4049" lane="2" entrytime="00:01:06.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="406" reactiontime="+74" swimtime="00:02:17.70" resultid="3154" heatid="4070" lane="2" entrytime="00:02:17.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:08.37" />
                    <SPLIT distance="150" swimtime="00:01:44.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="462" reactiontime="+78" swimtime="00:02:23.17" resultid="3155" heatid="4124" lane="4" entrytime="00:02:25.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:11.15" />
                    <SPLIT distance="150" swimtime="00:01:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="511" reactiontime="+74" swimtime="00:18:08.80" resultid="3156" heatid="4158" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="150" swimtime="00:01:48.37" />
                    <SPLIT distance="200" swimtime="00:02:25.13" />
                    <SPLIT distance="250" swimtime="00:03:02.05" />
                    <SPLIT distance="300" swimtime="00:03:38.86" />
                    <SPLIT distance="350" swimtime="00:04:15.50" />
                    <SPLIT distance="400" swimtime="00:04:52.04" />
                    <SPLIT distance="450" swimtime="00:05:28.63" />
                    <SPLIT distance="500" swimtime="00:06:05.20" />
                    <SPLIT distance="550" swimtime="00:06:41.92" />
                    <SPLIT distance="600" swimtime="00:07:18.48" />
                    <SPLIT distance="650" swimtime="00:07:55.16" />
                    <SPLIT distance="700" swimtime="00:08:31.58" />
                    <SPLIT distance="750" swimtime="00:09:08.14" />
                    <SPLIT distance="800" swimtime="00:09:44.56" />
                    <SPLIT distance="850" swimtime="00:10:21.23" />
                    <SPLIT distance="900" swimtime="00:10:57.92" />
                    <SPLIT distance="950" swimtime="00:11:34.28" />
                    <SPLIT distance="1000" swimtime="00:12:10.81" />
                    <SPLIT distance="1050" swimtime="00:12:47.15" />
                    <SPLIT distance="1100" swimtime="00:13:23.58" />
                    <SPLIT distance="1150" swimtime="00:14:00.01" />
                    <SPLIT distance="1200" swimtime="00:14:36.28" />
                    <SPLIT distance="1250" swimtime="00:15:12.55" />
                    <SPLIT distance="1300" swimtime="00:15:48.73" />
                    <SPLIT distance="1350" swimtime="00:16:24.72" />
                    <SPLIT distance="1400" swimtime="00:17:00.81" />
                    <SPLIT distance="1450" swimtime="00:17:36.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julita" lastname="Kossowska" birthdate="2005-07-20" gender="F" nation="POL" license="101605600153" swrid="5118469" athleteid="3162">
              <RESULTS>
                <RESULT eventid="1070" points="523" reactiontime="+81" swimtime="00:00:29.36" resultid="3163" heatid="4022" lane="6" entrytime="00:00:28.75" entrycourse="LCM" />
                <RESULT eventid="1281" points="635" reactiontime="+82" swimtime="00:02:11.38" resultid="3164" heatid="4065" lane="4" entrytime="00:02:10.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="100" swimtime="00:01:04.38" />
                    <SPLIT distance="150" swimtime="00:01:38.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="599" reactiontime="+83" swimtime="00:18:11.64" resultid="3165" heatid="4095" lane="5" entrytime="00:18:16.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:06.77" />
                    <SPLIT distance="150" swimtime="00:01:42.14" />
                    <SPLIT distance="200" swimtime="00:02:17.24" />
                    <SPLIT distance="250" swimtime="00:02:53.08" />
                    <SPLIT distance="300" swimtime="00:03:28.72" />
                    <SPLIT distance="350" swimtime="00:04:04.53" />
                    <SPLIT distance="400" swimtime="00:04:40.63" />
                    <SPLIT distance="450" swimtime="00:05:16.87" />
                    <SPLIT distance="500" swimtime="00:05:53.48" />
                    <SPLIT distance="550" swimtime="00:06:29.74" />
                    <SPLIT distance="600" swimtime="00:07:06.53" />
                    <SPLIT distance="650" swimtime="00:07:43.39" />
                    <SPLIT distance="700" swimtime="00:08:20.01" />
                    <SPLIT distance="750" swimtime="00:08:57.10" />
                    <SPLIT distance="800" swimtime="00:09:33.88" />
                    <SPLIT distance="850" swimtime="00:10:10.63" />
                    <SPLIT distance="900" swimtime="00:10:47.51" />
                    <SPLIT distance="950" swimtime="00:11:24.72" />
                    <SPLIT distance="1000" swimtime="00:12:01.80" />
                    <SPLIT distance="1050" swimtime="00:12:38.96" />
                    <SPLIT distance="1100" swimtime="00:13:16.27" />
                    <SPLIT distance="1150" swimtime="00:13:53.15" />
                    <SPLIT distance="1200" swimtime="00:14:30.21" />
                    <SPLIT distance="1250" swimtime="00:15:07.30" />
                    <SPLIT distance="1300" swimtime="00:15:44.77" />
                    <SPLIT distance="1350" swimtime="00:16:21.86" />
                    <SPLIT distance="1400" swimtime="00:16:59.48" />
                    <SPLIT distance="1450" swimtime="00:17:35.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="569" reactiontime="+78" swimtime="00:01:02.37" resultid="3166" heatid="4105" lane="5" entrytime="00:01:01.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="536" reactiontime="+81" swimtime="00:02:35.24" resultid="3167" heatid="4137" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:14.99" />
                    <SPLIT distance="150" swimtime="00:02:01.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="612" reactiontime="+80" swimtime="00:04:38.50" resultid="3168" heatid="4145" lane="5" entrytime="00:04:33.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:05.65" />
                    <SPLIT distance="150" swimtime="00:01:40.93" />
                    <SPLIT distance="200" swimtime="00:02:16.48" />
                    <SPLIT distance="250" swimtime="00:02:52.34" />
                    <SPLIT distance="300" swimtime="00:03:28.03" />
                    <SPLIT distance="350" swimtime="00:04:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="613" reactiontime="+80" swimtime="00:09:30.65" resultid="3169" heatid="4157" lane="5" entrytime="00:09:27.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:42.19" />
                    <SPLIT distance="200" swimtime="00:02:17.64" />
                    <SPLIT distance="250" swimtime="00:02:53.17" />
                    <SPLIT distance="300" swimtime="00:03:28.68" />
                    <SPLIT distance="350" swimtime="00:04:04.54" />
                    <SPLIT distance="400" swimtime="00:04:41.05" />
                    <SPLIT distance="450" swimtime="00:05:17.06" />
                    <SPLIT distance="500" swimtime="00:05:53.80" />
                    <SPLIT distance="550" swimtime="00:06:30.04" />
                    <SPLIT distance="600" swimtime="00:07:06.93" />
                    <SPLIT distance="650" swimtime="00:07:43.41" />
                    <SPLIT distance="700" swimtime="00:08:19.85" />
                    <SPLIT distance="750" swimtime="00:08:56.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Pacewicz" birthdate="2006-03-25" gender="M" nation="POL" license="101605700183" swrid="5170203" athleteid="3286">
              <RESULTS>
                <RESULT eventid="1258" points="551" reactiontime="+67" swimtime="00:00:29.27" resultid="3287" heatid="4060" lane="7" entrytime="00:00:29.25" entrycourse="LCM" />
                <RESULT eventid="1304" points="504" reactiontime="+69" swimtime="00:02:08.17" resultid="3288" heatid="4070" lane="3" entrytime="00:02:15.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="100" swimtime="00:01:02.32" />
                    <SPLIT distance="150" swimtime="00:01:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="542" reactiontime="+67" swimtime="00:00:27.30" resultid="3289" heatid="4093" lane="3" entrytime="00:00:27.46" entrycourse="LCM" />
                <RESULT eventid="1613" points="562" reactiontime="+65" swimtime="00:01:02.80" resultid="3290" heatid="4136" lane="3" entrytime="00:01:02.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="572" reactiontime="+62" swimtime="00:02:14.75" resultid="3291" heatid="4155" lane="6" entrytime="00:02:14.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:06.63" />
                    <SPLIT distance="150" swimtime="00:01:41.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Bednarek" birthdate="2009-04-26" gender="M" nation="POL" license="101605700242" swrid="5356127" athleteid="3212">
              <RESULTS>
                <RESULT eventid="1120" points="341" reactiontime="+78" swimtime="00:00:29.91" resultid="3213" heatid="4029" lane="9" entrytime="00:00:30.87" entrycourse="LCM" />
                <RESULT eventid="1258" points="319" reactiontime="+68" swimtime="00:00:35.09" resultid="3214" heatid="4059" lane="9" entrytime="00:00:36.05" entrycourse="LCM" />
                <RESULT eventid="1304" points="317" reactiontime="+60" swimtime="00:02:29.49" resultid="3215" heatid="4069" lane="5" entrytime="00:02:30.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                    <SPLIT distance="150" swimtime="00:01:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="352" reactiontime="+80" swimtime="00:01:06.39" resultid="3216" heatid="4112" lane="1" entrytime="00:01:06.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="313" reactiontime="+79" swimtime="00:01:16.32" resultid="3217" heatid="4135" lane="1" entrytime="00:01:15.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="314" reactiontime="+69" swimtime="00:02:44.50" resultid="3218" heatid="4154" lane="8" entrytime="00:02:50.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                    <SPLIT distance="150" swimtime="00:02:04.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Kacprzak" birthdate="2007-02-23" gender="M" nation="POL" license="101605700217" swrid="5198003" athleteid="3219">
              <RESULTS>
                <RESULT eventid="1120" points="439" reactiontime="+67" swimtime="00:00:27.50" resultid="3220" heatid="4030" lane="5" entrytime="00:00:27.25" entrycourse="LCM" />
                <RESULT eventid="1212" points="383" reactiontime="+68" swimtime="00:01:08.12" resultid="3221" heatid="4049" lane="6" entrytime="00:01:05.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="473" reactiontime="+68" swimtime="00:02:10.82" resultid="3222" heatid="4071" lane="3" entrytime="00:02:10.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="380" reactiontime="+60" swimtime="00:00:30.74" resultid="3223" heatid="4092" lane="5" entrytime="00:00:30.32" entrycourse="LCM" />
                <RESULT eventid="1475" points="468" reactiontime="+68" swimtime="00:01:00.38" resultid="3224" heatid="4113" lane="4" entrytime="00:00:58.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="483" reactiontime="+67" swimtime="00:04:40.36" resultid="3225" heatid="4147" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:08.78" />
                    <SPLIT distance="150" swimtime="00:01:44.92" />
                    <SPLIT distance="200" swimtime="00:02:21.22" />
                    <SPLIT distance="250" swimtime="00:02:57.16" />
                    <SPLIT distance="300" swimtime="00:03:33.10" />
                    <SPLIT distance="350" swimtime="00:04:08.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Stępka" birthdate="2008-02-25" gender="F" nation="POL" license="101605600233" swrid="5293172" athleteid="3233">
              <RESULTS>
                <RESULT eventid="1143" points="430" reactiontime="+74" swimtime="00:00:38.93" resultid="3234" heatid="4036" lane="5" entrytime="00:00:38.91" entrycourse="LCM" />
                <RESULT eventid="1327" points="379" reactiontime="+90" swimtime="00:01:28.57" resultid="3235" heatid="4075" lane="2" entrytime="00:01:27.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="302" reactiontime="+95" swimtime="00:00:36.38" resultid="3236" heatid="4084" lane="4" entrytime="00:00:42.63" entrycourse="LCM" />
                <RESULT eventid="1590" points="357" reactiontime="+74" swimtime="00:01:21.08" resultid="3237" heatid="4128" lane="5" entrytime="00:01:23.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="333" reactiontime="+84" swimtime="00:02:57.87" resultid="3238" heatid="4151" lane="0" entrytime="00:02:58.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:28.14" />
                    <SPLIT distance="150" swimtime="00:02:14.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Piekarska" birthdate="2006-09-26" gender="F" nation="POL" license="101605600298" swrid="5159131" athleteid="3111">
              <RESULTS>
                <RESULT eventid="1060" points="637" reactiontime="+76" swimtime="00:05:09.43" resultid="3112" heatid="4011" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:11.87" />
                    <SPLIT distance="150" swimtime="00:01:51.97" />
                    <SPLIT distance="200" swimtime="00:02:31.81" />
                    <SPLIT distance="250" swimtime="00:03:16.27" />
                    <SPLIT distance="300" swimtime="00:04:00.97" />
                    <SPLIT distance="350" swimtime="00:04:35.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="567" reactiontime="+71" swimtime="00:01:07.03" resultid="3113" heatid="4046" lane="4" entrytime="00:01:05.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="531" reactiontime="+72" swimtime="00:00:30.16" resultid="3114" heatid="4088" lane="4" entrytime="00:00:29.72" entrycourse="LCM" />
                <RESULT eventid="1544" points="602" reactiontime="+74" swimtime="00:02:24.20" resultid="3115" heatid="4123" lane="4" entrytime="00:02:23.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                    <SPLIT distance="100" swimtime="00:01:10.49" />
                    <SPLIT distance="150" swimtime="00:01:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="611" reactiontime="+71" swimtime="00:02:28.62" resultid="3116" heatid="4138" lane="5" entrytime="00:02:28.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:55.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="596" reactiontime="+76" swimtime="00:04:40.87" resultid="3117" heatid="4145" lane="8" entrytime="00:04:55.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:09.40" />
                    <SPLIT distance="150" swimtime="00:01:45.14" />
                    <SPLIT distance="200" swimtime="00:02:21.30" />
                    <SPLIT distance="250" swimtime="00:02:56.99" />
                    <SPLIT distance="300" swimtime="00:03:32.66" />
                    <SPLIT distance="350" swimtime="00:04:07.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Łuczak" birthdate="2008-01-29" gender="M" nation="POL" license="101605700237" swrid="4976843" athleteid="3182">
              <RESULTS>
                <RESULT eventid="1120" points="234" reactiontime="+84" swimtime="00:00:33.89" resultid="3183" heatid="4026" lane="3" entrytime="00:00:36.65" entrycourse="LCM" />
                <RESULT eventid="1258" points="219" swimtime="00:00:39.79" resultid="3184" heatid="4056" lane="3" />
                <RESULT eventid="1304" points="217" reactiontime="+86" swimtime="00:02:49.49" resultid="3185" heatid="4068" lane="5" entrytime="00:03:08.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:21.32" />
                    <SPLIT distance="150" swimtime="00:02:05.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="235" reactiontime="+84" swimtime="00:01:15.93" resultid="3186" heatid="4109" lane="3" entrytime="00:01:24.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="214" swimtime="00:01:26.67" resultid="3187" heatid="4131" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Franciszek" lastname="Jarczewski" birthdate="2005-12-10" gender="M" nation="POL" license="101605700239" swrid="5075910" athleteid="3125">
              <RESULTS>
                <RESULT eventid="1065" points="596" reactiontime="+73" swimtime="00:04:49.61" resultid="3126" heatid="4013" lane="3" entrytime="00:04:54.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="100" swimtime="00:01:04.63" />
                    <SPLIT distance="150" swimtime="00:01:42.39" />
                    <SPLIT distance="200" swimtime="00:02:19.39" />
                    <SPLIT distance="250" swimtime="00:03:00.96" />
                    <SPLIT distance="300" swimtime="00:03:42.86" />
                    <SPLIT distance="350" swimtime="00:04:16.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="499" reactiontime="+68" swimtime="00:01:02.38" resultid="3127" heatid="4049" lane="4" entrytime="00:01:01.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="549" reactiontime="+73" swimtime="00:09:11.97" resultid="3128" heatid="4096" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:06.49" />
                    <SPLIT distance="150" swimtime="00:01:41.28" />
                    <SPLIT distance="200" swimtime="00:02:16.27" />
                    <SPLIT distance="250" swimtime="00:02:50.90" />
                    <SPLIT distance="300" swimtime="00:03:25.48" />
                    <SPLIT distance="350" swimtime="00:04:00.22" />
                    <SPLIT distance="400" swimtime="00:04:34.93" />
                    <SPLIT distance="450" swimtime="00:05:09.64" />
                    <SPLIT distance="500" swimtime="00:05:44.28" />
                    <SPLIT distance="550" swimtime="00:06:18.85" />
                    <SPLIT distance="600" swimtime="00:06:53.61" />
                    <SPLIT distance="650" swimtime="00:07:28.63" />
                    <SPLIT distance="700" swimtime="00:08:04.15" />
                    <SPLIT distance="750" swimtime="00:08:38.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="534" reactiontime="+74" swimtime="00:02:16.47" resultid="3129" heatid="4125" lane="1" entrytime="00:02:16.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="100" swimtime="00:01:05.90" />
                    <SPLIT distance="150" swimtime="00:01:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="543" reactiontime="+71" swimtime="00:02:19.68" resultid="3130" heatid="4142" lane="6" entrytime="00:02:19.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:06.09" />
                    <SPLIT distance="150" swimtime="00:01:48.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="560" reactiontime="+72" swimtime="00:04:26.94" resultid="3131" heatid="4149" lane="1" entrytime="00:04:25.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                    <SPLIT distance="100" swimtime="00:01:03.60" />
                    <SPLIT distance="150" swimtime="00:01:37.31" />
                    <SPLIT distance="200" swimtime="00:02:11.59" />
                    <SPLIT distance="250" swimtime="00:02:45.51" />
                    <SPLIT distance="300" swimtime="00:03:19.86" />
                    <SPLIT distance="350" swimtime="00:03:53.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Wrzesińska" birthdate="2004-05-07" gender="F" nation="POL" license="101605600144" swrid="5034809" athleteid="3105">
              <RESULTS>
                <RESULT eventid="1060" points="635" reactiontime="+84" swimtime="00:05:09.78" resultid="3106" heatid="4011" lane="3" entrytime="00:05:14.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:01:52.19" />
                    <SPLIT distance="200" swimtime="00:02:33.04" />
                    <SPLIT distance="250" swimtime="00:03:16.69" />
                    <SPLIT distance="300" swimtime="00:03:59.69" />
                    <SPLIT distance="350" swimtime="00:04:35.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="640" reactiontime="+84" swimtime="00:17:47.85" resultid="3107" heatid="4095" lane="4" entrytime="00:17:40.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:06.60" />
                    <SPLIT distance="150" swimtime="00:01:41.85" />
                    <SPLIT distance="200" swimtime="00:02:16.79" />
                    <SPLIT distance="250" swimtime="00:02:52.28" />
                    <SPLIT distance="300" swimtime="00:03:27.96" />
                    <SPLIT distance="350" swimtime="00:04:03.31" />
                    <SPLIT distance="400" swimtime="00:04:38.78" />
                    <SPLIT distance="450" swimtime="00:05:14.31" />
                    <SPLIT distance="500" swimtime="00:05:50.10" />
                    <SPLIT distance="550" swimtime="00:06:25.72" />
                    <SPLIT distance="600" swimtime="00:07:01.31" />
                    <SPLIT distance="650" swimtime="00:07:36.97" />
                    <SPLIT distance="700" swimtime="00:08:12.86" />
                    <SPLIT distance="750" swimtime="00:08:48.63" />
                    <SPLIT distance="800" swimtime="00:09:24.26" />
                    <SPLIT distance="850" swimtime="00:10:00.08" />
                    <SPLIT distance="900" swimtime="00:10:36.45" />
                    <SPLIT distance="950" swimtime="00:11:12.42" />
                    <SPLIT distance="1000" swimtime="00:11:48.88" />
                    <SPLIT distance="1050" swimtime="00:12:25.06" />
                    <SPLIT distance="1100" swimtime="00:13:01.26" />
                    <SPLIT distance="1150" swimtime="00:13:37.59" />
                    <SPLIT distance="1200" swimtime="00:14:14.02" />
                    <SPLIT distance="1250" swimtime="00:14:49.85" />
                    <SPLIT distance="1300" swimtime="00:15:25.86" />
                    <SPLIT distance="1350" swimtime="00:16:01.79" />
                    <SPLIT distance="1400" swimtime="00:16:37.60" />
                    <SPLIT distance="1450" swimtime="00:17:12.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="555" reactiontime="+80" swimtime="00:02:49.25" resultid="3108" heatid="4116" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:02:05.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="650" reactiontime="+79" swimtime="00:04:32.88" resultid="3109" heatid="4145" lane="4" entrytime="00:04:30.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:05.53" />
                    <SPLIT distance="150" swimtime="00:01:40.49" />
                    <SPLIT distance="200" swimtime="00:02:15.37" />
                    <SPLIT distance="250" swimtime="00:02:49.81" />
                    <SPLIT distance="300" swimtime="00:03:24.42" />
                    <SPLIT distance="350" swimtime="00:03:58.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="653" reactiontime="+83" swimtime="00:09:18.60" resultid="3110" heatid="4157" lane="4" entrytime="00:09:19.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="150" swimtime="00:01:42.02" />
                    <SPLIT distance="200" swimtime="00:02:17.23" />
                    <SPLIT distance="250" swimtime="00:02:52.61" />
                    <SPLIT distance="300" swimtime="00:03:27.94" />
                    <SPLIT distance="350" swimtime="00:04:03.47" />
                    <SPLIT distance="400" swimtime="00:04:38.63" />
                    <SPLIT distance="450" swimtime="00:05:14.14" />
                    <SPLIT distance="500" swimtime="00:05:49.36" />
                    <SPLIT distance="550" swimtime="00:06:24.69" />
                    <SPLIT distance="600" swimtime="00:06:59.56" />
                    <SPLIT distance="650" swimtime="00:07:34.51" />
                    <SPLIT distance="700" swimtime="00:08:09.55" />
                    <SPLIT distance="750" swimtime="00:08:44.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Gomułka" birthdate="2004-07-02" gender="F" nation="POL" license="101605600143" swrid="5034811" athleteid="3239">
              <RESULTS>
                <RESULT eventid="1143" points="405" reactiontime="+69" swimtime="00:00:39.72" resultid="3240" heatid="4036" lane="7" entrytime="00:00:39.22" entrycourse="LCM" />
                <RESULT eventid="1327" points="422" reactiontime="+71" swimtime="00:01:25.46" resultid="3241" heatid="4076" lane="9" entrytime="00:01:22.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="487" reactiontime="+73" swimtime="00:02:56.74" resultid="3242" heatid="4118" lane="1" entrytime="00:02:56.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                    <SPLIT distance="100" swimtime="00:01:25.46" />
                    <SPLIT distance="150" swimtime="00:02:10.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="463" reactiontime="+78" swimtime="00:05:05.50" resultid="3243" heatid="4145" lane="0" entrytime="00:04:55.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:14.37" />
                    <SPLIT distance="150" swimtime="00:01:53.06" />
                    <SPLIT distance="200" swimtime="00:02:31.81" />
                    <SPLIT distance="250" swimtime="00:03:10.63" />
                    <SPLIT distance="300" swimtime="00:03:49.30" />
                    <SPLIT distance="350" swimtime="00:04:28.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Mańka" birthdate="2000-11-10" gender="M" nation="POL" license="101605700134" swrid="4630233" athleteid="3296">
              <RESULTS>
                <RESULT eventid="1613" points="609" reactiontime="+55" swimtime="00:01:01.15" resultid="3297" heatid="4132" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="616" reactiontime="+60" swimtime="00:02:11.48" resultid="3298" heatid="4155" lane="2" entrytime="00:02:15.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:06.57" />
                    <SPLIT distance="150" swimtime="00:01:39.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Woźniak" birthdate="2000-11-30" gender="M" nation="POL" license="101605700167" swrid="4630238" athleteid="3194">
              <RESULTS>
                <RESULT eventid="1120" points="626" reactiontime="+72" swimtime="00:00:24.44" resultid="3195" heatid="4032" lane="3" entrytime="00:00:24.31" entrycourse="LCM" />
                <RESULT eventid="1396" points="612" reactiontime="+72" swimtime="00:00:26.23" resultid="3196" heatid="4094" lane="3" entrytime="00:00:26.14" entrycourse="LCM" />
                <RESULT eventid="1446" status="DNS" swimtime="00:00:00.00" resultid="3197" heatid="4096" lane="2" />
                <RESULT eventid="1475" points="692" reactiontime="+71" swimtime="00:00:53.01" resultid="3198" heatid="4115" lane="5" entrytime="00:00:52.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="614" reactiontime="+74" swimtime="00:02:14.08" resultid="3199" heatid="4142" lane="4" entrytime="00:02:10.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                    <SPLIT distance="100" swimtime="00:01:02.85" />
                    <SPLIT distance="150" swimtime="00:01:42.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jagoda" lastname="Pawlak" birthdate="2009-01-03" gender="F" nation="POL" license="101605600244" swrid="5356913" athleteid="3157">
              <RESULTS>
                <RESULT eventid="1070" points="250" reactiontime="+83" swimtime="00:00:37.56" resultid="3158" heatid="4017" lane="7" entrytime="00:00:35.97" entrycourse="LCM" />
                <RESULT eventid="1143" points="238" reactiontime="+75" swimtime="00:00:47.39" resultid="3159" heatid="4034" lane="3" entrytime="00:00:47.39" entrycourse="LCM" />
                <RESULT eventid="1451" points="256" reactiontime="+86" swimtime="00:01:21.37" resultid="3160" heatid="4100" lane="4" entrytime="00:01:19.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="234" reactiontime="+95" swimtime="00:03:45.62" resultid="3161" heatid="4116" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.25" />
                    <SPLIT distance="100" swimtime="00:01:48.32" />
                    <SPLIT distance="150" swimtime="00:02:48.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Leśniak" birthdate="2004-09-28" gender="M" nation="POL" license="101605700176" swrid="5034907" athleteid="3206">
              <RESULTS>
                <RESULT eventid="1120" points="597" reactiontime="+66" swimtime="00:00:24.83" resultid="3207" heatid="4032" lane="2" entrytime="00:00:24.86" entrycourse="LCM" />
                <RESULT eventid="1304" points="620" reactiontime="+64" swimtime="00:01:59.61" resultid="3208" heatid="4072" lane="3" entrytime="00:01:58.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="100" swimtime="00:00:58.00" />
                    <SPLIT distance="150" swimtime="00:01:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="601" reactiontime="+65" swimtime="00:08:55.57" resultid="3209" heatid="4097" lane="3" entrytime="00:08:58.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                    <SPLIT distance="100" swimtime="00:01:03.93" />
                    <SPLIT distance="150" swimtime="00:01:37.97" />
                    <SPLIT distance="200" swimtime="00:02:11.88" />
                    <SPLIT distance="250" swimtime="00:02:45.44" />
                    <SPLIT distance="300" swimtime="00:03:19.25" />
                    <SPLIT distance="350" swimtime="00:03:52.42" />
                    <SPLIT distance="400" swimtime="00:04:26.15" />
                    <SPLIT distance="450" swimtime="00:05:00.32" />
                    <SPLIT distance="500" swimtime="00:05:34.06" />
                    <SPLIT distance="550" swimtime="00:06:07.75" />
                    <SPLIT distance="600" swimtime="00:06:41.59" />
                    <SPLIT distance="650" swimtime="00:07:15.45" />
                    <SPLIT distance="700" swimtime="00:07:49.47" />
                    <SPLIT distance="750" swimtime="00:08:22.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="646" reactiontime="+67" swimtime="00:00:54.25" resultid="3210" heatid="4115" lane="2" entrytime="00:00:53.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="627" reactiontime="+67" swimtime="00:04:17.02" resultid="3211" heatid="4149" lane="3" entrytime="00:04:13.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                    <SPLIT distance="100" swimtime="00:01:00.69" />
                    <SPLIT distance="150" swimtime="00:01:32.90" />
                    <SPLIT distance="200" swimtime="00:02:05.89" />
                    <SPLIT distance="250" swimtime="00:02:38.65" />
                    <SPLIT distance="300" swimtime="00:03:11.65" />
                    <SPLIT distance="350" swimtime="00:03:45.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Jarczewski" birthdate="2007-07-12" gender="M" nation="POL" license="101605700241" swrid="4901064" athleteid="3226">
              <RESULTS>
                <RESULT eventid="1120" points="296" reactiontime="+70" swimtime="00:00:31.37" resultid="3227" heatid="4028" lane="4" entrytime="00:00:31.10" entrycourse="LCM" />
                <RESULT eventid="1258" points="296" reactiontime="+64" swimtime="00:00:36.00" resultid="3228" heatid="4058" lane="4" entrytime="00:00:36.75" entrycourse="LCM" />
                <RESULT eventid="1304" points="359" reactiontime="+75" swimtime="00:02:23.41" resultid="3229" heatid="4070" lane="0" entrytime="00:02:26.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:09.62" />
                    <SPLIT distance="150" swimtime="00:01:47.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="329" reactiontime="+69" swimtime="00:01:07.90" resultid="3230" heatid="4111" lane="6" entrytime="00:01:08.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="314" reactiontime="+68" swimtime="00:02:47.64" resultid="3231" heatid="4141" lane="6" entrytime="00:02:46.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                    <SPLIT distance="100" swimtime="00:01:17.76" />
                    <SPLIT distance="150" swimtime="00:02:09.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="334" reactiontime="+60" swimtime="00:02:41.18" resultid="3232" heatid="4154" lane="6" entrytime="00:02:41.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                    <SPLIT distance="100" swimtime="00:01:19.57" />
                    <SPLIT distance="150" swimtime="00:02:01.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Kieruzel" birthdate="2005-12-11" gender="F" nation="POL" license="101605600263" swrid="5190452" athleteid="3170">
              <RESULTS>
                <RESULT eventid="1070" points="469" reactiontime="+72" swimtime="00:00:30.45" resultid="3171" heatid="4021" lane="9" entrytime="00:00:29.84" entrycourse="LCM" />
                <RESULT eventid="1281" points="524" reactiontime="+73" swimtime="00:02:20.09" resultid="3172" heatid="4064" lane="6" entrytime="00:02:21.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:07.97" />
                    <SPLIT distance="150" swimtime="00:01:44.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="464" reactiontime="+72" swimtime="00:19:48.13" resultid="3173" heatid="4095" lane="6" entrytime="00:19:37.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:15.14" />
                    <SPLIT distance="150" swimtime="00:01:55.56" />
                    <SPLIT distance="200" swimtime="00:02:35.81" />
                    <SPLIT distance="250" swimtime="00:03:15.22" />
                    <SPLIT distance="300" swimtime="00:03:55.08" />
                    <SPLIT distance="350" swimtime="00:04:35.06" />
                    <SPLIT distance="400" swimtime="00:05:14.68" />
                    <SPLIT distance="450" swimtime="00:05:54.50" />
                    <SPLIT distance="500" swimtime="00:06:34.42" />
                    <SPLIT distance="550" swimtime="00:07:14.42" />
                    <SPLIT distance="600" swimtime="00:07:54.41" />
                    <SPLIT distance="650" swimtime="00:08:34.19" />
                    <SPLIT distance="700" swimtime="00:09:14.26" />
                    <SPLIT distance="750" swimtime="00:09:53.88" />
                    <SPLIT distance="800" swimtime="00:10:33.90" />
                    <SPLIT distance="850" swimtime="00:11:14.01" />
                    <SPLIT distance="900" swimtime="00:11:53.96" />
                    <SPLIT distance="950" swimtime="00:12:33.93" />
                    <SPLIT distance="1000" swimtime="00:13:13.82" />
                    <SPLIT distance="1050" swimtime="00:13:53.20" />
                    <SPLIT distance="1100" swimtime="00:14:31.94" />
                    <SPLIT distance="1150" swimtime="00:15:11.78" />
                    <SPLIT distance="1200" swimtime="00:15:52.17" />
                    <SPLIT distance="1250" swimtime="00:16:32.78" />
                    <SPLIT distance="1300" swimtime="00:17:12.48" />
                    <SPLIT distance="1350" swimtime="00:17:51.77" />
                    <SPLIT distance="1400" swimtime="00:18:30.93" />
                    <SPLIT distance="1450" swimtime="00:19:10.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="470" reactiontime="+75" swimtime="00:01:06.50" resultid="3174" heatid="4103" lane="6" entrytime="00:01:05.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="517" reactiontime="+74" swimtime="00:04:54.53" resultid="3175" heatid="4145" lane="1" entrytime="00:04:53.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:10.27" />
                    <SPLIT distance="150" swimtime="00:01:47.43" />
                    <SPLIT distance="200" swimtime="00:02:25.21" />
                    <SPLIT distance="250" swimtime="00:03:02.74" />
                    <SPLIT distance="300" swimtime="00:03:40.77" />
                    <SPLIT distance="350" swimtime="00:04:18.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="489" reactiontime="+77" swimtime="00:10:15.26" resultid="3176" heatid="4157" lane="2" entrytime="00:10:10.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:14.48" />
                    <SPLIT distance="150" swimtime="00:01:54.25" />
                    <SPLIT distance="200" swimtime="00:02:33.50" />
                    <SPLIT distance="250" swimtime="00:03:11.64" />
                    <SPLIT distance="300" swimtime="00:03:49.85" />
                    <SPLIT distance="350" swimtime="00:04:27.90" />
                    <SPLIT distance="400" swimtime="00:05:06.49" />
                    <SPLIT distance="450" swimtime="00:05:45.58" />
                    <SPLIT distance="500" swimtime="00:06:24.44" />
                    <SPLIT distance="550" swimtime="00:07:03.71" />
                    <SPLIT distance="600" swimtime="00:07:42.63" />
                    <SPLIT distance="650" swimtime="00:08:21.85" />
                    <SPLIT distance="700" swimtime="00:09:01.01" />
                    <SPLIT distance="750" swimtime="00:09:38.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02805" nation="POL" region="05" clubid="2757" name="MUKS Zgierz">
          <ATHLETES>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-26" gender="F" nation="POL" license="502805600123" athleteid="2758">
              <RESULTS>
                <RESULT eventid="1070" points="53" swimtime="00:01:02.85" resultid="2759" heatid="4014" lane="4" />
                <RESULT eventid="1327" points="96" swimtime="00:02:19.99" resultid="2760" heatid="4073" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="72" swimtime="00:02:03.90" resultid="2761" heatid="4099" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Bednarek" birthdate="1951-03-24" gender="M" nation="POL" license="502805700052" athleteid="2792">
              <RESULTS>
                <RESULT eventid="1120" points="182" swimtime="00:00:36.84" resultid="2793" heatid="4026" lane="0" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="2794" heatid="4068" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" swrid="4992745" athleteid="2802">
              <RESULTS>
                <RESULT eventid="1189" points="457" reactiontime="+88" swimtime="00:01:12.01" resultid="2803" heatid="4044" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="442" reactiontime="+82" swimtime="00:00:32.06" resultid="2804" heatid="4084" lane="7" />
                <RESULT eventid="1544" points="330" reactiontime="+88" swimtime="00:02:56.12" resultid="2805" heatid="4123" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:21.42" />
                    <SPLIT distance="150" swimtime="00:02:07.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Błasiak" birthdate="1955-03-16" gender="M" nation="POL" license="502805700037" athleteid="2819">
              <RESULTS>
                <RESULT eventid="1304" points="90" reactiontime="+98" swimtime="00:03:47.10" resultid="2820" heatid="4066" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                    <SPLIT distance="100" swimtime="00:03:47.16" />
                    <SPLIT distance="150" swimtime="00:02:53.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="58" reactiontime="+96" swimtime="00:05:24.98" resultid="2821" heatid="4119" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.00" />
                    <SPLIT distance="100" swimtime="00:02:39.47" />
                    <SPLIT distance="150" swimtime="00:04:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="61" reactiontime="+97" swimtime="00:04:48.67" resultid="2822" heatid="4140" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.13" />
                    <SPLIT distance="100" swimtime="00:02:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="55" swimtime="00:04:54.06" resultid="2823" heatid="4153" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.02" />
                    <SPLIT distance="100" swimtime="00:02:27.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" swrid="4754660" athleteid="2762">
              <RESULTS>
                <RESULT eventid="1070" points="328" reactiontime="+88" swimtime="00:00:34.31" resultid="2763" heatid="4016" lane="8" />
                <RESULT eventid="1373" points="304" reactiontime="+96" swimtime="00:00:36.30" resultid="2764" heatid="4084" lane="9" />
                <RESULT eventid="1451" points="278" reactiontime="+92" swimtime="00:01:19.22" resultid="2765" heatid="4100" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="223" reactiontime="+88" swimtime="00:01:34.90" resultid="2766" heatid="4126" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Łatecki" birthdate="1957-05-25" gender="M" nation="POL" license="502805700022" athleteid="2816">
              <RESULTS>
                <RESULT eventid="1304" points="58" swimtime="00:04:22.65" resultid="2817" heatid="4067" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.39" />
                    <SPLIT distance="100" swimtime="00:02:03.68" />
                    <SPLIT distance="150" swimtime="00:03:14.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" status="DNS" swimtime="00:00:00.00" resultid="2818" heatid="4153" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Klusek" birthdate="1975-01-12" gender="F" nation="POL" license="502805600030" athleteid="2806">
              <RESULTS>
                <RESULT eventid="1189" points="245" swimtime="00:01:28.62" resultid="2807" heatid="4044" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="272" reactiontime="+99" swimtime="00:00:37.66" resultid="2808" heatid="4083" lane="7" />
                <RESULT eventid="1544" points="239" swimtime="00:03:16.22" resultid="2809" heatid="4123" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:29.75" />
                    <SPLIT distance="150" swimtime="00:02:21.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="294" swimtime="00:03:09.66" resultid="2810" heatid="4137" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="100" swimtime="00:01:31.49" />
                    <SPLIT distance="150" swimtime="00:02:25.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-01-05" gender="F" nation="POL" license="502805600055" swrid="4655158" athleteid="2795">
              <RESULTS>
                <RESULT eventid="1143" points="232" reactiontime="+65" swimtime="00:00:47.83" resultid="2796" heatid="4034" lane="0" />
                <RESULT eventid="1327" points="220" reactiontime="+87" swimtime="00:01:46.17" resultid="2797" heatid="4073" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="228" reactiontime="+73" swimtime="00:03:47.50" resultid="2798" heatid="4116" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.27" />
                    <SPLIT distance="100" swimtime="00:01:50.31" />
                    <SPLIT distance="150" swimtime="00:02:50.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Chwiałkowski" birthdate="1985-11-09" gender="M" nation="POL" license="502805700033" athleteid="2824">
              <RESULTS>
                <RESULT eventid="1304" points="240" swimtime="00:02:44.00" resultid="2825" heatid="4067" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="150" swimtime="00:01:59.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="234" reactiontime="+99" swimtime="00:05:57.11" resultid="2826" heatid="4147" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="100" swimtime="00:01:20.09" />
                    <SPLIT distance="150" swimtime="00:02:04.34" />
                    <SPLIT distance="200" swimtime="00:02:50.87" />
                    <SPLIT distance="250" swimtime="00:03:37.86" />
                    <SPLIT distance="300" swimtime="00:04:25.81" />
                    <SPLIT distance="350" swimtime="00:05:12.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Przytulski" birthdate="1957-01-09" gender="M" nation="POL" license="502805700049" swrid="4754657" athleteid="2811">
              <RESULTS>
                <RESULT eventid="1258" points="246" reactiontime="+87" swimtime="00:00:38.30" resultid="2812" heatid="4057" lane="8" />
                <RESULT eventid="1304" points="232" reactiontime="+91" swimtime="00:02:45.82" resultid="2813" heatid="4067" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:02:00.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="287" reactiontime="+94" swimtime="00:01:11.08" resultid="2814" heatid="4106" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="209" reactiontime="+83" swimtime="00:01:27.24" resultid="2815" heatid="4133" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Wiczel" birthdate="1948-01-22" gender="M" nation="POL" license="502805700021" swrid="4876444" athleteid="2799">
              <RESULTS>
                <RESULT eventid="1166" points="222" swimtime="00:00:42.83" resultid="2800" heatid="4039" lane="1" />
                <RESULT eventid="1350" points="180" reactiontime="+96" swimtime="00:01:40.59" resultid="2801" heatid="4077" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Gajda" birthdate="1978-02-23" gender="M" nation="POL" license="502805700059" swrid="5272788" athleteid="2787">
              <RESULTS>
                <RESULT eventid="1120" points="308" reactiontime="+84" swimtime="00:00:30.94" resultid="2788" heatid="4023" lane="5" />
                <RESULT eventid="1258" points="279" reactiontime="+73" swimtime="00:00:36.72" resultid="2789" heatid="4056" lane="7" />
                <RESULT eventid="1475" points="275" reactiontime="+87" swimtime="00:01:12.13" resultid="2790" heatid="4107" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="234" reactiontime="+74" swimtime="00:01:24.08" resultid="2791" heatid="4133" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Wojciechowski" birthdate="1949-02-07" gender="M" nation="POL" license="502805700047" swrid="5240290" athleteid="2779">
              <RESULTS>
                <RESULT eventid="1120" points="163" swimtime="00:00:38.26" resultid="2780" heatid="4025" lane="6" />
                <RESULT eventid="1166" points="219" swimtime="00:00:43.02" resultid="2781" heatid="4038" lane="6" />
                <RESULT eventid="1350" points="164" swimtime="00:01:43.72" resultid="2782" heatid="4078" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Maciejczyk" birthdate="1947-12-03" gender="M" nation="POL" license="502805700048" swrid="4302705" athleteid="2776">
              <RESULTS>
                <RESULT eventid="1120" points="191" reactiontime="+75" swimtime="00:00:36.29" resultid="2777" heatid="4026" lane="9" />
                <RESULT eventid="1396" status="DNS" swimtime="00:00:00.00" resultid="2778" heatid="4089" lane="5" />
                <RESULT eventid="1475" points="150" reactiontime="+96" swimtime="00:01:28.18" resultid="4226" heatid="4106" lane="8" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Węgrzycka" birthdate="1977-01-26" gender="F" nation="POL" license="502805600056" athleteid="2767">
              <RESULTS>
                <RESULT eventid="1070" points="164" swimtime="00:00:43.22" resultid="2768" heatid="4016" lane="7" />
                <RESULT eventid="1143" points="162" swimtime="00:00:53.91" resultid="2769" heatid="4034" lane="7" />
                <RESULT eventid="1451" points="141" swimtime="00:01:39.17" resultid="2770" heatid="4099" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Dziarek" birthdate="1959-02-19" gender="M" nation="POL" license="502805700029" swrid="4841500" athleteid="2771">
              <RESULTS>
                <RESULT eventid="1120" points="241" swimtime="00:00:33.56" resultid="2772" heatid="4025" lane="7" />
                <RESULT eventid="1304" points="215" swimtime="00:02:50.02" resultid="2773" heatid="4067" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="150" swimtime="00:02:03.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="230" swimtime="00:01:16.52" resultid="2774" heatid="4107" lane="0" />
                <RESULT eventid="1705" points="200" swimtime="00:06:15.96" resultid="2775" heatid="4147" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:26.69" />
                    <SPLIT distance="150" swimtime="00:02:13.95" />
                    <SPLIT distance="200" swimtime="00:03:01.91" />
                    <SPLIT distance="250" swimtime="00:03:50.88" />
                    <SPLIT distance="300" swimtime="00:06:15.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Maciejewski" birthdate="1974-04-11" gender="M" nation="POL" license="502805700028" swrid="5373991" athleteid="2783">
              <RESULTS>
                <RESULT eventid="1120" points="247" reactiontime="+92" swimtime="00:00:33.30" resultid="2784" heatid="4025" lane="8" />
                <RESULT eventid="1350" points="185" reactiontime="+96" swimtime="00:01:39.72" resultid="2785" heatid="4077" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="212" reactiontime="+93" swimtime="00:01:18.67" resultid="2786" heatid="4109" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10414" nation="POL" region="14" clubid="2109" name="Klub Sportowy Mako">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" license="510414700009" swrid="4655152" athleteid="2110">
              <RESULTS>
                <RESULT eventid="1166" points="185" reactiontime="+80" swimtime="00:00:45.48" resultid="2111" heatid="4038" lane="2" />
                <RESULT eventid="1350" points="153" reactiontime="+87" swimtime="00:01:46.31" resultid="2112" heatid="4077" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="127" reactiontime="+81" swimtime="00:01:33.17" resultid="2113" heatid="4108" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="129" reactiontime="+84" swimtime="00:07:15.30" resultid="2114" heatid="4146" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                    <SPLIT distance="100" swimtime="00:01:39.88" />
                    <SPLIT distance="150" swimtime="00:02:37.14" />
                    <SPLIT distance="200" swimtime="00:03:33.73" />
                    <SPLIT distance="250" swimtime="00:04:30.31" />
                    <SPLIT distance="300" swimtime="00:05:26.57" />
                    <SPLIT distance="350" swimtime="00:06:23.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00505" nation="POL" region="05" clubid="3054" name="TP Olimpijczyk Aleksandrów Łódzki">
          <ATHLETES>
            <ATHLETE firstname="Natalia" lastname="Mikuła" birthdate="2006-08-28" gender="F" nation="POL" license="100505600103" swrid="5113367" athleteid="3061">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1070" reactiontime="+48" status="DSQ" swimtime="00:00:30.40" resultid="3062" heatid="4020" lane="6" entrytime="00:00:29.96" entrycourse="LCM" />
                <RESULT eventid="1235" points="432" reactiontime="+74" swimtime="00:00:35.68" resultid="3063" heatid="4052" lane="1" />
                <RESULT eventid="1281" points="515" reactiontime="+77" swimtime="00:02:20.88" resultid="3064" heatid="4065" lane="0" entrytime="00:02:19.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="150" swimtime="00:01:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="444" reactiontime="+76" swimtime="00:01:07.74" resultid="3065" heatid="4103" lane="1" entrytime="00:01:05.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="528" reactiontime="+70" swimtime="00:09:59.76" resultid="3066" heatid="4157" lane="3" entrytime="00:09:58.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:44.58" />
                    <SPLIT distance="200" swimtime="00:02:21.38" />
                    <SPLIT distance="250" swimtime="00:02:58.52" />
                    <SPLIT distance="300" swimtime="00:03:35.84" />
                    <SPLIT distance="350" swimtime="00:04:13.73" />
                    <SPLIT distance="400" swimtime="00:04:51.72" />
                    <SPLIT distance="450" swimtime="00:05:30.10" />
                    <SPLIT distance="500" swimtime="00:06:08.53" />
                    <SPLIT distance="550" swimtime="00:06:47.30" />
                    <SPLIT distance="600" swimtime="00:07:26.36" />
                    <SPLIT distance="650" swimtime="00:08:05.45" />
                    <SPLIT distance="700" swimtime="00:08:44.16" />
                    <SPLIT distance="750" swimtime="00:09:22.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nadia" lastname="Walczak" birthdate="2006-05-30" gender="F" nation="POL" license="100505600200" swrid="5456469" athleteid="3095">
              <RESULTS>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="3096" heatid="4101" lane="5" entrytime="00:01:12.92" entrycourse="LCM" />
                <RESULT eventid="1682" status="DNS" swimtime="00:00:00.00" resultid="3097" heatid="4143" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Wisiałkowski" birthdate="2004-01-19" gender="M" nation="POL" license="100505700231" swrid="5034888" athleteid="3852">
              <RESULTS>
                <RESULT eventid="1166" status="DNS" swimtime="00:00:00.00" resultid="3853" heatid="4039" lane="0" />
                <RESULT eventid="1350" status="DNS" swimtime="00:00:00.00" resultid="3854" heatid="4077" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Oleski" birthdate="2003-12-28" gender="M" nation="POL" license="100505700195" swrid="5086155" athleteid="3089">
              <RESULTS>
                <RESULT eventid="1212" points="638" reactiontime="+69" swimtime="00:00:57.49" resultid="3090" heatid="4050" lane="3" entrytime="00:00:57.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" status="DNS" swimtime="00:00:00.00" resultid="3091" heatid="4094" lane="5" entrytime="00:00:25.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Pietrzyk" birthdate="2007-07-14" gender="F" nation="POL" license="100505600112" swrid="5164101" athleteid="3067">
              <RESULTS>
                <RESULT eventid="1143" points="586" reactiontime="+76" swimtime="00:00:35.12" resultid="3068" heatid="4037" lane="5" entrytime="00:00:34.73" entrycourse="LCM" />
                <RESULT eventid="1189" points="471" reactiontime="+82" swimtime="00:01:11.30" resultid="3069" heatid="4045" lane="3" entrytime="00:01:11.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1327" points="559" reactiontime="+77" swimtime="00:01:17.83" resultid="3070" heatid="4076" lane="5" entrytime="00:01:15.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="439" reactiontime="+76" swimtime="00:00:32.13" resultid="3071" heatid="4087" lane="5" entrytime="00:00:31.80" entrycourse="LCM" />
                <RESULT eventid="1498" points="575" reactiontime="+79" swimtime="00:02:47.20" resultid="3072" heatid="4118" lane="4" entrytime="00:02:44.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:01:20.55" />
                    <SPLIT distance="150" swimtime="00:02:04.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="536" reactiontime="+82" swimtime="00:02:35.24" resultid="3073" heatid="4138" lane="1" entrytime="00:02:34.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                    <SPLIT distance="150" swimtime="00:01:57.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sara" lastname="Motyl" birthdate="2003-09-16" gender="F" nation="POL" license="100505600193" swrid="4933042" athleteid="3074">
              <RESULTS>
                <RESULT eventid="1143" points="592" reactiontime="+67" swimtime="00:00:35.01" resultid="3075" heatid="4037" lane="3" entrytime="00:00:34.90" entrycourse="LCM" />
                <RESULT eventid="1327" points="570" reactiontime="+67" swimtime="00:01:17.31" resultid="3076" heatid="4076" lane="3" entrytime="00:01:16.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="482" reactiontime="+66" swimtime="00:00:31.14" resultid="3077" heatid="4088" lane="8" entrytime="00:00:30.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Dukowska" birthdate="2006-06-12" gender="F" nation="POL" license="100505600178" swrid="5183193" athleteid="3055">
              <RESULTS>
                <RESULT eventid="1070" points="492" reactiontime="+66" swimtime="00:00:29.97" resultid="3056" heatid="4020" lane="3" entrytime="00:00:29.93" entrycourse="LCM" />
                <RESULT eventid="1189" points="404" reactiontime="+64" swimtime="00:01:14.99" resultid="3057" heatid="4044" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="561" reactiontime="+77" swimtime="00:02:16.97" resultid="3058" heatid="4064" lane="3" entrytime="00:02:21.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:06.57" />
                    <SPLIT distance="150" swimtime="00:01:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="522" reactiontime="+65" swimtime="00:01:04.20" resultid="3059" heatid="4105" lane="9" entrytime="00:01:03.87" entrycourse="LCM" />
                <RESULT eventid="1636" points="499" reactiontime="+75" swimtime="00:02:38.95" resultid="3060" heatid="4137" lane="4" entrytime="00:02:38.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:15.28" />
                    <SPLIT distance="150" swimtime="00:02:02.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Łopaciński" birthdate="2005-04-19" gender="M" nation="POL" license="100505700232" swrid="5164097" athleteid="3078">
              <RESULTS>
                <RESULT eventid="1166" points="463" reactiontime="+73" swimtime="00:00:33.53" resultid="3079" heatid="4043" lane="9" entrytime="00:00:33.60" entrycourse="LCM" />
                <RESULT eventid="1350" points="453" reactiontime="+76" swimtime="00:01:14.01" resultid="3080" heatid="4081" lane="8" entrytime="00:01:13.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="451" reactiontime="+77" swimtime="00:01:01.14" resultid="3081" heatid="4113" lane="5" entrytime="00:00:59.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="481" reactiontime="+77" swimtime="00:02:40.86" resultid="3082" heatid="4122" lane="7" entrytime="00:02:39.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:18.64" />
                    <SPLIT distance="150" swimtime="00:02:00.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Trafalska" birthdate="2007-01-30" gender="F" nation="POL" license="100505600151" swrid="5220872" athleteid="3083">
              <RESULTS>
                <RESULT eventid="1189" points="352" reactiontime="+87" swimtime="00:01:18.53" resultid="3084" heatid="4044" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="509" reactiontime="+79" swimtime="00:02:21.41" resultid="3085" heatid="4064" lane="5" entrytime="00:02:20.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:09.68" />
                    <SPLIT distance="150" swimtime="00:01:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="383" reactiontime="+88" swimtime="00:00:33.62" resultid="3086" heatid="4083" lane="1" />
                <RESULT eventid="1451" points="479" reactiontime="+65" swimtime="00:01:06.08" resultid="3087" heatid="4103" lane="8" entrytime="00:01:06.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="500" reactiontime="+79" swimtime="00:10:10.62" resultid="3088" heatid="4157" lane="6" entrytime="00:09:59.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:09.34" />
                    <SPLIT distance="150" swimtime="00:01:46.59" />
                    <SPLIT distance="200" swimtime="00:02:24.63" />
                    <SPLIT distance="250" swimtime="00:03:02.60" />
                    <SPLIT distance="300" swimtime="00:03:41.29" />
                    <SPLIT distance="350" swimtime="00:04:20.16" />
                    <SPLIT distance="400" swimtime="00:04:59.61" />
                    <SPLIT distance="450" swimtime="00:05:38.35" />
                    <SPLIT distance="500" swimtime="00:06:17.68" />
                    <SPLIT distance="550" swimtime="00:06:56.36" />
                    <SPLIT distance="600" swimtime="00:07:35.63" />
                    <SPLIT distance="650" swimtime="00:08:14.41" />
                    <SPLIT distance="700" swimtime="00:08:54.15" />
                    <SPLIT distance="750" swimtime="00:09:33.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Ciesielski" birthdate="2004-04-04" gender="M" nation="POL" license="100505700190" swrid="5101081" athleteid="3098">
              <RESULTS>
                <RESULT eventid="1475" points="644" reactiontime="+72" swimtime="00:00:54.31" resultid="3099" heatid="4115" lane="3" entrytime="00:00:52.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Kilar" birthdate="2004-11-10" gender="M" nation="POL" license="100505700192" swrid="5034850" athleteid="3092">
              <RESULTS>
                <RESULT eventid="1304" points="535" reactiontime="+74" swimtime="00:02:05.63" resultid="3093" heatid="4072" lane="8" entrytime="00:02:04.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                    <SPLIT distance="100" swimtime="00:01:01.16" />
                    <SPLIT distance="150" swimtime="00:01:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="541" reactiontime="+57" swimtime="00:00:57.56" resultid="3094" heatid="4114" lane="2" entrytime="00:00:56.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00305" nation="POL" region="05" clubid="3312" name="UKS Nawa Skierniewice">
          <ATHLETES>
            <ATHLETE firstname="Kornelia" lastname="Walz" birthdate="2000-02-21" gender="F" nation="POL" license="100305600123" swrid="4648193" athleteid="3361">
              <RESULTS>
                <RESULT eventid="1070" points="578" reactiontime="+68" swimtime="00:00:28.40" resultid="3362" heatid="4015" lane="8" />
                <RESULT eventid="1235" points="515" reactiontime="+68" swimtime="00:00:33.65" resultid="3363" heatid="4051" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Maszewski" birthdate="2006-08-23" gender="M" nation="POL" license="100305700189" swrid="5075874" athleteid="3417">
              <RESULTS>
                <RESULT eventid="1120" points="461" reactiontime="+76" swimtime="00:00:27.06" resultid="3418" heatid="4030" lane="4" entrytime="00:00:26.97" entrycourse="LCM" />
                <RESULT eventid="1166" points="359" reactiontime="+74" swimtime="00:00:36.51" resultid="3419" heatid="4042" lane="9" entrytime="00:00:36.30" entrycourse="LCM" />
                <RESULT eventid="1304" points="385" reactiontime="+86" swimtime="00:02:20.13" resultid="3420" heatid="4070" lane="1" entrytime="00:02:19.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="150" swimtime="00:01:46.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="325" swimtime="00:01:22.65" resultid="3421" heatid="4079" lane="4" entrytime="00:01:22.91" entrycourse="LCM" />
                <RESULT eventid="1475" points="469" reactiontime="+81" swimtime="00:01:00.37" resultid="3422" heatid="4112" lane="5" entrytime="00:01:01.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Brodowski" birthdate="2007-04-10" gender="M" nation="POL" license="100305700209" swrid="5198024" athleteid="3446">
              <RESULTS>
                <RESULT eventid="1166" points="349" reactiontime="+80" swimtime="00:00:36.83" resultid="3447" heatid="4041" lane="3" entrytime="00:00:37.89" entrycourse="LCM" />
                <RESULT eventid="1304" points="283" reactiontime="+83" swimtime="00:02:35.27" resultid="3448" heatid="4069" lane="7" entrytime="00:02:37.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:57.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="325" reactiontime="+84" swimtime="00:01:22.70" resultid="3449" heatid="4080" lane="0" entrytime="00:01:21.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="339" reactiontime="+72" swimtime="00:01:07.27" resultid="3450" heatid="4112" lane="8" entrytime="00:01:06.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="353" reactiontime="+78" swimtime="00:02:58.39" resultid="3451" heatid="4121" lane="7" entrytime="00:03:00.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:27.76" />
                    <SPLIT distance="150" swimtime="00:02:13.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Inez" lastname="Sarna" birthdate="2007-03-05" gender="F" nation="POL" license="100305600208" swrid="5152517" athleteid="3349">
              <RESULTS>
                <RESULT eventid="1070" points="524" reactiontime="+78" swimtime="00:00:29.35" resultid="3350" heatid="4021" lane="3" entrytime="00:00:29.42" entrycourse="LCM" />
                <RESULT eventid="1235" points="495" reactiontime="+65" swimtime="00:00:34.10" resultid="3351" heatid="4055" lane="9" entrytime="00:00:33.30" entrycourse="LCM" />
                <RESULT eventid="1451" points="515" reactiontime="+81" swimtime="00:01:04.48" resultid="3352" heatid="4104" lane="9" entrytime="00:01:04.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="516" reactiontime="+65" swimtime="00:01:11.75" resultid="3353" heatid="4130" lane="1" entrytime="00:01:11.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="440" reactiontime="+64" swimtime="00:02:42.07" resultid="3354" heatid="4151" lane="3" entrytime="00:02:44.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:18.72" />
                    <SPLIT distance="150" swimtime="00:02:01.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nadia" lastname="Lipowska" birthdate="2006-11-01" gender="F" nation="POL" license="100305600187" swrid="5075872" athleteid="3337">
              <RESULTS>
                <RESULT eventid="1070" points="572" reactiontime="+83" swimtime="00:00:28.50" resultid="3338" heatid="4022" lane="0" entrytime="00:00:28.97" entrycourse="LCM" />
                <RESULT eventid="1281" points="617" reactiontime="+77" swimtime="00:02:12.70" resultid="3339" heatid="4065" lane="3" entrytime="00:02:14.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:04.35" />
                    <SPLIT distance="150" swimtime="00:01:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="574" reactiontime="+79" swimtime="00:01:02.19" resultid="3340" heatid="4105" lane="2" entrytime="00:01:02.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="548" reactiontime="+79" swimtime="00:04:48.87" resultid="3341" heatid="4145" lane="2" entrytime="00:04:48.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:08.58" />
                    <SPLIT distance="150" swimtime="00:01:45.62" />
                    <SPLIT distance="200" swimtime="00:02:22.79" />
                    <SPLIT distance="250" swimtime="00:03:00.17" />
                    <SPLIT distance="300" swimtime="00:03:37.43" />
                    <SPLIT distance="350" swimtime="00:04:14.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="492" reactiontime="+81" swimtime="00:10:13.94" resultid="3342" heatid="4157" lane="7" entrytime="00:10:23.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:52.70" />
                    <SPLIT distance="200" swimtime="00:02:32.05" />
                    <SPLIT distance="250" swimtime="00:03:11.64" />
                    <SPLIT distance="300" swimtime="00:03:51.54" />
                    <SPLIT distance="350" swimtime="00:04:30.55" />
                    <SPLIT distance="400" swimtime="00:05:09.97" />
                    <SPLIT distance="450" swimtime="00:05:48.87" />
                    <SPLIT distance="500" swimtime="00:06:28.27" />
                    <SPLIT distance="550" swimtime="00:07:07.20" />
                    <SPLIT distance="600" swimtime="00:07:46.40" />
                    <SPLIT distance="650" swimtime="00:08:25.11" />
                    <SPLIT distance="700" swimtime="00:09:03.66" />
                    <SPLIT distance="750" swimtime="00:09:39.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Lesiak" birthdate="2008-07-18" gender="F" nation="POL" license="100305600232" swrid="5244122" athleteid="3381">
              <RESULTS>
                <RESULT eventid="1070" points="493" reactiontime="+81" swimtime="00:00:29.95" resultid="3382" heatid="4019" lane="2" entrytime="00:00:31.68" entrycourse="LCM" />
                <RESULT eventid="1143" points="559" reactiontime="+71" swimtime="00:00:35.68" resultid="3383" heatid="4037" lane="7" entrytime="00:00:35.80" entrycourse="LCM" />
                <RESULT eventid="1281" points="445" reactiontime="+76" swimtime="00:02:27.93" resultid="3384" heatid="4062" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                    <SPLIT distance="150" swimtime="00:01:51.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1327" points="539" reactiontime="+76" swimtime="00:01:18.78" resultid="3385" heatid="4076" lane="7" entrytime="00:01:18.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="378" reactiontime="+78" swimtime="00:00:33.78" resultid="3386" heatid="4087" lane="1" entrytime="00:00:32.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michalina" lastname="Rutkowska" birthdate="2006-01-07" gender="F" nation="POL" license="100305600270" swrid="4949149" athleteid="3343">
              <RESULTS>
                <RESULT eventid="1070" points="477" reactiontime="+82" swimtime="00:00:30.28" resultid="3344" heatid="4021" lane="8" entrytime="00:00:29.72" entrycourse="LCM" />
                <RESULT eventid="1143" points="429" reactiontime="+86" swimtime="00:00:38.97" resultid="3345" heatid="4036" lane="2" entrytime="00:00:39.15" entrycourse="LCM" />
                <RESULT eventid="1281" points="463" reactiontime="+85" swimtime="00:02:25.95" resultid="3346" heatid="4064" lane="0" entrytime="00:02:25.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="336" reactiontime="+79" swimtime="00:00:35.13" resultid="3347" heatid="4082" lane="4" />
                <RESULT eventid="1451" points="489" reactiontime="+79" swimtime="00:01:05.60" resultid="3348" heatid="4103" lane="2" entrytime="00:01:05.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Petrykowska" birthdate="2008-02-19" gender="F" nation="POL" license="100305600236" swrid="5244132" athleteid="3364">
              <RESULTS>
                <RESULT eventid="1070" points="354" reactiontime="+82" swimtime="00:00:33.46" resultid="3365" heatid="4018" lane="3" entrytime="00:00:33.57" entrycourse="LCM" />
                <RESULT eventid="1143" points="418" reactiontime="+88" swimtime="00:00:39.29" resultid="3366" heatid="4036" lane="1" entrytime="00:00:40.10" entrycourse="LCM" />
                <RESULT eventid="1281" points="295" reactiontime="+90" swimtime="00:02:49.71" resultid="3367" heatid="4062" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="100" swimtime="00:01:20.86" />
                    <SPLIT distance="150" swimtime="00:02:06.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1327" points="351" reactiontime="+89" swimtime="00:01:30.83" resultid="3368" heatid="4075" lane="8" entrytime="00:01:28.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="249" reactiontime="+90" swimtime="00:00:38.83" resultid="3369" heatid="4084" lane="5" entrytime="00:00:46.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Górska" birthdate="2005-05-31" gender="F" nation="POL" license="100305600140" swrid="5075861" athleteid="3331">
              <RESULTS>
                <RESULT eventid="1070" points="604" reactiontime="+74" swimtime="00:00:27.99" resultid="3332" heatid="4022" lane="4" entrytime="00:00:28.10" entrycourse="LCM" />
                <RESULT eventid="1235" points="644" reactiontime="+63" swimtime="00:00:31.24" resultid="3333" heatid="4055" lane="5" entrytime="00:00:31.34" entrycourse="LCM" />
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="3334" heatid="4105" lane="6" entrytime="00:01:02.24" entrycourse="LCM" />
                <RESULT eventid="1590" status="DNS" swimtime="00:00:00.00" resultid="3335" heatid="4130" lane="6" entrytime="00:01:08.32" entrycourse="LCM" />
                <RESULT eventid="1728" status="DNS" swimtime="00:00:00.00" resultid="3336" heatid="4152" lane="1" entrytime="00:02:31.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julian" lastname="Pietrowski" birthdate="2008-02-01" gender="M" nation="POL" license="100305700246" swrid="4976715" athleteid="3423">
              <RESULTS>
                <RESULT eventid="1120" points="346" reactiontime="+87" swimtime="00:00:29.76" resultid="3424" heatid="4029" lane="2" entrytime="00:00:30.09" entrycourse="LCM" />
                <RESULT eventid="1212" points="269" reactiontime="+86" swimtime="00:01:16.66" resultid="3425" heatid="4048" lane="6" entrytime="00:01:15.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="283" reactiontime="+87" swimtime="00:02:35.19" resultid="3426" heatid="4069" lane="2" entrytime="00:02:36.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                    <SPLIT distance="100" swimtime="00:01:17.25" />
                    <SPLIT distance="150" swimtime="00:01:58.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="344" reactiontime="+87" swimtime="00:00:31.76" resultid="3427" heatid="4092" lane="0" entrytime="00:00:32.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Lesiński" birthdate="2005-01-16" gender="M" nation="POL" license="100305700179" swrid="4896433" athleteid="3393">
              <RESULTS>
                <RESULT eventid="1120" points="511" reactiontime="+72" swimtime="00:00:26.14" resultid="3394" heatid="4031" lane="2" entrytime="00:00:26.36" entrycourse="LCM" />
                <RESULT eventid="1258" points="493" reactiontime="+67" swimtime="00:00:30.37" resultid="3395" heatid="4060" lane="0" entrytime="00:00:29.62" entrycourse="LCM" />
                <RESULT eventid="1396" points="504" reactiontime="+69" swimtime="00:00:27.97" resultid="3396" heatid="4093" lane="8" entrytime="00:00:28.09" entrycourse="LCM" />
                <RESULT eventid="1613" points="473" reactiontime="+60" swimtime="00:01:06.53" resultid="3397" heatid="4136" lane="9" entrytime="00:01:04.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="452" reactiontime="+60" swimtime="00:02:25.78" resultid="3398" heatid="4155" lane="8" entrytime="00:02:24.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:11.44" />
                    <SPLIT distance="150" swimtime="00:01:49.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Goździk" birthdate="2005-11-07" gender="M" nation="POL" license="100305700176" swrid="5075862" athleteid="3399">
              <RESULTS>
                <RESULT eventid="1120" points="329" reactiontime="+82" swimtime="00:00:30.28" resultid="3400" heatid="4029" lane="5" entrytime="00:00:29.65" entrycourse="LCM" />
                <RESULT eventid="1304" points="334" reactiontime="+88" swimtime="00:02:26.96" resultid="3401" heatid="4070" lane="8" entrytime="00:02:23.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:09.77" />
                    <SPLIT distance="150" swimtime="00:01:49.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="346" reactiontime="+92" swimtime="00:10:43.50" resultid="3402" heatid="4096" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:14.78" />
                    <SPLIT distance="150" swimtime="00:01:55.97" />
                    <SPLIT distance="200" swimtime="00:02:36.60" />
                    <SPLIT distance="250" swimtime="00:03:18.13" />
                    <SPLIT distance="300" swimtime="00:03:59.39" />
                    <SPLIT distance="350" swimtime="00:04:41.53" />
                    <SPLIT distance="400" swimtime="00:05:22.19" />
                    <SPLIT distance="450" swimtime="00:06:03.14" />
                    <SPLIT distance="500" swimtime="00:06:44.16" />
                    <SPLIT distance="550" swimtime="00:07:24.43" />
                    <SPLIT distance="600" swimtime="00:08:05.27" />
                    <SPLIT distance="650" swimtime="00:08:45.26" />
                    <SPLIT distance="700" swimtime="00:09:24.67" />
                    <SPLIT distance="750" swimtime="00:10:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="349" reactiontime="+82" swimtime="00:01:06.60" resultid="3403" heatid="4112" lane="7" entrytime="00:01:06.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="348" reactiontime="+87" swimtime="00:05:12.66" resultid="3404" heatid="4148" lane="2" entrytime="00:05:11.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                    <SPLIT distance="150" swimtime="00:01:54.09" />
                    <SPLIT distance="200" swimtime="00:02:34.39" />
                    <SPLIT distance="250" swimtime="00:03:14.68" />
                    <SPLIT distance="300" swimtime="00:03:54.73" />
                    <SPLIT distance="350" swimtime="00:04:34.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Stefanowski" birthdate="2003-04-03" gender="M" nation="POL" license="100305700152" swrid="4844962" athleteid="3411">
              <RESULTS>
                <RESULT eventid="1120" points="541" reactiontime="+61" swimtime="00:00:25.66" resultid="3412" heatid="4032" lane="8" entrytime="00:00:25.37" entrycourse="LCM" />
                <RESULT eventid="1212" points="637" reactiontime="+66" swimtime="00:00:57.51" resultid="3413" heatid="4050" lane="5" entrytime="00:00:57.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="626" reactiontime="+69" swimtime="00:00:26.03" resultid="3414" heatid="4094" lane="2" entrytime="00:00:26.25" entrycourse="LCM" />
                <RESULT eventid="1567" points="490" reactiontime="+67" swimtime="00:02:20.41" resultid="3415" heatid="4125" lane="6" entrytime="00:02:12.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:05.37" />
                    <SPLIT distance="150" swimtime="00:01:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="546" reactiontime="+62" swimtime="00:04:29.13" resultid="3416" heatid="4149" lane="8" entrytime="00:04:29.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="150" swimtime="00:01:40.45" />
                    <SPLIT distance="200" swimtime="00:02:14.80" />
                    <SPLIT distance="250" swimtime="00:02:49.48" />
                    <SPLIT distance="300" swimtime="00:03:23.91" />
                    <SPLIT distance="350" swimtime="00:03:58.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Dudek" birthdate="2006-11-28" gender="F" nation="POL" license="100305600188" swrid="5195531" athleteid="3472">
              <RESULTS>
                <RESULT eventid="1235" points="546" reactiontime="+62" swimtime="00:00:33.00" resultid="3473" heatid="4054" lane="5" entrytime="00:00:34.18" entrycourse="LCM" />
                <RESULT eventid="1281" points="509" reactiontime="+80" swimtime="00:02:21.44" resultid="3474" heatid="4064" lane="8" entrytime="00:02:23.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:08.30" />
                    <SPLIT distance="150" swimtime="00:01:44.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="454" reactiontime="+74" swimtime="00:00:31.78" resultid="3475" heatid="4086" lane="5" entrytime="00:00:33.88" entrycourse="LCM" />
                <RESULT eventid="1590" points="504" reactiontime="+64" swimtime="00:01:12.34" resultid="3476" heatid="4130" lane="9" entrytime="00:01:13.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="482" reactiontime="+67" swimtime="00:02:37.25" resultid="3477" heatid="4151" lane="4" entrytime="00:02:39.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:17.28" />
                    <SPLIT distance="150" swimtime="00:01:57.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gracjan" lastname="Kostański" birthdate="2005-06-11" gender="M" nation="POL" license="100305700180" swrid="5075869" athleteid="3405">
              <RESULTS>
                <RESULT eventid="1120" points="496" reactiontime="+68" swimtime="00:00:26.40" resultid="3406" heatid="4031" lane="7" entrytime="00:00:26.37" entrycourse="LCM" />
                <RESULT eventid="1166" points="468" reactiontime="+68" swimtime="00:00:33.40" resultid="3407" heatid="4043" lane="1" entrytime="00:00:32.99" entrycourse="LCM" />
                <RESULT eventid="1212" points="418" reactiontime="+69" swimtime="00:01:06.19" resultid="3408" heatid="4049" lane="8" entrytime="00:01:06.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="429" reactiontime="+65" swimtime="00:01:15.38" resultid="3409" heatid="4081" lane="9" entrytime="00:01:15.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="502" reactiontime="+68" swimtime="00:00:58.99" resultid="3410" heatid="4113" lane="2" entrytime="00:01:00.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pola" lastname="Drążkiewicz" birthdate="2007-07-25" gender="F" nation="POL" license="100305600212" swrid="5198017" athleteid="3355">
              <RESULTS>
                <RESULT eventid="1070" points="428" reactiontime="+81" swimtime="00:00:31.40" resultid="3356" heatid="4020" lane="0" entrytime="00:00:30.87" entrycourse="LCM" />
                <RESULT eventid="1143" points="571" reactiontime="+83" swimtime="00:00:35.42" resultid="3357" heatid="4037" lane="2" entrytime="00:00:35.37" entrycourse="LCM" />
                <RESULT eventid="1327" points="541" reactiontime="+83" swimtime="00:01:18.66" resultid="3358" heatid="4076" lane="2" entrytime="00:01:18.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="522" reactiontime="+83" swimtime="00:02:52.69" resultid="3359" heatid="4118" lane="3" entrytime="00:02:52.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                    <SPLIT distance="100" swimtime="00:01:23.46" />
                    <SPLIT distance="150" swimtime="00:02:08.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="418" reactiontime="+94" swimtime="00:05:16.05" resultid="3360" heatid="4144" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:01:55.09" />
                    <SPLIT distance="200" swimtime="00:02:36.55" />
                    <SPLIT distance="250" swimtime="00:03:16.92" />
                    <SPLIT distance="300" swimtime="00:03:57.99" />
                    <SPLIT distance="350" swimtime="00:04:38.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Jankiewicz Delgado" birthdate="2006-06-14" gender="M" nation="POL" license="100305700191" swrid="5075865" athleteid="3325">
              <RESULTS>
                <RESULT eventid="1065" points="420" reactiontime="+81" swimtime="00:05:25.46" resultid="3326" heatid="4013" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:54.99" />
                    <SPLIT distance="200" swimtime="00:02:37.06" />
                    <SPLIT distance="250" swimtime="00:03:23.93" />
                    <SPLIT distance="300" swimtime="00:04:11.39" />
                    <SPLIT distance="350" swimtime="00:04:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="338" reactiontime="+81" swimtime="00:00:37.23" resultid="3327" heatid="4041" lane="2" entrytime="00:00:39.46" entrycourse="LCM" />
                <RESULT eventid="1258" points="342" reactiontime="+69" swimtime="00:00:34.29" resultid="3328" heatid="4059" lane="7" entrytime="00:00:33.50" entrycourse="LCM" />
                <RESULT eventid="1304" points="425" reactiontime="+84" swimtime="00:02:15.60" resultid="3329" heatid="4070" lane="7" entrytime="00:02:17.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                    <SPLIT distance="150" swimtime="00:01:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="436" reactiontime="+83" swimtime="00:09:55.87" resultid="3330" heatid="4097" lane="9" entrytime="00:10:11.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                    <SPLIT distance="150" swimtime="00:01:47.25" />
                    <SPLIT distance="200" swimtime="00:02:25.28" />
                    <SPLIT distance="250" swimtime="00:03:03.03" />
                    <SPLIT distance="300" swimtime="00:03:40.99" />
                    <SPLIT distance="350" swimtime="00:04:19.00" />
                    <SPLIT distance="400" swimtime="00:04:56.93" />
                    <SPLIT distance="450" swimtime="00:05:34.54" />
                    <SPLIT distance="500" swimtime="00:06:12.00" />
                    <SPLIT distance="550" swimtime="00:06:49.56" />
                    <SPLIT distance="600" swimtime="00:07:27.31" />
                    <SPLIT distance="650" swimtime="00:08:04.97" />
                    <SPLIT distance="700" swimtime="00:08:42.18" />
                    <SPLIT distance="750" swimtime="00:09:19.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Michalik" birthdate="2007-10-29" gender="F" nation="POL" license="100305600250" swrid="5303137" athleteid="3434">
              <RESULTS>
                <RESULT eventid="1143" points="440" reactiontime="+79" swimtime="00:00:38.64" resultid="3435" heatid="4037" lane="0" entrytime="00:00:37.97" entrycourse="LCM" />
                <RESULT eventid="1281" points="427" reactiontime="+81" swimtime="00:02:29.99" resultid="3436" heatid="4061" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:12.59" />
                    <SPLIT distance="150" swimtime="00:01:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1327" points="420" reactiontime="+77" swimtime="00:01:25.61" resultid="3437" heatid="4075" lane="4" entrytime="00:01:22.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="424" reactiontime="+78" swimtime="00:03:05.04" resultid="3438" heatid="4118" lane="9" entrytime="00:03:01.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                    <SPLIT distance="100" swimtime="00:01:29.67" />
                    <SPLIT distance="150" swimtime="00:02:19.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="474" reactiontime="+80" swimtime="00:02:41.65" resultid="3439" heatid="4137" lane="5" entrytime="00:02:40.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:16.87" />
                    <SPLIT distance="150" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Celina" lastname="Trzeciak" birthdate="2007-06-20" gender="F" nation="POL" license="100305600241" swrid="4976864" athleteid="3370">
              <RESULTS>
                <RESULT eventid="1070" points="264" reactiontime="+87" swimtime="00:00:36.88" resultid="3371" heatid="4016" lane="4" entrytime="00:00:37.73" entrycourse="LCM" />
                <RESULT eventid="1143" points="250" reactiontime="+77" swimtime="00:00:46.64" resultid="3372" heatid="4035" lane="9" entrytime="00:00:46.58" entrycourse="LCM" />
                <RESULT eventid="1327" points="244" reactiontime="+78" swimtime="00:01:42.57" resultid="3373" heatid="4074" lane="0" entrytime="00:01:42.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="113" reactiontime="+96" swimtime="00:00:50.40" resultid="3374" heatid="4083" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Zakrzewska" birthdate="2007-04-20" gender="F" nation="POL" license="100305600222" swrid="5152529" athleteid="3464">
              <RESULTS>
                <RESULT eventid="1189" points="444" reactiontime="+75" swimtime="00:01:12.68" resultid="3465" heatid="4045" lane="2" entrytime="00:01:13.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="544" reactiontime="+59" swimtime="00:00:33.05" resultid="3466" heatid="4055" lane="8" entrytime="00:00:32.89" entrycourse="LCM" />
                <RESULT eventid="1281" points="469" reactiontime="+73" swimtime="00:02:25.38" resultid="3467" heatid="4061" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:09.58" />
                    <SPLIT distance="150" swimtime="00:01:47.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="546" reactiontime="+60" swimtime="00:01:10.40" resultid="3468" heatid="4130" lane="7" entrytime="00:01:10.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="489" reactiontime="+61" swimtime="00:02:36.55" resultid="3469" heatid="4152" lane="8" entrytime="00:02:36.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:16.92" />
                    <SPLIT distance="150" swimtime="00:01:57.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaja" lastname="Nowak" birthdate="2008-03-30" gender="F" nation="POL" license="100305600233" swrid="4133140" athleteid="3375">
              <RESULTS>
                <RESULT eventid="1070" points="354" reactiontime="+85" swimtime="00:00:33.45" resultid="3376" heatid="4018" lane="9" entrytime="00:00:34.48" entrycourse="LCM" />
                <RESULT eventid="1189" points="228" reactiontime="+73" swimtime="00:01:30.72" resultid="3377" heatid="4044" lane="3" entrytime="00:01:31.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="264" reactiontime="+77" swimtime="00:00:42.05" resultid="3378" heatid="4052" lane="4" entrytime="00:00:43.28" entrycourse="LCM" />
                <RESULT eventid="1281" points="345" reactiontime="+93" swimtime="00:02:40.97" resultid="3379" heatid="4063" lane="0" entrytime="00:02:38.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                    <SPLIT distance="150" swimtime="00:02:00.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="228" reactiontime="+72" swimtime="00:00:39.97" resultid="3380" heatid="4085" lane="7" entrytime="00:00:38.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Rodziewicz" birthdate="2008-01-03" gender="F" nation="POL" license="100305600234" swrid="5198022" athleteid="3387">
              <RESULTS>
                <RESULT eventid="1070" points="540" reactiontime="+62" swimtime="00:00:29.06" resultid="3388" heatid="4015" lane="3" />
                <RESULT eventid="1189" points="570" reactiontime="+69" swimtime="00:01:06.90" resultid="3389" heatid="4046" lane="6" entrytime="00:01:07.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="545" reactiontime="+74" swimtime="00:00:33.01" resultid="3390" heatid="4055" lane="1" entrytime="00:00:32.86" entrycourse="LCM" />
                <RESULT eventid="1281" points="527" reactiontime="+62" swimtime="00:02:19.85" resultid="3391" heatid="4064" lane="9" entrytime="00:02:25.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:44.09" />
                    <SPLIT distance="100" swimtime="00:01:08.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="523" reactiontime="+57" swimtime="00:00:30.31" resultid="3392" heatid="4088" lane="7" entrytime="00:00:30.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Denisiewicz" birthdate="2007-09-24" gender="F" nation="POL" license="100305600272" swrid="5152497" athleteid="3313">
              <RESULTS>
                <RESULT eventid="1060" points="534" reactiontime="+72" swimtime="00:05:28.20" resultid="3314" heatid="4011" lane="8" entrytime="00:05:35.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:17.03" />
                    <SPLIT distance="150" swimtime="00:01:56.62" />
                    <SPLIT distance="200" swimtime="00:02:36.27" />
                    <SPLIT distance="250" swimtime="00:03:22.89" />
                    <SPLIT distance="300" swimtime="00:04:09.26" />
                    <SPLIT distance="350" swimtime="00:04:49.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="450" reactiontime="+72" swimtime="00:01:12.39" resultid="3315" heatid="4045" lane="5" entrytime="00:01:10.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="488" reactiontime="+77" swimtime="00:02:23.46" resultid="3316" heatid="4064" lane="2" entrytime="00:02:21.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:10.29" />
                    <SPLIT distance="150" swimtime="00:01:47.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="565" reactiontime="+70" swimtime="00:02:32.54" resultid="3317" heatid="4138" lane="7" entrytime="00:02:31.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                    <SPLIT distance="150" swimtime="00:01:56.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="531" reactiontime="+61" swimtime="00:02:32.25" resultid="3318" heatid="4152" lane="7" entrytime="00:02:30.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:15.31" />
                    <SPLIT distance="150" swimtime="00:01:54.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Karwat" birthdate="2008-01-12" gender="M" nation="POL" license="100305700235" swrid="5269117" athleteid="3428">
              <RESULTS>
                <RESULT eventid="1120" points="393" reactiontime="+67" swimtime="00:00:28.54" resultid="3429" heatid="4025" lane="2" />
                <RESULT eventid="1212" points="379" reactiontime="+68" swimtime="00:01:08.37" resultid="3430" heatid="4048" lane="4" entrytime="00:01:11.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="418" reactiontime="+67" swimtime="00:00:32.08" resultid="3431" heatid="4059" lane="6" entrytime="00:00:32.81" entrycourse="LCM" />
                <RESULT eventid="1304" points="382" reactiontime="+68" swimtime="00:02:20.50" resultid="3432" heatid="4066" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="150" swimtime="00:01:45.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="390" reactiontime="+66" swimtime="00:00:30.48" resultid="3433" heatid="4092" lane="7" entrytime="00:00:31.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Głowacki" birthdate="2007-02-17" gender="M" nation="POL" license="100305700271" swrid="5230709" athleteid="3440">
              <RESULTS>
                <RESULT eventid="1166" points="378" reactiontime="+70" swimtime="00:00:35.88" resultid="3441" heatid="4042" lane="8" entrytime="00:00:35.90" entrycourse="LCM" />
                <RESULT eventid="1304" points="423" reactiontime="+74" swimtime="00:02:15.86" resultid="3442" heatid="4070" lane="6" entrytime="00:02:16.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:07.30" />
                    <SPLIT distance="150" swimtime="00:01:42.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="409" reactiontime="+76" swimtime="00:01:16.61" resultid="3443" heatid="4080" lane="3" entrytime="00:01:17.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="443" reactiontime="+80" swimtime="00:02:45.32" resultid="3444" heatid="4122" lane="0" entrytime="00:02:44.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:20.62" />
                    <SPLIT distance="150" swimtime="00:02:03.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="417" reactiontime="+72" swimtime="00:04:54.35" resultid="3445" heatid="4148" lane="6" entrytime="00:04:57.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                    <SPLIT distance="200" swimtime="00:02:27.02" />
                    <SPLIT distance="250" swimtime="00:03:04.90" />
                    <SPLIT distance="300" swimtime="00:03:42.71" />
                    <SPLIT distance="350" swimtime="00:04:19.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Ulicka" birthdate="2001-05-16" gender="F" nation="POL" license="100305600206" swrid="4484714" athleteid="3470">
              <RESULTS>
                <RESULT eventid="1235" points="662" reactiontime="+57" swimtime="00:00:30.95" resultid="3471" heatid="4055" lane="4" entrytime="00:00:30.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Świderska" birthdate="2005-08-14" gender="F" nation="POL" license="100305600175" swrid="5075883" athleteid="3452">
              <RESULTS>
                <RESULT eventid="1189" points="585" reactiontime="+81" swimtime="00:01:06.31" resultid="3453" heatid="4046" lane="5" entrytime="00:01:05.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1327" points="377" reactiontime="+84" swimtime="00:01:28.77" resultid="3454" heatid="4075" lane="3" entrytime="00:01:25.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="535" reactiontime="+80" swimtime="00:00:30.08" resultid="3455" heatid="4088" lane="3" entrytime="00:00:29.81" entrycourse="LCM" />
                <RESULT eventid="1544" points="506" reactiontime="+87" swimtime="00:02:32.78" resultid="3456" heatid="4123" lane="3" entrytime="00:02:29.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="150" swimtime="00:01:53.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="443" reactiontime="+91" swimtime="00:02:45.44" resultid="3457" heatid="4138" lane="0" entrytime="00:02:38.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="150" swimtime="00:02:06.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Michalak" birthdate="2003-02-06" gender="M" nation="POL" license="100305700149" swrid="4939878" athleteid="3319">
              <RESULTS>
                <RESULT eventid="1065" points="625" reactiontime="+76" swimtime="00:04:45.08" resultid="3320" heatid="4013" lane="4" entrytime="00:04:40.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                    <SPLIT distance="100" swimtime="00:01:04.38" />
                    <SPLIT distance="150" swimtime="00:01:40.17" />
                    <SPLIT distance="200" swimtime="00:02:17.06" />
                    <SPLIT distance="250" swimtime="00:02:57.97" />
                    <SPLIT distance="300" swimtime="00:03:39.11" />
                    <SPLIT distance="350" swimtime="00:04:12.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="554" reactiontime="+78" swimtime="00:02:04.17" resultid="3321" heatid="4072" lane="0" entrytime="00:02:04.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                    <SPLIT distance="100" swimtime="00:01:01.17" />
                    <SPLIT distance="150" swimtime="00:01:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="511" reactiontime="+76" swimtime="00:00:58.67" resultid="3322" heatid="4109" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="484" reactiontime="+81" swimtime="00:02:40.54" resultid="3323" heatid="4122" lane="3" entrytime="00:02:30.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:16.31" />
                    <SPLIT distance="150" swimtime="00:01:58.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="543" reactiontime="+72" swimtime="00:01:03.55" resultid="3324" heatid="4133" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Furmańska" birthdate="2006-12-16" gender="F" nation="POL" license="100305600186" swrid="5075860" athleteid="3458">
              <RESULTS>
                <RESULT eventid="1189" points="472" reactiontime="+77" swimtime="00:01:11.24" resultid="3459" heatid="4045" lane="6" entrytime="00:01:12.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="492" reactiontime="+84" swimtime="00:02:23.04" resultid="3460" heatid="4064" lane="1" entrytime="00:02:22.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:10.99" />
                    <SPLIT distance="150" swimtime="00:01:48.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="457" reactiontime="+72" swimtime="00:02:38.13" resultid="3461" heatid="4123" lane="7" entrytime="00:02:39.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:57.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="490" reactiontime="+81" swimtime="00:04:59.89" resultid="3462" heatid="4144" lane="4" entrytime="00:05:02.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:11.96" />
                    <SPLIT distance="150" swimtime="00:01:50.32" />
                    <SPLIT distance="200" swimtime="00:02:28.74" />
                    <SPLIT distance="250" swimtime="00:03:07.26" />
                    <SPLIT distance="300" swimtime="00:03:45.60" />
                    <SPLIT distance="350" swimtime="00:04:23.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="473" reactiontime="+85" swimtime="00:10:21.77" resultid="3463" heatid="4157" lane="1" entrytime="00:10:24.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:14.58" />
                    <SPLIT distance="150" swimtime="00:01:54.03" />
                    <SPLIT distance="200" swimtime="00:02:33.50" />
                    <SPLIT distance="250" swimtime="00:03:12.81" />
                    <SPLIT distance="300" swimtime="00:03:51.35" />
                    <SPLIT distance="350" swimtime="00:04:30.40" />
                    <SPLIT distance="400" swimtime="00:05:09.99" />
                    <SPLIT distance="450" swimtime="00:05:49.36" />
                    <SPLIT distance="500" swimtime="00:06:28.73" />
                    <SPLIT distance="550" swimtime="00:07:08.07" />
                    <SPLIT distance="600" swimtime="00:07:47.65" />
                    <SPLIT distance="650" swimtime="00:08:27.04" />
                    <SPLIT distance="700" swimtime="00:09:06.05" />
                    <SPLIT distance="750" swimtime="00:09:44.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02705" nation="POL" region="05" clubid="2827" name="OLIMPIJCZYK Tomaszów Mazowiecki">
          <ATHLETES>
            <ATHLETE firstname="Łucja" lastname="Mielnicka" birthdate="2006-12-29" gender="F" nation="POL" license="102705600062" swrid="4951776" athleteid="2841">
              <RESULTS>
                <RESULT eventid="1070" points="463" reactiontime="+66" swimtime="00:00:30.59" resultid="2842" heatid="4020" lane="9" entrytime="00:00:30.94" entrycourse="LCM" />
                <RESULT eventid="1235" points="487" reactiontime="+74" swimtime="00:00:34.28" resultid="2843" heatid="4054" lane="2" entrytime="00:00:34.56" entrycourse="LCM" />
                <RESULT eventid="1373" points="388" swimtime="00:00:33.48" resultid="2844" heatid="4087" lane="0" entrytime="00:00:33.32" entrycourse="LCM" />
                <RESULT eventid="1590" points="479" reactiontime="+72" swimtime="00:01:13.55" resultid="2845" heatid="4129" lane="5" entrytime="00:01:15.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="418" reactiontime="+72" swimtime="00:02:44.86" resultid="2846" heatid="4151" lane="2" entrytime="00:02:47.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                    <SPLIT distance="100" swimtime="00:01:20.56" />
                    <SPLIT distance="150" swimtime="00:02:03.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Wieczorek" birthdate="2009-09-10" gender="M" nation="POL" license="102705700063" swrid="5253996" athleteid="2866">
              <RESULTS>
                <RESULT eventid="1120" points="299" swimtime="00:00:31.27" resultid="2867" heatid="4029" lane="0" entrytime="00:00:30.76" entrycourse="LCM" />
                <RESULT eventid="1212" points="276" swimtime="00:01:16.01" resultid="2868" heatid="4048" lane="3" entrytime="00:01:14.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="281" reactiontime="+95" swimtime="00:00:33.99" resultid="2869" heatid="4091" lane="4" entrytime="00:00:34.93" entrycourse="LCM" />
                <RESULT eventid="1475" points="334" reactiontime="+72" swimtime="00:01:07.56" resultid="2870" heatid="4111" lane="3" entrytime="00:01:07.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="278" reactiontime="+86" swimtime="00:02:54.57" resultid="2871" heatid="4141" lane="8" entrytime="00:02:55.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                    <SPLIT distance="150" swimtime="00:02:17.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Biernacka" birthdate="2007-07-27" gender="F" nation="POL" license="102705600058" swrid="5214004" athleteid="2828">
              <RESULTS>
                <RESULT eventid="1070" points="527" reactiontime="+79" swimtime="00:00:29.30" resultid="2829" heatid="4021" lane="6" entrytime="00:00:29.48" entrycourse="LCM" />
                <RESULT eventid="1189" points="476" reactiontime="+82" swimtime="00:01:11.03" resultid="2830" heatid="4046" lane="0" entrytime="00:01:08.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="512" reactiontime="+74" swimtime="00:00:30.52" resultid="2831" heatid="4088" lane="2" entrytime="00:00:30.14" entrycourse="LCM" />
                <RESULT eventid="1451" points="520" reactiontime="+79" swimtime="00:01:04.27" resultid="2832" heatid="4103" lane="4" entrytime="00:01:05.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="488" reactiontime="+68" swimtime="00:01:13.09" resultid="2833" heatid="4129" lane="2" entrytime="00:01:18.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Gąsiorowski" birthdate="2009-07-06" gender="M" nation="POL" license="102705700048" swrid="5405807" athleteid="2853">
              <RESULTS>
                <RESULT eventid="1120" points="177" reactiontime="+82" swimtime="00:00:37.22" resultid="2854" heatid="4026" lane="4" entrytime="00:00:35.92" entrycourse="LCM" />
                <RESULT eventid="1166" points="107" reactiontime="+78" swimtime="00:00:54.57" resultid="2855" heatid="4038" lane="7" />
                <RESULT eventid="1258" points="163" reactiontime="+74" swimtime="00:00:43.92" resultid="2856" heatid="4058" lane="9" entrytime="00:00:42.98" entrycourse="LCM" />
                <RESULT eventid="1475" points="177" swimtime="00:01:23.46" resultid="2857" heatid="4109" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="159" reactiontime="+66" swimtime="00:01:35.70" resultid="2858" heatid="4132" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michalina" lastname="Jasińska" birthdate="2006-02-19" gender="F" nation="POL" license="102705600060" swrid="5200924" athleteid="2834">
              <RESULTS>
                <RESULT eventid="1070" points="621" reactiontime="+71" swimtime="00:00:27.74" resultid="2835" heatid="4022" lane="7" entrytime="00:00:28.85" entrycourse="LCM" />
                <RESULT eventid="1235" points="620" reactiontime="+67" swimtime="00:00:31.63" resultid="2836" heatid="4055" lane="2" entrytime="00:00:32.59" entrycourse="LCM" />
                <RESULT eventid="1281" points="565" reactiontime="+84" swimtime="00:02:16.61" resultid="2837" heatid="4065" lane="1" entrytime="00:02:18.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="150" swimtime="00:01:42.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="593" reactiontime="+83" swimtime="00:01:01.52" resultid="2838" heatid="4105" lane="0" entrytime="00:01:03.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="574" reactiontime="+76" swimtime="00:01:09.25" resultid="2839" heatid="4129" lane="4" entrytime="00:01:13.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="512" reactiontime="+66" swimtime="00:02:34.09" resultid="2840" heatid="4152" lane="0" entrytime="00:02:38.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:16.18" />
                    <SPLIT distance="150" swimtime="00:01:55.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Rodzik" birthdate="2007-11-16" gender="F" nation="POL" license="102705600065" swrid="5198060" athleteid="2847">
              <RESULTS>
                <RESULT eventid="1070" points="386" swimtime="00:00:32.49" resultid="2848" heatid="4019" lane="7" entrytime="00:00:31.88" entrycourse="LCM" />
                <RESULT eventid="1143" points="328" swimtime="00:00:42.62" resultid="2849" heatid="4035" lane="5" entrytime="00:00:42.35" entrycourse="LCM" />
                <RESULT eventid="1373" points="356" reactiontime="+72" swimtime="00:00:34.44" resultid="2850" heatid="4086" lane="4" entrytime="00:00:33.85" entrycourse="LCM" />
                <RESULT eventid="1451" points="339" swimtime="00:01:14.11" resultid="2851" heatid="4102" lane="0" entrytime="00:01:11.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="218" reactiontime="+68" swimtime="00:03:22.38" resultid="2852" heatid="4123" lane="1" entrytime="00:03:20.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:24.73" />
                    <SPLIT distance="150" swimtime="00:02:23.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Kowalski" birthdate="2008-10-18" gender="M" nation="POL" license="102705700051" swrid="5356892" athleteid="2859">
              <RESULTS>
                <RESULT eventid="1120" points="264" reactiontime="+83" swimtime="00:00:32.57" resultid="2860" heatid="4027" lane="6" entrytime="00:00:33.32" entrycourse="LCM" />
                <RESULT eventid="1304" points="258" reactiontime="+86" swimtime="00:02:40.15" resultid="2861" heatid="4068" lane="4" entrytime="00:03:03.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:20.35" />
                    <SPLIT distance="150" swimtime="00:02:01.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="167" reactiontime="+84" swimtime="00:00:40.43" resultid="2862" heatid="4090" lane="2" />
                <RESULT eventid="1475" points="269" reactiontime="+85" swimtime="00:01:12.60" resultid="2863" heatid="4110" lane="6" entrytime="00:01:12.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="286" reactiontime="+88" swimtime="00:05:33.85" resultid="2864" heatid="4148" lane="1" entrytime="00:06:02.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:18.36" />
                    <SPLIT distance="150" swimtime="00:02:02.10" />
                    <SPLIT distance="200" swimtime="00:02:45.32" />
                    <SPLIT distance="250" swimtime="00:03:28.34" />
                    <SPLIT distance="300" swimtime="00:04:11.93" />
                    <SPLIT distance="350" swimtime="00:04:54.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="271" reactiontime="+76" swimtime="00:02:52.90" resultid="2865" heatid="4153" lane="4" entrytime="00:03:06.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                    <SPLIT distance="100" swimtime="00:01:27.42" />
                    <SPLIT distance="150" swimtime="00:02:11.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00605" nation="POL" region="05" clubid="3587" name="UKS SP-149 Łódź">
          <ATHLETES>
            <ATHLETE firstname="Kamila" lastname="Haładyn" birthdate="2004-12-02" gender="F" nation="POL" license="100605600389" swrid="5034904" athleteid="3591">
              <RESULTS>
                <RESULT eventid="1060" points="538" reactiontime="+70" swimtime="00:05:27.31" resultid="3592" heatid="4011" lane="7" entrytime="00:05:30.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:10.27" />
                    <SPLIT distance="150" swimtime="00:01:53.44" />
                    <SPLIT distance="200" swimtime="00:02:35.58" />
                    <SPLIT distance="250" swimtime="00:03:24.83" />
                    <SPLIT distance="300" swimtime="00:04:14.30" />
                    <SPLIT distance="350" swimtime="00:04:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="552" reactiontime="+72" swimtime="00:18:41.74" resultid="3593" heatid="4095" lane="3" entrytime="00:18:20.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:09.50" />
                    <SPLIT distance="150" swimtime="00:01:45.75" />
                    <SPLIT distance="200" swimtime="00:02:22.49" />
                    <SPLIT distance="250" swimtime="00:02:59.21" />
                    <SPLIT distance="300" swimtime="00:03:35.91" />
                    <SPLIT distance="350" swimtime="00:04:12.95" />
                    <SPLIT distance="400" swimtime="00:04:49.45" />
                    <SPLIT distance="450" swimtime="00:05:26.50" />
                    <SPLIT distance="500" swimtime="00:06:03.91" />
                    <SPLIT distance="550" swimtime="00:06:41.36" />
                    <SPLIT distance="600" swimtime="00:07:19.41" />
                    <SPLIT distance="650" swimtime="00:07:57.02" />
                    <SPLIT distance="700" swimtime="00:08:34.98" />
                    <SPLIT distance="750" swimtime="00:09:12.69" />
                    <SPLIT distance="800" swimtime="00:09:50.52" />
                    <SPLIT distance="850" swimtime="00:10:28.22" />
                    <SPLIT distance="900" swimtime="00:11:06.14" />
                    <SPLIT distance="950" swimtime="00:11:44.48" />
                    <SPLIT distance="1000" swimtime="00:12:23.11" />
                    <SPLIT distance="1050" swimtime="00:13:01.59" />
                    <SPLIT distance="1100" swimtime="00:13:40.04" />
                    <SPLIT distance="1150" swimtime="00:14:18.54" />
                    <SPLIT distance="1200" swimtime="00:14:57.61" />
                    <SPLIT distance="1250" swimtime="00:15:35.83" />
                    <SPLIT distance="1300" swimtime="00:16:13.92" />
                    <SPLIT distance="1350" swimtime="00:16:52.41" />
                    <SPLIT distance="1400" swimtime="00:17:31.18" />
                    <SPLIT distance="1450" swimtime="00:18:08.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="574" reactiontime="+72" swimtime="00:02:26.51" resultid="3594" heatid="4123" lane="5" entrytime="00:02:26.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:10.05" />
                    <SPLIT distance="150" swimtime="00:01:47.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="565" reactiontime="+71" swimtime="00:04:45.98" resultid="3595" heatid="4145" lane="6" entrytime="00:04:45.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:08.36" />
                    <SPLIT distance="150" swimtime="00:01:44.28" />
                    <SPLIT distance="200" swimtime="00:02:21.29" />
                    <SPLIT distance="250" swimtime="00:02:57.97" />
                    <SPLIT distance="300" swimtime="00:03:35.23" />
                    <SPLIT distance="350" swimtime="00:04:11.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Wentland" birthdate="2007-03-04" gender="M" nation="POL" license="100605700338" swrid="4838034" athleteid="3632">
              <RESULTS>
                <RESULT eventid="1166" points="378" reactiontime="+74" swimtime="00:00:35.88" resultid="3633" heatid="4042" lane="2" entrytime="00:00:35.64" entrycourse="LCM" />
                <RESULT eventid="1350" points="353" reactiontime="+73" swimtime="00:01:20.42" resultid="3634" heatid="4080" lane="2" entrytime="00:01:19.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="385" reactiontime="+68" swimtime="00:00:30.61" resultid="3635" heatid="4092" lane="6" entrytime="00:00:30.55" entrycourse="LCM" />
                <RESULT eventid="1659" points="444" reactiontime="+68" swimtime="00:02:29.37" resultid="3636" heatid="4141" lane="4" entrytime="00:02:31.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="100" swimtime="00:01:09.87" />
                    <SPLIT distance="150" swimtime="00:01:53.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="510" reactiontime="+72" swimtime="00:18:09.94" resultid="3637" heatid="4158" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:46.47" />
                    <SPLIT distance="200" swimtime="00:02:23.70" />
                    <SPLIT distance="250" swimtime="00:03:00.52" />
                    <SPLIT distance="300" swimtime="00:03:38.24" />
                    <SPLIT distance="350" swimtime="00:04:14.98" />
                    <SPLIT distance="400" swimtime="00:04:52.09" />
                    <SPLIT distance="450" swimtime="00:05:28.36" />
                    <SPLIT distance="500" swimtime="00:06:05.91" />
                    <SPLIT distance="550" swimtime="00:06:42.64" />
                    <SPLIT distance="600" swimtime="00:07:19.68" />
                    <SPLIT distance="650" swimtime="00:07:56.21" />
                    <SPLIT distance="700" swimtime="00:08:33.21" />
                    <SPLIT distance="750" swimtime="00:09:10.07" />
                    <SPLIT distance="800" swimtime="00:09:46.67" />
                    <SPLIT distance="850" swimtime="00:10:22.39" />
                    <SPLIT distance="900" swimtime="00:10:59.05" />
                    <SPLIT distance="950" swimtime="00:11:35.79" />
                    <SPLIT distance="1000" swimtime="00:12:12.54" />
                    <SPLIT distance="1050" swimtime="00:12:48.71" />
                    <SPLIT distance="1100" swimtime="00:13:25.25" />
                    <SPLIT distance="1150" swimtime="00:14:01.61" />
                    <SPLIT distance="1200" swimtime="00:14:37.81" />
                    <SPLIT distance="1250" swimtime="00:15:14.00" />
                    <SPLIT distance="1300" swimtime="00:15:50.07" />
                    <SPLIT distance="1350" swimtime="00:16:25.61" />
                    <SPLIT distance="1400" swimtime="00:17:01.82" />
                    <SPLIT distance="1450" swimtime="00:17:36.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Polińska" birthdate="2007-03-28" gender="F" nation="POL" license="100605600346" swrid="4837139" athleteid="3669">
              <RESULTS>
                <RESULT eventid="1235" points="369" reactiontime="+95" swimtime="00:00:37.59" resultid="3670" heatid="4054" lane="0" entrytime="00:00:37.12" entrycourse="LCM" />
                <RESULT eventid="1281" points="357" reactiontime="+84" swimtime="00:02:39.12" resultid="3671" heatid="4062" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:01:59.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="354" reactiontime="+49" swimtime="00:02:54.35" resultid="3672" heatid="4151" lane="1" entrytime="00:02:52.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                    <SPLIT distance="100" swimtime="00:01:26.27" />
                    <SPLIT distance="150" swimtime="00:02:11.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="351" reactiontime="+84" swimtime="00:11:26.71" resultid="3673" heatid="4157" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:21.09" />
                    <SPLIT distance="150" swimtime="00:02:04.39" />
                    <SPLIT distance="200" swimtime="00:02:48.22" />
                    <SPLIT distance="250" swimtime="00:03:32.03" />
                    <SPLIT distance="300" swimtime="00:04:16.17" />
                    <SPLIT distance="350" swimtime="00:05:00.07" />
                    <SPLIT distance="400" swimtime="00:05:43.90" />
                    <SPLIT distance="450" swimtime="00:06:27.77" />
                    <SPLIT distance="500" swimtime="00:07:11.48" />
                    <SPLIT distance="550" swimtime="00:07:55.08" />
                    <SPLIT distance="600" swimtime="00:08:39.04" />
                    <SPLIT distance="650" swimtime="00:09:20.97" />
                    <SPLIT distance="700" swimtime="00:10:04.97" />
                    <SPLIT distance="750" swimtime="00:10:47.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Czerbniak" birthdate="2008-11-21" gender="M" nation="POL" license="100605700393" swrid="5353540" athleteid="3619">
              <RESULTS>
                <RESULT eventid="1120" points="244" reactiontime="+73" swimtime="00:00:33.46" resultid="3620" heatid="4027" lane="3" entrytime="00:00:33.25" entrycourse="LCM" />
                <RESULT eventid="1212" points="232" reactiontime="+91" swimtime="00:01:20.54" resultid="3621" heatid="4048" lane="8" entrytime="00:01:26.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="260" reactiontime="+88" swimtime="00:02:39.64" resultid="3622" heatid="4069" lane="1" entrytime="00:02:39.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:18.11" />
                    <SPLIT distance="150" swimtime="00:02:00.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="227" reactiontime="+74" swimtime="00:01:24.99" resultid="3623" heatid="4134" lane="3" entrytime="00:01:23.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="245" reactiontime="+93" swimtime="00:03:01.94" resultid="3624" heatid="4141" lane="0" entrytime="00:03:00.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:25.06" />
                    <SPLIT distance="150" swimtime="00:02:21.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Rutkowska" birthdate="2007-02-03" gender="F" nation="POL" license="100605600336" swrid="5159189" athleteid="3601">
              <RESULTS>
                <RESULT eventid="1070" points="522" reactiontime="+72" swimtime="00:00:29.38" resultid="3602" heatid="4021" lane="5" entrytime="00:00:29.42" entrycourse="LCM" />
                <RESULT eventid="1281" points="463" reactiontime="+76" swimtime="00:02:26.02" resultid="3603" heatid="4064" lane="4" entrytime="00:02:19.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="150" swimtime="00:01:47.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="523" reactiontime="+81" swimtime="00:01:04.17" resultid="3604" heatid="4104" lane="2" entrytime="00:01:04.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="450" reactiontime="+77" swimtime="00:05:08.40" resultid="3605" heatid="4144" lane="5" entrytime="00:05:05.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                    <SPLIT distance="150" swimtime="00:01:52.16" />
                    <SPLIT distance="200" swimtime="00:02:31.70" />
                    <SPLIT distance="250" swimtime="00:03:11.55" />
                    <SPLIT distance="300" swimtime="00:03:51.14" />
                    <SPLIT distance="350" swimtime="00:04:30.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Porada" birthdate="2008-04-16" gender="M" nation="POL" license="100605700366" swrid="5094196" athleteid="3644">
              <RESULTS>
                <RESULT eventid="1212" points="308" reactiontime="+84" swimtime="00:01:13.22" resultid="3645" heatid="4048" lane="5" entrytime="00:01:13.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="275" swimtime="00:01:27.42" resultid="3646" heatid="4079" lane="5" entrytime="00:01:25.14" entrycourse="LCM" />
                <RESULT eventid="1396" points="265" reactiontime="+87" swimtime="00:00:34.64" resultid="3647" heatid="4089" lane="3" />
                <RESULT eventid="1521" points="334" reactiontime="+91" swimtime="00:03:01.67" resultid="3648" heatid="4121" lane="1" entrytime="00:03:04.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:01:29.27" />
                    <SPLIT distance="150" swimtime="00:02:15.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="345" reactiontime="+98" swimtime="00:05:13.56" resultid="3649" heatid="4147" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:17.28" />
                    <SPLIT distance="150" swimtime="00:01:57.34" />
                    <SPLIT distance="200" swimtime="00:02:37.61" />
                    <SPLIT distance="250" swimtime="00:03:17.33" />
                    <SPLIT distance="300" swimtime="00:03:57.08" />
                    <SPLIT distance="350" swimtime="00:04:36.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Albert" lastname="Ferraretto" birthdate="2008-08-02" gender="M" nation="POL" license="100605700373" swrid="4977094" athleteid="3684">
              <RESULTS>
                <RESULT eventid="1258" points="183" reactiontime="+62" swimtime="00:00:42.23" resultid="3685" heatid="4057" lane="5" entrytime="00:00:43.50" entrycourse="LCM" />
                <RESULT eventid="1304" points="246" reactiontime="+56" swimtime="00:02:42.58" resultid="3686" heatid="4069" lane="9" entrytime="00:02:50.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                    <SPLIT distance="100" swimtime="00:01:21.80" />
                    <SPLIT distance="150" swimtime="00:02:04.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="124" reactiontime="+57" swimtime="00:00:44.60" resultid="3687" heatid="4091" lane="9" entrytime="00:00:45.27" entrycourse="LCM" />
                <RESULT eventid="1705" points="291" reactiontime="+65" swimtime="00:05:31.94" resultid="3688" heatid="4148" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:04.02" />
                    <SPLIT distance="200" swimtime="00:02:46.65" />
                    <SPLIT distance="250" swimtime="00:03:28.97" />
                    <SPLIT distance="300" swimtime="00:04:11.66" />
                    <SPLIT distance="350" swimtime="00:04:53.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Drelich" birthdate="2009-02-09" gender="M" nation="POL" license="100605700394" swrid="5254133" athleteid="3657">
              <RESULTS>
                <RESULT eventid="1212" points="232" reactiontime="+49" swimtime="00:01:20.55" resultid="3658" heatid="4048" lane="7" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="248" reactiontime="+62" swimtime="00:00:38.18" resultid="3659" heatid="4056" lane="0" />
                <RESULT eventid="1350" points="255" swimtime="00:01:29.68" resultid="3660" heatid="4079" lane="1" entrytime="00:01:30.98" entrycourse="LCM" />
                <RESULT eventid="1396" points="223" reactiontime="+55" swimtime="00:00:36.72" resultid="3661" heatid="4090" lane="9" />
                <RESULT eventid="1613" points="257" reactiontime="+61" swimtime="00:01:21.53" resultid="3662" heatid="4134" lane="4" entrytime="00:01:21.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="298" reactiontime="+52" swimtime="00:03:08.70" resultid="4009" heatid="4121" lane="8" entrytime="00:03:07.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:32.74" />
                    <SPLIT distance="150" swimtime="00:02:20.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="293" reactiontime="+61" swimtime="00:02:48.36" resultid="4010" heatid="4154" lane="7" entrytime="00:02:48.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:24.30" />
                    <SPLIT distance="150" swimtime="00:02:07.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Grabarczyk" birthdate="2008-05-30" gender="F" nation="POL" license="100605600360" swrid="5096073" athleteid="3663">
              <RESULTS>
                <RESULT eventid="1235" points="437" reactiontime="+66" swimtime="00:00:35.53" resultid="3664" heatid="4054" lane="8" entrytime="00:00:36.15" entrycourse="LCM" />
                <RESULT eventid="1281" points="417" reactiontime="+71" swimtime="00:02:31.19" resultid="3665" heatid="4063" lane="7" entrytime="00:02:33.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:14.70" />
                    <SPLIT distance="150" swimtime="00:01:53.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="297" reactiontime="+74" swimtime="00:00:36.58" resultid="3666" heatid="4084" lane="6" />
                <RESULT eventid="1590" points="462" reactiontime="+67" swimtime="00:01:14.47" resultid="3667" heatid="4129" lane="6" entrytime="00:01:16.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="483" reactiontime="+76" swimtime="00:02:37.15" resultid="3668" heatid="4151" lane="6" entrytime="00:02:45.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                    <SPLIT distance="150" swimtime="00:01:59.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Rudnicka" birthdate="2009-10-19" gender="F" nation="POL" license="100605600398" swrid="4976834" athleteid="3679">
              <RESULTS>
                <RESULT eventid="1235" points="187" swimtime="00:00:47.16" resultid="3680" heatid="4052" lane="3" entrytime="00:00:47.07" entrycourse="LCM" />
                <RESULT eventid="1281" points="268" swimtime="00:02:55.12" resultid="3681" heatid="4062" lane="6" entrytime="00:03:01.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:01:26.03" />
                    <SPLIT distance="150" swimtime="00:02:10.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="239" swimtime="00:01:23.29" resultid="3682" heatid="4100" lane="6" entrytime="00:01:24.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="267" swimtime="00:06:06.82" resultid="3683" heatid="4144" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:01:27.05" />
                    <SPLIT distance="150" swimtime="00:02:14.33" />
                    <SPLIT distance="200" swimtime="00:03:01.90" />
                    <SPLIT distance="250" swimtime="00:03:48.08" />
                    <SPLIT distance="300" swimtime="00:04:34.97" />
                    <SPLIT distance="350" swimtime="00:05:20.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Mikołajczyk" birthdate="2004-04-16" gender="F" nation="POL" license="100605600245" swrid="4934154" athleteid="3588">
              <RESULTS>
                <RESULT eventid="1060" points="611" reactiontime="+72" swimtime="00:05:13.84" resultid="3589" heatid="4011" lane="6" entrytime="00:05:15.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:12.32" />
                    <SPLIT distance="150" swimtime="00:01:54.08" />
                    <SPLIT distance="200" swimtime="00:02:35.19" />
                    <SPLIT distance="250" swimtime="00:03:19.75" />
                    <SPLIT distance="300" swimtime="00:04:03.07" />
                    <SPLIT distance="350" swimtime="00:04:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="558" reactiontime="+77" swimtime="00:02:27.95" resultid="3590" heatid="4123" lane="6" entrytime="00:02:30.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:11.95" />
                    <SPLIT distance="150" swimtime="00:01:50.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Thim" birthdate="2008-12-18" gender="M" nation="POL" license="100605700379" swrid="5254074" athleteid="3650">
              <RESULTS>
                <RESULT eventid="1212" points="160" reactiontime="+74" swimtime="00:01:31.05" resultid="3651" heatid="4048" lane="0" entrytime="00:01:47.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="233" reactiontime="+77" swimtime="00:00:39.00" resultid="3652" heatid="4058" lane="8" entrytime="00:00:41.83" entrycourse="LCM" />
                <RESULT eventid="1396" points="145" reactiontime="+80" swimtime="00:00:42.35" resultid="3653" heatid="4090" lane="4" entrytime="00:00:46.48" entrycourse="LCM" />
                <RESULT eventid="1613" points="233" reactiontime="+68" swimtime="00:01:24.26" resultid="3654" heatid="4134" lane="7" entrytime="00:01:32.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="199" reactiontime="+82" swimtime="00:03:15.17" resultid="3655" heatid="4140" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="100" swimtime="00:01:34.06" />
                    <SPLIT distance="150" swimtime="00:02:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="259" reactiontime="+68" swimtime="00:02:55.45" resultid="3656" heatid="4153" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="100" swimtime="00:01:27.99" />
                    <SPLIT distance="150" swimtime="00:02:13.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Patyra" birthdate="2009-08-21" gender="F" nation="POL" license="100605600416" swrid="5356901" athleteid="3625">
              <RESULTS>
                <RESULT eventid="1143" points="283" reactiontime="+89" swimtime="00:00:44.78" resultid="3626" heatid="4035" lane="8" entrytime="00:00:45.52" entrycourse="LCM" />
                <RESULT eventid="1235" points="215" swimtime="00:00:44.99" resultid="3627" heatid="4052" lane="2" />
                <RESULT eventid="1327" points="286" reactiontime="+88" swimtime="00:01:37.31" resultid="3628" heatid="4074" lane="6" entrytime="00:01:35.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="225" reactiontime="+75" swimtime="00:01:25.00" resultid="3629" heatid="4098" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="310" reactiontime="+69" swimtime="00:03:25.40" resultid="3630" heatid="4117" lane="7" entrytime="00:03:18.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="100" swimtime="00:01:38.15" />
                    <SPLIT distance="150" swimtime="00:02:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="264" reactiontime="+84" swimtime="00:03:16.36" resultid="3631" heatid="4137" lane="7" entrytime="00:03:20.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                    <SPLIT distance="100" swimtime="00:01:37.39" />
                    <SPLIT distance="150" swimtime="00:02:30.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Rutkowska" birthdate="2009-09-30" gender="F" nation="POL" license="100605600417" swrid="5269131" athleteid="3606">
              <RESULTS>
                <RESULT eventid="1070" points="502" reactiontime="+68" swimtime="00:00:29.77" resultid="3607" heatid="4019" lane="6" entrytime="00:00:31.46" entrycourse="LCM" />
                <RESULT eventid="1189" points="463" reactiontime="+63" swimtime="00:01:11.67" resultid="3608" heatid="4045" lane="7" entrytime="00:01:14.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="469" reactiontime="+66" swimtime="00:02:25.40" resultid="3609" heatid="4063" lane="2" entrytime="00:02:30.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:12.40" />
                    <SPLIT distance="150" swimtime="00:01:50.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="436" reactiontime="+61" swimtime="00:00:32.21" resultid="3610" heatid="4087" lane="9" entrytime="00:00:33.49" entrycourse="LCM" />
                <RESULT eventid="1451" points="499" reactiontime="+60" swimtime="00:01:05.17" resultid="3611" heatid="4103" lane="7" entrytime="00:01:05.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="483" reactiontime="+64" swimtime="00:05:01.36" resultid="3612" heatid="4143" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:12.02" />
                    <SPLIT distance="150" swimtime="00:01:50.68" />
                    <SPLIT distance="200" swimtime="00:02:29.70" />
                    <SPLIT distance="250" swimtime="00:03:08.49" />
                    <SPLIT distance="300" swimtime="00:03:47.68" />
                    <SPLIT distance="350" swimtime="00:04:25.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Jekiel" birthdate="2009-06-05" gender="F" nation="POL" license="100605600395" swrid="5254045" athleteid="3613">
              <RESULTS>
                <RESULT eventid="1070" points="347" reactiontime="+65" swimtime="00:00:33.68" resultid="3614" heatid="4018" lane="6" entrytime="00:00:33.75" entrycourse="LCM" />
                <RESULT eventid="1235" points="309" reactiontime="+91" swimtime="00:00:39.88" resultid="3615" heatid="4053" lane="8" entrytime="00:00:42.03" entrycourse="LCM" />
                <RESULT eventid="1373" points="304" reactiontime="+71" swimtime="00:00:36.32" resultid="3616" heatid="4085" lane="2" entrytime="00:00:37.97" entrycourse="LCM" />
                <RESULT eventid="1451" points="347" reactiontime="+73" swimtime="00:01:13.54" resultid="3617" heatid="4102" lane="9" entrytime="00:01:11.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="312" reactiontime="+95" swimtime="00:01:24.87" resultid="3618" heatid="4128" lane="4" entrytime="00:01:23.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anika" lastname="Łuczak" birthdate="2009-02-12" gender="F" nation="POL" license="100605600400" swrid="5254097" athleteid="3638">
              <RESULTS>
                <RESULT eventid="1189" points="256" reactiontime="+77" swimtime="00:01:27.35" resultid="3639" heatid="4044" lane="5" entrytime="00:01:26.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="370" reactiontime="+79" swimtime="00:02:37.30" resultid="3640" heatid="4062" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                    <SPLIT distance="150" swimtime="00:01:56.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="254" reactiontime="+85" swimtime="00:00:38.57" resultid="3641" heatid="4085" lane="1" entrytime="00:00:39.61" entrycourse="LCM" />
                <RESULT eventid="1590" points="323" reactiontime="+82" swimtime="00:01:23.86" resultid="3642" heatid="4128" lane="7" entrytime="00:01:25.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="334" reactiontime="+75" swimtime="00:02:57.78" resultid="3643" heatid="4151" lane="9" entrytime="00:03:02.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="100" swimtime="00:01:27.24" />
                    <SPLIT distance="150" swimtime="00:02:13.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Fornal" birthdate="2006-07-05" gender="F" nation="POL" license="100605600308" swrid="5159198" athleteid="3674">
              <RESULTS>
                <RESULT eventid="1235" points="333" reactiontime="+63" swimtime="00:00:38.91" resultid="3675" heatid="4052" lane="8" />
                <RESULT eventid="1373" points="371" reactiontime="+75" swimtime="00:00:33.98" resultid="3676" heatid="4086" lane="7" entrytime="00:00:35.36" entrycourse="LCM" />
                <RESULT eventid="1636" points="413" reactiontime="+77" swimtime="00:02:49.27" resultid="3677" heatid="4137" lane="2" entrytime="00:02:53.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:20.13" />
                    <SPLIT distance="150" swimtime="00:02:10.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="374" reactiontime="+67" swimtime="00:02:51.08" resultid="3678" heatid="4151" lane="7" entrytime="00:02:48.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:01:24.17" />
                    <SPLIT distance="150" swimtime="00:02:08.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Boruszewski" birthdate="2007-06-06" gender="M" nation="POL" license="100605700337" swrid="5159195" athleteid="3596">
              <RESULTS>
                <RESULT eventid="1065" points="505" reactiontime="+80" swimtime="00:05:06.06" resultid="3597" heatid="4013" lane="8" entrytime="00:05:16.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:12.06" />
                    <SPLIT distance="150" swimtime="00:01:51.72" />
                    <SPLIT distance="200" swimtime="00:02:30.29" />
                    <SPLIT distance="250" swimtime="00:03:11.80" />
                    <SPLIT distance="300" swimtime="00:03:55.87" />
                    <SPLIT distance="350" swimtime="00:04:32.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="445" reactiontime="+78" swimtime="00:09:52.18" resultid="3598" heatid="4096" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:12.63" />
                    <SPLIT distance="150" swimtime="00:01:50.40" />
                    <SPLIT distance="200" swimtime="00:02:28.08" />
                    <SPLIT distance="250" swimtime="00:03:05.79" />
                    <SPLIT distance="300" swimtime="00:03:44.10" />
                    <SPLIT distance="350" swimtime="00:04:21.53" />
                    <SPLIT distance="400" swimtime="00:04:59.06" />
                    <SPLIT distance="450" swimtime="00:05:36.69" />
                    <SPLIT distance="500" swimtime="00:06:13.68" />
                    <SPLIT distance="550" swimtime="00:06:50.89" />
                    <SPLIT distance="600" swimtime="00:07:29.26" />
                    <SPLIT distance="650" swimtime="00:08:05.52" />
                    <SPLIT distance="700" swimtime="00:08:41.53" />
                    <SPLIT distance="750" swimtime="00:09:16.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="422" reactiontime="+74" swimtime="00:02:48.07" resultid="3599" heatid="4121" lane="3" entrytime="00:02:56.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:22.94" />
                    <SPLIT distance="150" swimtime="00:02:07.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="488" reactiontime="+77" swimtime="00:18:26.10" resultid="3600" heatid="4158" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:51.51" />
                    <SPLIT distance="100" swimtime="00:01:13.12" />
                    <SPLIT distance="150" swimtime="00:03:06.61" />
                    <SPLIT distance="200" swimtime="00:02:28.97" />
                    <SPLIT distance="250" swimtime="00:04:21.78" />
                    <SPLIT distance="300" swimtime="00:03:44.41" />
                    <SPLIT distance="350" swimtime="00:05:36.09" />
                    <SPLIT distance="400" swimtime="00:04:58.86" />
                    <SPLIT distance="450" swimtime="00:06:49.74" />
                    <SPLIT distance="500" swimtime="00:06:13.02" />
                    <SPLIT distance="550" swimtime="00:08:03.46" />
                    <SPLIT distance="600" swimtime="00:07:26.39" />
                    <SPLIT distance="650" swimtime="00:09:17.61" />
                    <SPLIT distance="700" swimtime="00:08:40.33" />
                    <SPLIT distance="750" swimtime="00:10:31.32" />
                    <SPLIT distance="800" swimtime="00:09:54.47" />
                    <SPLIT distance="850" swimtime="00:11:45.13" />
                    <SPLIT distance="900" swimtime="00:11:08.31" />
                    <SPLIT distance="950" swimtime="00:12:58.85" />
                    <SPLIT distance="1000" swimtime="00:12:21.90" />
                    <SPLIT distance="1050" swimtime="00:14:12.65" />
                    <SPLIT distance="1100" swimtime="00:13:36.10" />
                    <SPLIT distance="1150" swimtime="00:15:25.31" />
                    <SPLIT distance="1200" swimtime="00:14:49.19" />
                    <SPLIT distance="1250" swimtime="00:16:38.18" />
                    <SPLIT distance="1300" swimtime="00:16:02.54" />
                    <SPLIT distance="1350" swimtime="00:17:50.31" />
                    <SPLIT distance="1400" swimtime="00:17:14.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05114" nation="POL" region="14" clubid="3308" name="UKS G-8 Bielany Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Rafał" lastname="Żółtowski" birthdate="2005-08-28" gender="M" nation="POL" license="105114700344" swrid="4993430" athleteid="3309">
              <RESULTS>
                <RESULT eventid="1212" points="460" reactiontime="+81" swimtime="00:01:04.11" resultid="3310" heatid="4047" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="452" reactiontime="+78" swimtime="00:02:12.85" resultid="3311" heatid="4068" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:05.41" />
                    <SPLIT distance="150" swimtime="00:01:39.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01905" nation="POL" region="05" clubid="2643" name="MUKS Wodnik Łask">
          <ATHLETES>
            <ATHLETE firstname="Oliwier" lastname="Piotrowski" birthdate="2009-09-18" gender="M" nation="POL" license="101905700153" swrid="5356893" athleteid="2718">
              <RESULTS>
                <RESULT eventid="1120" points="122" reactiontime="+90" swimtime="00:00:42.09" resultid="2719" heatid="4026" lane="1" entrytime="00:00:42.11" entrycourse="LCM" />
                <RESULT eventid="1166" status="DNS" swimtime="00:00:00.00" resultid="2720" heatid="4039" lane="7" entrytime="00:01:04.05" entrycourse="LCM" />
                <RESULT eventid="1258" points="73" reactiontime="+87" swimtime="00:00:57.34" resultid="2721" heatid="4057" lane="1" entrytime="00:00:54.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Gawlik" birthdate="2008-01-09" gender="M" nation="POL" license="101905700138" swrid="4976794" athleteid="2712">
              <RESULTS>
                <RESULT eventid="1120" points="376" reactiontime="+69" swimtime="00:00:28.96" resultid="2713" heatid="4029" lane="6" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1166" points="323" reactiontime="+69" swimtime="00:00:37.82" resultid="2714" heatid="4041" lane="7" entrytime="00:00:40.08" entrycourse="LCM" />
                <RESULT eventid="1350" points="281" reactiontime="+79" swimtime="00:01:26.77" resultid="2715" heatid="4077" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="389" reactiontime="+68" swimtime="00:01:04.23" resultid="2716" heatid="4111" lane="5" entrytime="00:01:07.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="276" reactiontime="+72" swimtime="00:01:19.60" resultid="2717" heatid="4131" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Romański" birthdate="2007-04-27" gender="M" nation="POL" license="101905700134" swrid="4977187" athleteid="2695">
              <RESULTS>
                <RESULT eventid="1120" points="370" reactiontime="+73" swimtime="00:00:29.12" resultid="2696" heatid="4030" lane="9" entrytime="00:00:29.18" entrycourse="LCM" />
                <RESULT eventid="1166" points="337" reactiontime="+92" swimtime="00:00:37.28" resultid="2697" heatid="4041" lane="5" entrytime="00:00:37.39" entrycourse="LCM" />
                <RESULT eventid="1396" points="337" reactiontime="+77" swimtime="00:00:31.98" resultid="2698" heatid="4092" lane="2" entrytime="00:00:30.97" entrycourse="LCM" />
                <RESULT eventid="1475" points="370" reactiontime="+80" swimtime="00:01:05.31" resultid="2699" heatid="4112" lane="2" entrytime="00:01:04.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="305" reactiontime="+99" swimtime="00:03:07.17" resultid="2700" heatid="4121" lane="2" entrytime="00:02:59.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                    <SPLIT distance="100" swimtime="00:01:30.63" />
                    <SPLIT distance="150" swimtime="00:02:19.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Sysio" birthdate="2004-06-21" gender="F" nation="POL" license="101905600079" swrid="5009631" athleteid="2668">
              <RESULTS>
                <RESULT eventid="1070" points="466" reactiontime="+67" swimtime="00:00:30.51" resultid="2669" heatid="4020" lane="7" entrytime="00:00:30.16" entrycourse="LCM" />
                <RESULT eventid="1235" points="462" reactiontime="+62" swimtime="00:00:34.90" resultid="2670" heatid="4054" lane="7" entrytime="00:00:34.83" entrycourse="LCM" />
                <RESULT eventid="1281" points="435" reactiontime="+85" swimtime="00:02:29.00" resultid="2671" heatid="4062" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:52.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="487" reactiontime="+67" swimtime="00:01:05.69" resultid="2672" heatid="4099" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="433" reactiontime="+62" swimtime="00:01:16.06" resultid="2673" heatid="4127" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Wasielewska" birthdate="2008-06-19" gender="F" nation="POL" license="101905600136" swrid="5254109" athleteid="2650">
              <RESULTS>
                <RESULT eventid="1070" points="292" reactiontime="+84" swimtime="00:00:35.66" resultid="2651" heatid="4017" lane="6" entrytime="00:00:35.49" entrycourse="LCM" />
                <RESULT eventid="1143" points="288" reactiontime="+86" swimtime="00:00:44.51" resultid="2652" heatid="4035" lane="3" entrytime="00:00:42.84" entrycourse="LCM" />
                <RESULT eventid="1451" points="280" reactiontime="+91" swimtime="00:01:18.97" resultid="2653" heatid="4101" lane="2" entrytime="00:01:18.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="296" reactiontime="+91" swimtime="00:03:28.52" resultid="2654" heatid="4117" lane="1" entrytime="00:03:29.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                    <SPLIT distance="100" swimtime="00:01:37.14" />
                    <SPLIT distance="150" swimtime="00:02:32.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Nawrocka" birthdate="2008-06-17" gender="F" nation="POL" license="101905600128" swrid="5179197" athleteid="2644">
              <RESULTS>
                <RESULT eventid="1070" points="325" reactiontime="+44" swimtime="00:00:34.41" resultid="2645" heatid="4018" lane="7" entrytime="00:00:33.87" entrycourse="LCM" />
                <RESULT eventid="1235" points="307" reactiontime="+65" swimtime="00:00:39.96" resultid="2646" heatid="4053" lane="5" entrytime="00:00:38.45" entrycourse="LCM" />
                <RESULT eventid="1281" points="308" swimtime="00:02:47.17" resultid="2647" heatid="4062" lane="5" entrytime="00:02:51.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:21.70" />
                    <SPLIT distance="150" swimtime="00:02:07.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="343" reactiontime="+65" swimtime="00:01:13.83" resultid="2648" heatid="4101" lane="6" entrytime="00:01:15.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="291" reactiontime="+76" swimtime="00:01:26.81" resultid="2649" heatid="4128" lane="1" entrytime="00:01:25.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Ulas" birthdate="2007-05-12" gender="M" nation="POL" license="101905700145" swrid="5128620" athleteid="2701">
              <RESULTS>
                <RESULT eventid="1120" points="425" reactiontime="+78" swimtime="00:00:27.81" resultid="2702" heatid="4030" lane="3" entrytime="00:00:27.41" entrycourse="LCM" />
                <RESULT eventid="1258" points="396" reactiontime="+73" swimtime="00:00:32.67" resultid="2703" heatid="4059" lane="3" entrytime="00:00:31.87" entrycourse="LCM" />
                <RESULT eventid="1396" points="400" reactiontime="+72" swimtime="00:00:30.20" resultid="2704" heatid="4092" lane="3" entrytime="00:00:30.32" entrycourse="LCM" />
                <RESULT eventid="1475" points="468" reactiontime="+80" swimtime="00:01:00.41" resultid="2705" heatid="4113" lane="8" entrytime="00:01:01.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="368" reactiontime="+74" swimtime="00:01:12.29" resultid="2706" heatid="4135" lane="2" entrytime="00:01:13.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Kowal" birthdate="2005-04-25" gender="F" nation="POL" license="101905600071" swrid="5009628" athleteid="2728">
              <RESULTS>
                <RESULT eventid="1143" points="474" reactiontime="+85" swimtime="00:00:37.70" resultid="2729" heatid="4037" lane="8" entrytime="00:00:37.41" entrycourse="LCM" />
                <RESULT eventid="1327" points="454" reactiontime="+87" swimtime="00:01:23.42" resultid="2730" heatid="4076" lane="8" entrytime="00:01:21.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="468" reactiontime="+85" swimtime="00:02:59.05" resultid="2731" heatid="4118" lane="2" entrytime="00:02:55.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                    <SPLIT distance="100" swimtime="00:01:26.84" />
                    <SPLIT distance="150" swimtime="00:02:13.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Jura" birthdate="2009-10-14" gender="F" nation="POL" license="101905600154" swrid="5356898" athleteid="2674">
              <RESULTS>
                <RESULT eventid="1070" points="145" reactiontime="+73" swimtime="00:00:45.04" resultid="2675" heatid="4016" lane="2" entrytime="00:00:43.84" entrycourse="LCM" />
                <RESULT eventid="1235" points="166" reactiontime="+85" swimtime="00:00:49.01" resultid="2676" heatid="4052" lane="6" entrytime="00:00:48.57" entrycourse="LCM" />
                <RESULT comment="M4 - Pływak wykonał nierównoczesne ruchy ramion." eventid="1373" reactiontime="+82" status="DSQ" swimtime="00:01:02.39" resultid="2677" heatid="4083" lane="8" />
                <RESULT eventid="1451" points="128" swimtime="00:01:42.34" resultid="2678" heatid="4100" lane="0" entrytime="00:01:42.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="166" reactiontime="+66" swimtime="00:01:44.62" resultid="2679" heatid="4127" lane="3" entrytime="00:01:46.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Drewicz" birthdate="2009-09-06" gender="F" nation="POL" license="101905600156" swrid="5398853" athleteid="2732">
              <RESULTS>
                <RESULT eventid="1143" points="159" reactiontime="+94" swimtime="00:00:54.21" resultid="2733" heatid="4034" lane="6" entrytime="00:00:53.99" entrycourse="LCM" />
                <RESULT eventid="1327" points="164" reactiontime="+96" swimtime="00:01:57.00" resultid="2734" heatid="4073" lane="4" entrytime="00:02:11.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="185" swimtime="00:04:04.04" resultid="2735" heatid="4116" lane="5" entrytime="00:04:26.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.91" />
                    <SPLIT distance="100" swimtime="00:01:58.62" />
                    <SPLIT distance="150" swimtime="00:03:02.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="114" reactiontime="+76" swimtime="00:01:58.42" resultid="2736" heatid="4126" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Piechowski" birthdate="2008-02-04" gender="M" nation="POL" license="101905700139" swrid="5269106" athleteid="2680">
              <RESULTS>
                <RESULT eventid="1120" points="230" reactiontime="+86" swimtime="00:00:34.10" resultid="2681" heatid="4024" lane="3" />
                <RESULT eventid="1396" points="130" reactiontime="+92" swimtime="00:00:43.85" resultid="2682" heatid="4089" lane="6" />
                <RESULT eventid="1475" points="211" reactiontime="+81" swimtime="00:01:18.76" resultid="2683" heatid="4106" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="148" reactiontime="+89" swimtime="00:01:37.86" resultid="2684" heatid="4132" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Kraćkowska" birthdate="2008-01-15" gender="F" nation="POL" license="101905600158" swrid="5356891" athleteid="2655">
              <RESULTS>
                <RESULT eventid="1070" points="291" reactiontime="+79" swimtime="00:00:35.69" resultid="2656" heatid="4017" lane="5" entrytime="00:00:34.73" entrycourse="LCM" />
                <RESULT eventid="1235" points="272" swimtime="00:00:41.59" resultid="2657" heatid="4053" lane="0" entrytime="00:00:43.19" entrycourse="LCM" />
                <RESULT eventid="1451" points="275" reactiontime="+93" swimtime="00:01:19.47" resultid="2658" heatid="4101" lane="0" entrytime="00:01:19.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="241" swimtime="00:01:32.49" resultid="2659" heatid="4126" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Szubert" birthdate="2009-08-21" gender="F" nation="POL" license="101905600148" swrid="4976729" athleteid="2751">
              <RESULTS>
                <RESULT eventid="1451" points="246" reactiontime="+85" swimtime="00:01:22.48" resultid="2752" heatid="4100" lane="3" entrytime="00:01:22.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="227" swimtime="00:01:34.33" resultid="2753" heatid="4127" lane="4" entrytime="00:01:36.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Grzegorzewski" birthdate="2004-03-07" gender="M" nation="POL" license="101905700101" swrid="5113399" athleteid="2737">
              <RESULTS>
                <RESULT eventid="1166" points="579" reactiontime="+71" swimtime="00:00:31.13" resultid="2738" heatid="4043" lane="5" entrytime="00:00:31.21" entrycourse="LCM" />
                <RESULT eventid="1350" points="524" reactiontime="+76" swimtime="00:01:10.55" resultid="2739" heatid="4081" lane="2" entrytime="00:01:10.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="579" reactiontime="+75" swimtime="00:00:56.26" resultid="2740" heatid="4114" lane="3" entrytime="00:00:56.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Kucharska" birthdate="2008-07-07" gender="F" nation="POL" license="101905600142" swrid="4976933" athleteid="2663">
              <RESULTS>
                <RESULT eventid="1070" points="354" reactiontime="+65" swimtime="00:00:33.43" resultid="2664" heatid="4017" lane="3" entrytime="00:00:35.15" entrycourse="LCM" />
                <RESULT eventid="1235" points="259" reactiontime="+77" swimtime="00:00:42.29" resultid="2665" heatid="4053" lane="9" entrytime="00:00:43.19" entrycourse="LCM" />
                <RESULT eventid="1373" points="224" reactiontime="+65" swimtime="00:00:40.20" resultid="2666" heatid="4085" lane="9" entrytime="00:00:42.16" entrycourse="LCM" />
                <RESULT eventid="1451" points="338" reactiontime="+67" swimtime="00:01:14.17" resultid="2667" heatid="4101" lane="7" entrytime="00:01:18.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Lewandowski" birthdate="2003-10-11" gender="M" nation="POL" license="101905700323" swrid="4982310" athleteid="2707">
              <RESULTS>
                <RESULT eventid="1120" points="520" reactiontime="+78" swimtime="00:00:26.00" resultid="2708" heatid="4025" lane="5" />
                <RESULT eventid="1166" points="416" reactiontime="+83" swimtime="00:00:34.75" resultid="2709" heatid="4038" lane="5" />
                <RESULT eventid="1258" points="400" reactiontime="+86" swimtime="00:00:32.56" resultid="2710" heatid="4057" lane="0" />
                <RESULT eventid="1396" points="449" reactiontime="+85" swimtime="00:00:29.07" resultid="2711" heatid="4090" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Olejnik" birthdate="2009-01-19" gender="M" nation="POL" license="101905700175" swrid="5456467" athleteid="2741">
              <RESULTS>
                <RESULT eventid="1166" points="126" swimtime="00:00:51.71" resultid="2742" heatid="4039" lane="2" entrytime="00:00:54.91" entrycourse="LCM" />
                <RESULT eventid="1350" points="112" reactiontime="+99" swimtime="00:01:57.73" resultid="2743" heatid="4078" lane="0" entrytime="00:02:01.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="134" swimtime="00:04:06.34" resultid="2744" heatid="4120" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.06" />
                    <SPLIT distance="100" swimtime="00:01:58.66" />
                    <SPLIT distance="150" swimtime="00:03:04.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="75" reactiontime="+44" swimtime="00:02:02.80" resultid="2745" heatid="4132" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Makówka" birthdate="2006-09-08" gender="M" nation="POL" license="101905700109" swrid="5195515" athleteid="2754">
              <RESULTS>
                <RESULT eventid="1475" points="274" reactiontime="+75" swimtime="00:01:12.16" resultid="2755" heatid="4110" lane="3" entrytime="00:01:12.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="184" reactiontime="+70" swimtime="00:03:41.50" resultid="2756" heatid="4119" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.99" />
                    <SPLIT distance="100" swimtime="00:01:47.87" />
                    <SPLIT distance="150" swimtime="00:02:45.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Klęk" birthdate="2007-10-21" gender="M" nation="POL" license="101905700178" swrid="4132544" athleteid="2690">
              <RESULTS>
                <RESULT eventid="1120" points="293" swimtime="00:00:31.47" resultid="2691" heatid="4028" lane="8" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1166" points="258" reactiontime="+78" swimtime="00:00:40.73" resultid="2692" heatid="4040" lane="8" entrytime="00:00:45.79" entrycourse="LCM" />
                <RESULT eventid="1396" points="260" reactiontime="+83" swimtime="00:00:34.86" resultid="2693" heatid="4091" lane="7" entrytime="00:00:37.43" entrycourse="LCM" />
                <RESULT eventid="1475" points="295" reactiontime="+79" swimtime="00:01:10.41" resultid="2694" heatid="4110" lane="7" entrytime="00:01:14.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nikola" lastname="Błażejewska" birthdate="2003-01-16" gender="F" nation="POL" license="101905600105" swrid="4982307" athleteid="2722">
              <RESULTS>
                <RESULT eventid="1143" points="661" reactiontime="+68" swimtime="00:00:33.75" resultid="2723" heatid="4037" lane="4" entrytime="00:00:33.88" entrycourse="LCM" />
                <RESULT eventid="1327" points="638" reactiontime="+72" swimtime="00:01:14.46" resultid="2724" heatid="4076" lane="4" entrytime="00:01:14.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="480" reactiontime="+76" swimtime="00:00:31.18" resultid="2725" heatid="4087" lane="4" entrytime="00:00:31.05" entrycourse="LCM" />
                <RESULT eventid="1498" points="574" reactiontime="+80" swimtime="00:02:47.34" resultid="2726" heatid="4118" lane="5" entrytime="00:02:45.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                    <SPLIT distance="100" swimtime="00:01:21.66" />
                    <SPLIT distance="150" swimtime="00:02:05.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="573" reactiontime="+74" swimtime="00:02:31.76" resultid="2727" heatid="4138" lane="6" entrytime="00:02:31.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:13.73" />
                    <SPLIT distance="150" swimtime="00:01:56.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Berbelski" birthdate="2009-04-15" gender="M" nation="POL" license="101905700149" swrid="4955510" athleteid="2685">
              <RESULTS>
                <RESULT eventid="1120" points="155" reactiontime="+83" swimtime="00:00:38.92" resultid="2686" heatid="4025" lane="4" />
                <RESULT eventid="1166" points="119" reactiontime="+79" swimtime="00:00:52.69" resultid="2687" heatid="4039" lane="9" />
                <RESULT eventid="1475" points="169" reactiontime="+58" swimtime="00:01:24.78" resultid="2688" heatid="4106" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="124" reactiontime="+71" swimtime="00:01:43.89" resultid="2689" heatid="4133" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Urban" birthdate="2007-12-17" gender="F" nation="POL" license="101905600120" swrid="5254041" athleteid="2660">
              <RESULTS>
                <RESULT eventid="1070" points="318" reactiontime="+89" swimtime="00:00:34.67" resultid="2661" heatid="4018" lane="1" entrytime="00:00:34.15" entrycourse="LCM" />
                <RESULT eventid="1373" points="210" reactiontime="+85" swimtime="00:00:41.07" resultid="2662" heatid="4085" lane="0" entrytime="00:00:40.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Dębkowska" birthdate="2004-10-31" gender="F" nation="POL" license="101905600068" swrid="5101075" athleteid="2746">
              <RESULTS>
                <RESULT eventid="1189" points="532" reactiontime="+83" swimtime="00:01:08.46" resultid="2747" heatid="4046" lane="1" entrytime="00:01:08.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="479" reactiontime="+76" swimtime="00:00:31.21" resultid="2748" heatid="4088" lane="9" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="1544" points="505" reactiontime="+83" swimtime="00:02:32.95" resultid="2749" heatid="4123" lane="2" entrytime="00:02:34.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:12.59" />
                    <SPLIT distance="150" swimtime="00:01:52.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="533" reactiontime="+78" swimtime="00:02:35.49" resultid="2750" heatid="4138" lane="8" entrytime="00:02:35.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:01:59.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03905" nation="POL" region="05" clubid="2030" name="Champion Tomaszów Maz.">
          <ATHLETES>
            <ATHLETE firstname="Laura" lastname="Stępień" birthdate="2008-01-29" gender="F" nation="POL" license="103905600006" swrid="5356112" athleteid="2041">
              <RESULTS>
                <RESULT eventid="1070" points="359" swimtime="00:00:33.28" resultid="2042" heatid="4019" lane="9" entrytime="00:00:32.75" entrycourse="LCM" />
                <RESULT eventid="1235" points="341" reactiontime="+57" swimtime="00:00:38.60" resultid="2043" heatid="4054" lane="9" entrytime="00:00:37.90" entrycourse="LCM" />
                <RESULT eventid="1373" points="271" reactiontime="+58" swimtime="00:00:37.71" resultid="2044" heatid="4085" lane="6" entrytime="00:00:37.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ada" lastname="Lewandowska" birthdate="2009-12-29" gender="F" nation="POL" license="103905600002" swrid="4977027" athleteid="2037">
              <RESULTS>
                <RESULT eventid="1070" points="499" reactiontime="+55" swimtime="00:00:29.83" resultid="2038" heatid="4021" lane="7" entrytime="00:00:29.64" entrycourse="LCM" />
                <RESULT eventid="1235" points="477" reactiontime="+70" swimtime="00:00:34.51" resultid="2039" heatid="4054" lane="6" entrytime="00:00:34.47" entrycourse="LCM" />
                <RESULT eventid="1373" points="442" reactiontime="+63" swimtime="00:00:32.06" resultid="2040" heatid="4087" lane="6" entrytime="00:00:32.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Świnoga" birthdate="2009-03-05" gender="F" nation="POL" license="103905600001" swrid="5356116" athleteid="2045">
              <RESULTS>
                <RESULT eventid="1070" points="328" reactiontime="+73" swimtime="00:00:34.32" resultid="2046" heatid="4018" lane="2" entrytime="00:00:33.75" entrycourse="LCM" />
                <RESULT eventid="1235" points="282" reactiontime="+66" swimtime="00:00:41.11" resultid="2047" heatid="4051" lane="6" />
                <RESULT eventid="1373" points="206" reactiontime="+74" swimtime="00:00:41.32" resultid="2048" heatid="4085" lane="8" entrytime="00:00:40.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marika" lastname="Lesiewicz" birthdate="2004-06-14" gender="F" nation="POL" license="103905600012" swrid="5175104" athleteid="2031">
              <RESULTS>
                <RESULT eventid="1070" points="522" reactiontime="+69" swimtime="00:00:29.38" resultid="2032" heatid="4022" lane="3" entrytime="00:00:28.69" entrycourse="LCM" />
                <RESULT eventid="1235" points="472" reactiontime="+62" swimtime="00:00:34.65" resultid="2033" heatid="4054" lane="3" entrytime="00:00:34.36" entrycourse="LCM" />
                <RESULT eventid="1373" points="467" reactiontime="+71" swimtime="00:00:31.48" resultid="2034" heatid="4088" lane="0" entrytime="00:00:30.98" entrycourse="LCM" />
                <RESULT eventid="1451" points="508" reactiontime="+65" swimtime="00:01:04.80" resultid="2035" heatid="4104" lane="8" entrytime="00:01:04.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="405" reactiontime="+67" swimtime="00:01:17.75" resultid="2036" heatid="4129" lane="3" entrytime="00:01:15.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01014" nation="POL" region="14" clubid="2156" name="KS ,,1&apos;&apos; Ożarów Mazowiecki">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Sobiecka" birthdate="2006-02-22" gender="F" nation="POL" license="101014600118" swrid="5161554" athleteid="2164">
              <RESULTS>
                <RESULT eventid="1070" points="518" reactiontime="+74" swimtime="00:00:29.47" resultid="2165" heatid="4021" lane="1" entrytime="00:00:29.72" entrycourse="LCM" />
                <RESULT eventid="1235" points="524" reactiontime="+70" swimtime="00:00:33.45" resultid="2166" heatid="4054" lane="4" entrytime="00:00:33.61" entrycourse="LCM" />
                <RESULT eventid="1373" points="434" reactiontime="+73" swimtime="00:00:32.25" resultid="2167" heatid="4087" lane="8" entrytime="00:00:32.85" entrycourse="LCM" />
                <RESULT eventid="1451" points="522" reactiontime="+76" swimtime="00:01:04.19" resultid="2168" heatid="4098" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="477" reactiontime="+75" swimtime="00:01:13.65" resultid="2169" heatid="4130" lane="0" entrytime="00:01:13.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Popow" birthdate="2006-04-09" gender="M" nation="POL" license="101014700117" swrid="5161556" athleteid="2170">
              <RESULTS>
                <RESULT eventid="1258" points="555" reactiontime="+85" swimtime="00:00:29.20" resultid="2171" heatid="4060" lane="2" entrytime="00:00:29.11" entrycourse="LCM" />
                <RESULT eventid="1304" points="487" reactiontime="+76" swimtime="00:02:09.59" resultid="2172" heatid="4068" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:01:01.19" />
                    <SPLIT distance="150" swimtime="00:01:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="477" reactiontime="+82" swimtime="00:00:28.49" resultid="2173" heatid="4090" lane="0" />
                <RESULT eventid="1475" points="536" reactiontime="+81" swimtime="00:00:57.72" resultid="2174" heatid="4107" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="569" reactiontime="+77" swimtime="00:01:02.55" resultid="2175" heatid="4136" lane="8" entrytime="00:01:03.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="471" reactiontime="+85" swimtime="00:04:42.72" resultid="2176" heatid="4146" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:05.64" />
                    <SPLIT distance="150" swimtime="00:01:41.71" />
                    <SPLIT distance="200" swimtime="00:02:18.34" />
                    <SPLIT distance="250" swimtime="00:02:55.28" />
                    <SPLIT distance="300" swimtime="00:03:31.93" />
                    <SPLIT distance="350" swimtime="00:04:08.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Adamczyk" birthdate="2006-04-28" gender="F" nation="POL" license="101014600111" swrid="5056861" athleteid="2157">
              <RESULTS>
                <RESULT eventid="1070" points="568" reactiontime="+78" swimtime="00:00:28.57" resultid="2158" heatid="4022" lane="2" entrytime="00:00:28.82" entrycourse="LCM" />
                <RESULT eventid="1189" points="436" reactiontime="+81" swimtime="00:01:13.15" resultid="2159" heatid="4046" lane="7" entrytime="00:01:08.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="564" reactiontime="+78" swimtime="00:02:16.68" resultid="2160" heatid="4065" lane="5" entrytime="00:02:14.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:05.59" />
                    <SPLIT distance="150" swimtime="00:01:41.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="576" reactiontime="+79" swimtime="00:01:02.13" resultid="2161" heatid="4104" lane="3" entrytime="00:01:04.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="452" reactiontime="+78" swimtime="00:03:01.26" resultid="2162" heatid="4116" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:26.82" />
                    <SPLIT distance="150" swimtime="00:02:13.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="522" reactiontime="+80" swimtime="00:04:53.65" resultid="2163" heatid="4145" lane="7" entrytime="00:04:53.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:48.35" />
                    <SPLIT distance="200" swimtime="00:02:26.11" />
                    <SPLIT distance="250" swimtime="00:03:03.27" />
                    <SPLIT distance="300" swimtime="00:03:40.67" />
                    <SPLIT distance="350" swimtime="00:04:17.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00105" nation="POL" region="05" clubid="2876" name="SKS 137 Delfin Łódź">
          <ATHLETES>
            <ATHLETE firstname="Bianka" lastname="Cieplucha" birthdate="2008-09-06" gender="F" nation="POL" license="100105600297" swrid="5254092" athleteid="2971">
              <RESULTS>
                <RESULT eventid="1143" points="405" reactiontime="+85" swimtime="00:00:39.73" resultid="2972" heatid="4035" lane="1" entrytime="00:00:45.21" entrycourse="LCM" />
                <RESULT eventid="1235" points="422" reactiontime="+80" swimtime="00:00:35.95" resultid="2973" heatid="4054" lane="1" entrytime="00:00:35.96" entrycourse="LCM" />
                <RESULT eventid="1327" points="397" reactiontime="+83" swimtime="00:01:27.21" resultid="2974" heatid="4075" lane="6" entrytime="00:01:25.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2975" heatid="4118" lane="8" entrytime="00:02:58.23" entrycourse="LCM" />
                <RESULT eventid="1728" status="DNS" swimtime="00:00:00.00" resultid="2976" heatid="4151" lane="5" entrytime="00:02:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Jeziorska" birthdate="2007-07-27" gender="F" nation="POL" license="100105600268" swrid="5197990" athleteid="2966">
              <RESULTS>
                <RESULT eventid="1143" points="397" reactiontime="+75" swimtime="00:00:39.97" resultid="2967" heatid="4036" lane="8" entrytime="00:00:40.27" entrycourse="LCM" />
                <RESULT eventid="1327" points="403" reactiontime="+83" swimtime="00:01:26.79" resultid="2968" heatid="4075" lane="1" entrytime="00:01:27.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="363" reactiontime="+85" swimtime="00:00:34.22" resultid="2969" heatid="4086" lane="2" entrytime="00:00:35.36" entrycourse="LCM" />
                <RESULT eventid="1498" points="399" reactiontime="+92" swimtime="00:03:08.82" resultid="2970" heatid="4117" lane="4" entrytime="00:03:06.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                    <SPLIT distance="100" swimtime="00:01:31.65" />
                    <SPLIT distance="150" swimtime="00:02:20.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Augustyniak" birthdate="2009-02-01" gender="F" nation="POL" license="100105600324" swrid="4976654" athleteid="3026">
              <RESULTS>
                <RESULT eventid="1498" points="279" reactiontime="+83" swimtime="00:03:32.64" resultid="3027" heatid="4117" lane="8" entrytime="00:03:30.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.41" />
                    <SPLIT distance="100" swimtime="00:01:43.52" />
                    <SPLIT distance="150" swimtime="00:02:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="202" reactiontime="+78" swimtime="00:01:38.00" resultid="3028" heatid="4126" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Strzemecki" birthdate="2008-06-28" gender="M" nation="POL" license="100105700287" swrid="5254059" athleteid="2920">
              <RESULTS>
                <RESULT eventid="1120" points="279" reactiontime="+82" swimtime="00:00:32.00" resultid="2921" heatid="4025" lane="9" />
                <RESULT eventid="1350" points="251" reactiontime="+78" swimtime="00:01:30.06" resultid="2922" heatid="4077" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="243" reactiontime="+79" swimtime="00:01:15.17" resultid="2923" heatid="4107" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="281" reactiontime="+86" swimtime="00:03:12.46" resultid="2924" heatid="4120" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                    <SPLIT distance="100" swimtime="00:01:33.93" />
                    <SPLIT distance="150" swimtime="00:02:23.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="245" reactiontime="+80" swimtime="00:00:41.46" resultid="4161" heatid="4038" lane="8" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sergiusz" lastname="Foryś" birthdate="2008-04-21" gender="M" nation="POL" license="100105700327" swrid="5398852" athleteid="2993">
              <RESULTS>
                <RESULT eventid="1166" points="201" reactiontime="+83" swimtime="00:00:44.27" resultid="2994" heatid="4039" lane="4" entrytime="00:00:48.15" entrycourse="LCM" />
                <RESULT eventid="1350" points="166" reactiontime="+69" swimtime="00:01:43.32" resultid="2995" heatid="4078" lane="1" entrytime="00:01:49.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="185" reactiontime="+64" swimtime="00:03:41.21" resultid="2996" heatid="4119" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                    <SPLIT distance="100" swimtime="00:01:48.13" />
                    <SPLIT distance="150" swimtime="00:02:48.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Adamczyk" birthdate="2006-08-01" gender="F" nation="POL" license="100105600238" swrid="5159129" athleteid="2877">
              <RESULTS>
                <RESULT eventid="1070" points="547" reactiontime="+78" swimtime="00:00:28.94" resultid="2878" heatid="4022" lane="8" entrytime="00:00:28.95" entrycourse="LCM" />
                <RESULT eventid="1189" points="483" reactiontime="+79" swimtime="00:01:10.70" resultid="2879" heatid="4045" lane="4" entrytime="00:01:09.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="497" reactiontime="+82" swimtime="00:00:30.83" resultid="2880" heatid="4088" lane="1" entrytime="00:00:30.62" entrycourse="LCM" />
                <RESULT eventid="1451" points="506" reactiontime="+76" swimtime="00:01:04.85" resultid="2881" heatid="4104" lane="5" entrytime="00:01:03.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Mikołajczyk" birthdate="2007-06-16" gender="M" nation="POL" license="100105700272" swrid="5197985" athleteid="2960">
              <RESULTS>
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="2961" heatid="4030" lane="2" entrytime="00:00:28.08" entrycourse="LCM" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="2962" heatid="4071" lane="8" entrytime="00:02:13.43" entrycourse="LCM" />
                <RESULT eventid="1446" status="DNS" swimtime="00:00:00.00" resultid="2963" heatid="4097" lane="0" entrytime="00:09:57.94" entrycourse="LCM" />
                <RESULT eventid="1475" status="DNS" swimtime="00:00:00.00" resultid="2964" heatid="4113" lane="1" entrytime="00:01:00.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jagoda" lastname="Krystek" birthdate="2008-11-26" gender="F" nation="POL" license="100105600283" swrid="5264120" athleteid="2977">
              <RESULTS>
                <RESULT eventid="1143" points="373" reactiontime="+73" swimtime="00:00:40.83" resultid="2978" heatid="4036" lane="0" entrytime="00:00:40.87" entrycourse="LCM" />
                <RESULT eventid="1281" points="423" reactiontime="+66" swimtime="00:02:30.41" resultid="2979" heatid="4063" lane="8" entrytime="00:02:37.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1327" points="363" reactiontime="+72" swimtime="00:01:29.86" resultid="2980" heatid="4075" lane="0" entrytime="00:01:28.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="396" reactiontime="+62" swimtime="00:03:09.41" resultid="2981" heatid="4117" lane="3" entrytime="00:03:09.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                    <SPLIT distance="100" swimtime="00:01:33.25" />
                    <SPLIT distance="150" swimtime="00:02:22.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="382" reactiontime="+64" swimtime="00:05:25.74" resultid="2982" heatid="4144" lane="3" entrytime="00:05:39.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:01:57.51" />
                    <SPLIT distance="200" swimtime="00:02:39.52" />
                    <SPLIT distance="250" swimtime="00:03:22.33" />
                    <SPLIT distance="300" swimtime="00:04:04.36" />
                    <SPLIT distance="350" swimtime="00:04:46.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Bazler" birthdate="2009-03-30" gender="M" nation="POL" license="100105700316" swrid="5356104" athleteid="2931">
              <RESULTS>
                <RESULT eventid="1120" points="297" reactiontime="+67" swimtime="00:00:31.31" resultid="2932" heatid="4027" lane="4" entrytime="00:00:32.54" entrycourse="LCM" />
                <RESULT eventid="1258" points="271" reactiontime="+69" swimtime="00:00:37.06" resultid="2933" heatid="4058" lane="3" entrytime="00:00:37.60" entrycourse="LCM" />
                <RESULT eventid="1475" points="303" reactiontime="+69" swimtime="00:01:09.80" resultid="2934" heatid="4108" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="283" reactiontime="+75" swimtime="00:01:18.91" resultid="2935" heatid="4135" lane="0" entrytime="00:01:21.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="279" reactiontime="+68" swimtime="00:02:51.15" resultid="2936" heatid="4154" lane="0" entrytime="00:02:54.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:08.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymoteusz" lastname="Borowski" birthdate="2007-04-21" gender="M" nation="POL" license="100105700280" swrid="5264162" athleteid="2910">
              <RESULTS>
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="2911" heatid="4024" lane="8" />
                <RESULT eventid="1258" status="DNS" swimtime="00:00:00.00" resultid="2912" heatid="4056" lane="4" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="2913" heatid="4067" lane="1" />
                <RESULT eventid="1475" status="DNS" swimtime="00:00:00.00" resultid="2914" heatid="4106" lane="2" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="2915" heatid="4131" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Grocholińska" birthdate="2006-03-28" gender="F" nation="POL" license="100105600345" swrid="5170199" athleteid="2882">
              <RESULTS>
                <RESULT eventid="1070" points="238" reactiontime="+92" swimtime="00:00:38.19" resultid="2883" heatid="4016" lane="5" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1235" points="252" reactiontime="+90" swimtime="00:00:42.70" resultid="2884" heatid="4053" lane="7" entrytime="00:00:40.78" entrycourse="LCM" />
                <RESULT eventid="1451" points="203" reactiontime="+97" swimtime="00:01:27.95" resultid="2885" heatid="4100" lane="2" entrytime="00:01:24.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="225" reactiontime="+94" swimtime="00:01:34.53" resultid="2886" heatid="4128" lane="9" entrytime="00:01:32.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Kowalski" birthdate="2008-06-02" gender="M" nation="POL" license="100105700308" swrid="5334758" athleteid="2916">
              <RESULTS>
                <RESULT eventid="1120" points="209" reactiontime="+81" swimtime="00:00:35.20" resultid="2917" heatid="4024" lane="2" />
                <RESULT eventid="1350" points="165" reactiontime="+79" swimtime="00:01:43.62" resultid="2918" heatid="4077" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="189" reactiontime="+92" swimtime="00:03:39.61" resultid="2919" heatid="4120" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.87" />
                    <SPLIT distance="100" swimtime="00:01:45.66" />
                    <SPLIT distance="150" swimtime="00:02:43.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Gajda" birthdate="2007-06-26" gender="M" nation="POL" license="100105700263" swrid="5159126" athleteid="2948">
              <RESULTS>
                <RESULT eventid="1120" points="487" reactiontime="+79" swimtime="00:00:26.56" resultid="2949" heatid="4031" lane="1" entrytime="00:00:26.53" entrycourse="LCM" />
                <RESULT eventid="1212" points="518" reactiontime="+74" swimtime="00:01:01.61" resultid="2950" heatid="4050" lane="8" entrytime="00:01:01.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="460" reactiontime="+83" swimtime="00:02:12.04" resultid="2951" heatid="4071" lane="0" entrytime="00:02:13.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:41.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="502" reactiontime="+82" swimtime="00:00:28.02" resultid="2952" heatid="4093" lane="1" entrytime="00:00:27.92" entrycourse="LCM" />
                <RESULT eventid="1475" points="523" reactiontime="+77" swimtime="00:00:58.22" resultid="2953" heatid="4114" lane="8" entrytime="00:00:58.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="475" reactiontime="+84" swimtime="00:02:21.87" resultid="2954" heatid="4125" lane="8" entrytime="00:02:19.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:46.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="337" reactiontime="+82" swimtime="00:05:16.01" resultid="4227" heatid="4148" lane="5" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:11.70" />
                    <SPLIT distance="150" swimtime="00:01:52.29" />
                    <SPLIT distance="200" swimtime="00:02:33.97" />
                    <SPLIT distance="250" swimtime="00:03:15.08" />
                    <SPLIT distance="300" swimtime="00:03:57.22" />
                    <SPLIT distance="350" swimtime="00:04:39.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Lesiak" birthdate="2009-08-17" gender="M" nation="POL" license="100105700323" swrid="5254046" athleteid="3003">
              <RESULTS>
                <RESULT eventid="1166" points="270" reactiontime="+84" swimtime="00:00:40.14" resultid="3004" heatid="4038" lane="3" />
                <RESULT eventid="1258" points="273" reactiontime="+85" swimtime="00:00:36.98" resultid="3005" heatid="4056" lane="5" />
                <RESULT eventid="1350" points="280" swimtime="00:01:26.93" resultid="3006" heatid="4079" lane="3" entrytime="00:01:27.19" entrycourse="LCM" />
                <RESULT eventid="1521" points="278" reactiontime="+74" swimtime="00:03:13.18" resultid="3007" heatid="4119" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:01:31.51" />
                    <SPLIT distance="150" swimtime="00:02:22.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="286" reactiontime="+72" swimtime="00:02:52.96" resultid="3008" heatid="4141" lane="7" entrytime="00:02:48.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:21.60" />
                    <SPLIT distance="150" swimtime="00:02:11.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Rozwadowska" birthdate="2009-02-07" gender="F" nation="POL" license="100105600312" swrid="5254131" athleteid="2988">
              <RESULTS>
                <RESULT eventid="1143" points="351" reactiontime="+73" swimtime="00:00:41.66" resultid="2989" heatid="4035" lane="2" entrytime="00:00:43.46" entrycourse="LCM" />
                <RESULT eventid="1327" points="377" reactiontime="+74" swimtime="00:01:28.74" resultid="2990" heatid="4074" lane="5" entrytime="00:01:30.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="384" reactiontime="+80" swimtime="00:03:11.31" resultid="2991" heatid="4117" lane="2" entrytime="00:03:13.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.43" />
                    <SPLIT distance="100" swimtime="00:01:33.29" />
                    <SPLIT distance="150" swimtime="00:02:22.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="349" reactiontime="+86" swimtime="00:02:55.18" resultid="2992" heatid="4150" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="100" swimtime="00:01:26.83" />
                    <SPLIT distance="150" swimtime="00:02:12.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystian" lastname="Mierczyński" birthdate="2008-12-30" gender="M" nation="POL" license="100105700305" swrid="5334764" athleteid="2937">
              <RESULTS>
                <RESULT eventid="1120" points="275" reactiontime="+76" swimtime="00:00:32.14" resultid="2938" heatid="4027" lane="2" entrytime="00:00:33.70" entrycourse="LCM" />
                <RESULT eventid="1304" points="255" reactiontime="+79" swimtime="00:02:40.65" resultid="2939" heatid="4069" lane="8" entrytime="00:02:44.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:19.05" />
                    <SPLIT distance="150" swimtime="00:02:02.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="284" reactiontime="+78" swimtime="00:01:11.32" resultid="2940" heatid="4110" lane="1" entrytime="00:01:15.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="197" reactiontime="+69" swimtime="00:01:29.11" resultid="2941" heatid="4134" lane="9" entrytime="00:01:38.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Woźniak" birthdate="2009-05-12" gender="F" nation="POL" license="100105600313" swrid="5254142" athleteid="3012">
              <RESULTS>
                <RESULT eventid="1189" points="308" reactiontime="+67" swimtime="00:01:22.11" resultid="3013" heatid="4045" lane="1" entrytime="00:01:21.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="299" reactiontime="+75" swimtime="00:00:40.34" resultid="3014" heatid="4053" lane="6" entrytime="00:00:39.82" entrycourse="LCM" />
                <RESULT eventid="1373" points="322" reactiontime="+65" swimtime="00:00:35.63" resultid="3015" heatid="4086" lane="9" entrytime="00:00:35.85" entrycourse="LCM" />
                <RESULT eventid="1590" points="322" reactiontime="+71" swimtime="00:01:23.91" resultid="3016" heatid="4128" lane="3" entrytime="00:01:24.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="280" reactiontime="+84" swimtime="00:06:01.21" resultid="3017" heatid="4143" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:01:27.15" />
                    <SPLIT distance="150" swimtime="00:02:14.01" />
                    <SPLIT distance="200" swimtime="00:03:00.96" />
                    <SPLIT distance="250" swimtime="00:03:47.31" />
                    <SPLIT distance="300" swimtime="00:04:32.93" />
                    <SPLIT distance="350" swimtime="00:05:18.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Lamenta" birthdate="2008-08-06" gender="M" nation="POL" license="100105700307" swrid="5334757" athleteid="2925">
              <RESULTS>
                <RESULT eventid="1120" points="385" reactiontime="+66" swimtime="00:00:28.72" resultid="2926" heatid="4029" lane="3" entrytime="00:00:29.75" entrycourse="LCM" />
                <RESULT eventid="1258" points="372" reactiontime="+76" swimtime="00:00:33.37" resultid="2927" heatid="4059" lane="8" entrytime="00:00:35.08" entrycourse="LCM" />
                <RESULT eventid="1396" points="319" reactiontime="+68" swimtime="00:00:32.59" resultid="2928" heatid="4092" lane="1" entrytime="00:00:32.11" entrycourse="LCM" />
                <RESULT eventid="1613" points="366" reactiontime="+69" swimtime="00:01:12.47" resultid="2929" heatid="4135" lane="7" entrytime="00:01:14.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="364" reactiontime="+69" swimtime="00:02:36.73" resultid="2930" heatid="4154" lane="3" entrytime="00:02:40.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:01:58.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Janczak" birthdate="2009-01-27" gender="F" nation="POL" license="100105600315" swrid="5254151" athleteid="2983">
              <RESULTS>
                <RESULT eventid="1143" points="374" reactiontime="+84" swimtime="00:00:40.77" resultid="2984" heatid="4035" lane="4" entrytime="00:00:41.97" entrycourse="LCM" />
                <RESULT eventid="1327" points="393" reactiontime="+86" swimtime="00:01:27.54" resultid="2985" heatid="4074" lane="4" entrytime="00:01:30.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="372" swimtime="00:03:13.27" resultid="2986" heatid="4117" lane="6" entrytime="00:03:10.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                    <SPLIT distance="100" swimtime="00:01:34.69" />
                    <SPLIT distance="150" swimtime="00:02:24.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="313" swimtime="00:05:47.96" resultid="2987" heatid="4143" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="100" swimtime="00:01:21.83" />
                    <SPLIT distance="150" swimtime="00:02:06.66" />
                    <SPLIT distance="200" swimtime="00:02:51.46" />
                    <SPLIT distance="250" swimtime="00:03:35.92" />
                    <SPLIT distance="300" swimtime="00:04:20.89" />
                    <SPLIT distance="350" swimtime="00:05:05.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Kotulska" birthdate="2008-11-06" gender="F" nation="POL" license="100105600288" swrid="5264166" athleteid="2893">
              <RESULTS>
                <RESULT eventid="1070" points="306" reactiontime="+87" swimtime="00:00:35.09" resultid="2894" heatid="4017" lane="1" entrytime="00:00:36.76" entrycourse="LCM" />
                <RESULT eventid="1143" points="271" reactiontime="+94" swimtime="00:00:45.41" resultid="2895" heatid="4034" lane="5" entrytime="00:00:47.02" entrycourse="LCM" />
                <RESULT eventid="1327" points="271" reactiontime="+90" swimtime="00:01:39.07" resultid="2896" heatid="4073" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="252" reactiontime="+95" swimtime="00:03:40.20" resultid="2897" heatid="4116" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.09" />
                    <SPLIT distance="100" swimtime="00:01:43.41" />
                    <SPLIT distance="150" swimtime="00:02:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="292" reactiontime="+76" swimtime="00:03:05.86" resultid="2898" heatid="4150" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                    <SPLIT distance="100" swimtime="00:01:28.45" />
                    <SPLIT distance="150" swimtime="00:02:17.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymon" lastname="Brzeziński" birthdate="2009-07-15" gender="M" nation="POL" license="100105700317" swrid="5254144" athleteid="3018">
              <RESULTS>
                <RESULT eventid="1258" points="264" reactiontime="+92" swimtime="00:00:37.40" resultid="3019" heatid="4058" lane="1" entrytime="00:00:38.87" entrycourse="LCM" />
                <RESULT eventid="1396" points="210" reactiontime="+82" swimtime="00:00:37.43" resultid="3020" heatid="4091" lane="2" entrytime="00:00:36.94" entrycourse="LCM" />
                <RESULT eventid="1613" points="279" reactiontime="+81" swimtime="00:01:19.28" resultid="3021" heatid="4134" lane="2" entrytime="00:01:24.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="236" reactiontime="+83" swimtime="00:03:01.06" resultid="3022" heatid="4154" lane="9" entrytime="00:03:05.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                    <SPLIT distance="100" swimtime="00:01:32.54" />
                    <SPLIT distance="150" swimtime="00:02:20.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Goniszewski" birthdate="2008-07-26" gender="M" nation="POL" license="100105700286" swrid="5197988" athleteid="2955">
              <RESULTS>
                <RESULT eventid="1120" points="239" reactiontime="+76" swimtime="00:00:33.66" resultid="2956" heatid="4028" lane="0" entrytime="00:00:32.15" entrycourse="LCM" />
                <RESULT eventid="1258" points="217" reactiontime="+80" swimtime="00:00:39.91" resultid="2957" heatid="4058" lane="7" entrytime="00:00:38.56" entrycourse="LCM" />
                <RESULT eventid="1475" points="259" reactiontime="+71" swimtime="00:01:13.52" resultid="2958" heatid="4110" lane="4" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="262" reactiontime="+72" swimtime="00:05:43.67" resultid="2959" heatid="4146" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:01:20.65" />
                    <SPLIT distance="150" swimtime="00:02:03.98" />
                    <SPLIT distance="200" swimtime="00:02:48.50" />
                    <SPLIT distance="250" swimtime="00:03:33.74" />
                    <SPLIT distance="300" swimtime="00:04:18.35" />
                    <SPLIT distance="350" swimtime="00:05:02.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Jałkiewicz" birthdate="2008-01-07" gender="M" nation="POL" license="100105700294" swrid="5197979" athleteid="2997">
              <RESULTS>
                <RESULT eventid="1166" points="343" reactiontime="+70" swimtime="00:00:37.07" resultid="2998" heatid="4041" lane="6" entrytime="00:00:38.67" entrycourse="LCM" />
                <RESULT eventid="1258" points="267" reactiontime="+67" swimtime="00:00:37.25" resultid="2999" heatid="4058" lane="6" entrytime="00:00:37.64" entrycourse="LCM" />
                <RESULT eventid="1350" points="285" swimtime="00:01:26.39" resultid="3000" heatid="4079" lane="6" entrytime="00:01:27.95" entrycourse="LCM" />
                <RESULT eventid="1521" points="290" reactiontime="+75" swimtime="00:03:10.35" resultid="3001" heatid="4121" lane="0" entrytime="00:03:07.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                    <SPLIT distance="100" swimtime="00:01:32.20" />
                    <SPLIT distance="150" swimtime="00:02:22.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="242" reactiontime="+70" swimtime="00:01:23.15" resultid="3002" heatid="4134" lane="5" entrytime="00:01:21.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Kowalska" birthdate="2008-01-03" gender="F" nation="POL" license="100105600293" swrid="5190604" athleteid="3023">
              <RESULTS>
                <RESULT eventid="1451" points="278" reactiontime="+73" swimtime="00:01:19.17" resultid="3024" heatid="4101" lane="9" entrytime="00:01:19.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="298" reactiontime="+86" swimtime="00:05:53.92" resultid="3025" heatid="4143" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:09.79" />
                    <SPLIT distance="200" swimtime="00:02:55.28" />
                    <SPLIT distance="250" swimtime="00:03:41.27" />
                    <SPLIT distance="300" swimtime="00:04:26.89" />
                    <SPLIT distance="350" swimtime="00:05:13.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Lichański" birthdate="2008-04-14" gender="M" nation="POL" license="100105700295" swrid="5197983" athleteid="2942">
              <RESULTS>
                <RESULT eventid="1120" points="287" reactiontime="+68" swimtime="00:00:31.69" resultid="2943" heatid="4028" lane="1" entrytime="00:00:31.82" entrycourse="LCM" />
                <RESULT eventid="1166" points="237" reactiontime="+74" swimtime="00:00:41.89" resultid="2944" heatid="4040" lane="4" entrytime="00:00:42.48" entrycourse="LCM" />
                <RESULT eventid="1396" points="191" reactiontime="+66" swimtime="00:00:38.67" resultid="2945" heatid="4091" lane="5" entrytime="00:00:36.57" entrycourse="LCM" />
                <RESULT eventid="1475" points="294" reactiontime="+66" swimtime="00:01:10.50" resultid="2946" heatid="4111" lane="9" entrytime="00:01:10.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="238" reactiontime="+69" swimtime="00:03:03.82" resultid="2947" heatid="4140" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:30.22" />
                    <SPLIT distance="150" swimtime="00:02:24.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Śliwińska" birthdate="2009-04-17" gender="F" nation="POL" license="100105600320" swrid="5254067" athleteid="2899">
              <RESULTS>
                <RESULT eventid="1070" points="289" reactiontime="+95" swimtime="00:00:35.79" resultid="2900" heatid="4017" lane="0" entrytime="00:00:37.33" entrycourse="LCM" />
                <RESULT eventid="1327" points="245" reactiontime="+97" swimtime="00:01:42.35" resultid="2901" heatid="4073" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="259" reactiontime="+92" swimtime="00:01:21.11" resultid="2902" heatid="4098" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="248" reactiontime="+53" swimtime="00:03:41.25" resultid="2903" heatid="4117" lane="9" entrytime="00:03:42.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.31" />
                    <SPLIT distance="100" swimtime="00:01:47.37" />
                    <SPLIT distance="150" swimtime="00:02:45.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymoteusz" lastname="Ogiński" birthdate="2009-01-23" gender="M" nation="POL" license="100105700319" swrid="5254140" athleteid="3009">
              <RESULTS>
                <RESULT eventid="1166" points="209" reactiontime="+60" swimtime="00:00:43.71" resultid="3010" heatid="4040" lane="3" entrytime="00:00:43.02" entrycourse="LCM" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1350" status="DSQ" swimtime="00:01:37.39" resultid="3011" heatid="4079" lane="8" entrytime="00:01:34.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Płuciennikowska" birthdate="2009-08-25" gender="F" nation="POL" license="100105600314" swrid="5293164" athleteid="2887">
              <RESULTS>
                <RESULT eventid="1070" points="450" reactiontime="+75" swimtime="00:00:30.88" resultid="2888" heatid="4019" lane="5" entrytime="00:00:31.13" entrycourse="LCM" />
                <RESULT eventid="1235" points="355" reactiontime="+87" swimtime="00:00:38.08" resultid="2889" heatid="4053" lane="4" entrytime="00:00:38.19" entrycourse="LCM" />
                <RESULT eventid="1373" points="360" reactiontime="+74" swimtime="00:00:34.33" resultid="2890" heatid="4086" lane="3" entrytime="00:00:34.54" entrycourse="LCM" />
                <RESULT eventid="1590" points="354" reactiontime="+99" swimtime="00:01:21.35" resultid="2891" heatid="4129" lane="0" entrytime="00:01:20.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="352" reactiontime="+85" swimtime="00:02:54.66" resultid="2892" heatid="4150" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="150" swimtime="00:02:12.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Adamczyk" birthdate="2009-08-12" gender="F" nation="POL" license="100105600311" swrid="5214020" athleteid="2904">
              <RESULTS>
                <RESULT eventid="1070" points="309" reactiontime="+79" swimtime="00:00:35.00" resultid="2905" heatid="4017" lane="4" entrytime="00:00:34.57" entrycourse="LCM" />
                <RESULT eventid="1235" points="273" reactiontime="+80" swimtime="00:00:41.57" resultid="2906" heatid="4053" lane="1" entrytime="00:00:40.89" entrycourse="LCM" />
                <RESULT eventid="1281" points="312" swimtime="00:02:46.43" resultid="2907" heatid="4063" lane="9" entrytime="00:02:44.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:04.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="282" reactiontime="+75" swimtime="00:01:27.70" resultid="2908" heatid="4128" lane="8" entrytime="00:01:27.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="309" swimtime="00:05:49.49" resultid="2909" heatid="4143" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:22.31" />
                    <SPLIT distance="150" swimtime="00:02:07.52" />
                    <SPLIT distance="200" swimtime="00:02:53.02" />
                    <SPLIT distance="250" swimtime="00:03:38.25" />
                    <SPLIT distance="300" swimtime="00:04:23.42" />
                    <SPLIT distance="350" swimtime="00:05:07.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01105" nation="POL" region="05" clubid="2258" name="MKS Jedynka Łódź">
          <ATHLETES>
            <ATHLETE firstname="Justyna" lastname="Poznańska" birthdate="2005-12-29" gender="F" nation="POL" license="101105600275" swrid="5014386" athleteid="2259">
              <RESULTS>
                <RESULT eventid="1060" points="666" reactiontime="+76" swimtime="00:05:04.95" resultid="2260" heatid="4011" lane="4" entrytime="00:04:55.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:08.90" />
                    <SPLIT distance="150" swimtime="00:01:47.10" />
                    <SPLIT distance="200" swimtime="00:02:23.60" />
                    <SPLIT distance="250" swimtime="00:03:08.55" />
                    <SPLIT distance="300" swimtime="00:03:54.07" />
                    <SPLIT distance="350" swimtime="00:04:30.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="632" reactiontime="+76" swimtime="00:01:04.63" resultid="2261" heatid="4046" lane="3" entrytime="00:01:05.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="678" reactiontime="+73" swimtime="00:02:08.59" resultid="2262" heatid="4062" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="100" swimtime="00:01:03.36" />
                    <SPLIT distance="150" swimtime="00:01:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1327" points="586" reactiontime="+75" swimtime="00:01:16.60" resultid="2263" heatid="4076" lane="6" entrytime="00:01:17.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="578" reactiontime="+77" swimtime="00:02:46.98" resultid="2264" heatid="4116" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:22.06" />
                    <SPLIT distance="150" swimtime="00:02:04.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="682" reactiontime="+60" swimtime="00:01:05.38" resultid="2265" heatid="4130" lane="4" entrytime="00:01:06.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="622" reactiontime="+74" swimtime="00:02:27.67" resultid="2266" heatid="4138" lane="4" entrytime="00:02:19.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:53.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Rudzki" birthdate="2005-03-05" gender="M" nation="POL" license="101105700131" swrid="5118420" athleteid="2368">
              <RESULTS>
                <RESULT eventid="1120" points="541" reactiontime="+70" swimtime="00:00:25.66" resultid="2369" heatid="4031" lane="3" entrytime="00:00:25.87" entrycourse="LCM" />
                <RESULT eventid="1212" points="482" reactiontime="+76" swimtime="00:01:03.09" resultid="2370" heatid="4049" lane="5" entrytime="00:01:03.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="433" reactiontime="+69" swimtime="00:00:31.70" resultid="2371" heatid="4056" lane="6" />
                <RESULT eventid="1304" points="434" reactiontime="+74" swimtime="00:02:14.64" resultid="2372" heatid="4071" lane="4" entrytime="00:02:08.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                    <SPLIT distance="100" swimtime="00:01:03.15" />
                    <SPLIT distance="150" swimtime="00:01:38.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="530" reactiontime="+71" swimtime="00:00:27.51" resultid="2373" heatid="4093" lane="6" entrytime="00:00:27.50" entrycourse="LCM" />
                <RESULT eventid="1475" points="550" reactiontime="+74" swimtime="00:00:57.25" resultid="2374" heatid="4114" lane="5" entrytime="00:00:56.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="513" reactiontime="+70" swimtime="00:02:22.40" resultid="2375" heatid="4140" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:07.99" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Potemka" birthdate="2004-04-24" gender="F" nation="POL" license="101105600243" swrid="5075840" athleteid="2414">
              <RESULTS>
                <RESULT eventid="1451" points="461" reactiontime="+71" swimtime="00:01:06.92" resultid="2415" heatid="4099" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="477" reactiontime="+75" swimtime="00:05:02.55" resultid="2416" heatid="4143" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:49.13" />
                    <SPLIT distance="200" swimtime="00:02:27.95" />
                    <SPLIT distance="250" swimtime="00:03:06.86" />
                    <SPLIT distance="300" swimtime="00:03:45.88" />
                    <SPLIT distance="350" swimtime="00:04:24.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymoteusz" lastname="Jóźwiak" birthdate="2008-04-27" gender="M" nation="POL" license="101105700278" swrid="5180509" athleteid="2345">
              <RESULTS>
                <RESULT eventid="1120" points="479" reactiontime="+87" swimtime="00:00:26.72" resultid="2346" heatid="4031" lane="0" entrytime="00:00:26.96" entrycourse="LCM" />
                <RESULT eventid="1212" points="535" reactiontime="+80" swimtime="00:01:00.94" resultid="2347" heatid="4050" lane="9" entrytime="00:01:01.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="515" reactiontime="+80" swimtime="00:02:07.23" resultid="2348" heatid="4071" lane="5" entrytime="00:02:09.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                    <SPLIT distance="100" swimtime="00:01:02.14" />
                    <SPLIT distance="150" swimtime="00:01:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="513" reactiontime="+76" swimtime="00:00:27.81" resultid="2349" heatid="4093" lane="7" entrytime="00:00:27.81" entrycourse="LCM" />
                <RESULT eventid="1475" points="511" reactiontime="+81" swimtime="00:00:58.67" resultid="2350" heatid="4114" lane="9" entrytime="00:00:58.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="521" reactiontime="+85" swimtime="00:04:33.48" resultid="2351" heatid="4148" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="150" swimtime="00:01:39.14" />
                    <SPLIT distance="200" swimtime="00:02:14.26" />
                    <SPLIT distance="250" swimtime="00:02:49.45" />
                    <SPLIT distance="300" swimtime="00:03:24.29" />
                    <SPLIT distance="350" swimtime="00:03:59.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marianna" lastname="Oberbecka" birthdate="2006-06-14" gender="F" nation="POL" license="101105600306" swrid="5159152" athleteid="2303">
              <RESULTS>
                <RESULT eventid="1070" points="376" reactiontime="+92" swimtime="00:00:32.79" resultid="2304" heatid="4016" lane="1" />
                <RESULT eventid="1451" points="321" reactiontime="+99" swimtime="00:01:15.50" resultid="2305" heatid="4098" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Arent" birthdate="2005-05-05" gender="M" nation="POL" license="101105700215" swrid="5118473" athleteid="2276">
              <RESULTS>
                <RESULT eventid="1065" points="554" reactiontime="+63" swimtime="00:04:56.75" resultid="2277" heatid="4012" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:08.98" />
                    <SPLIT distance="150" swimtime="00:01:48.69" />
                    <SPLIT distance="200" swimtime="00:02:27.21" />
                    <SPLIT distance="250" swimtime="00:03:07.17" />
                    <SPLIT distance="300" swimtime="00:03:48.55" />
                    <SPLIT distance="350" swimtime="00:04:23.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="487" reactiontime="+66" swimtime="00:02:09.58" resultid="2278" heatid="4072" lane="9" entrytime="00:02:06.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:03.03" />
                    <SPLIT distance="150" swimtime="00:01:36.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="579" reactiontime="+67" swimtime="00:09:02.15" resultid="2279" heatid="4097" lane="6" entrytime="00:09:05.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                    <SPLIT distance="100" swimtime="00:01:05.65" />
                    <SPLIT distance="150" swimtime="00:01:40.23" />
                    <SPLIT distance="200" swimtime="00:02:14.91" />
                    <SPLIT distance="250" swimtime="00:02:49.68" />
                    <SPLIT distance="300" swimtime="00:03:24.20" />
                    <SPLIT distance="350" swimtime="00:03:58.40" />
                    <SPLIT distance="400" swimtime="00:04:33.29" />
                    <SPLIT distance="450" swimtime="00:05:07.41" />
                    <SPLIT distance="500" swimtime="00:05:41.53" />
                    <SPLIT distance="550" swimtime="00:06:15.28" />
                    <SPLIT distance="600" swimtime="00:06:49.19" />
                    <SPLIT distance="650" swimtime="00:07:22.96" />
                    <SPLIT distance="700" swimtime="00:07:56.78" />
                    <SPLIT distance="750" swimtime="00:08:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="546" reactiontime="+71" swimtime="00:02:19.45" resultid="2280" heatid="4140" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:07.61" />
                    <SPLIT distance="150" swimtime="00:01:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="546" reactiontime="+66" swimtime="00:04:29.13" resultid="2281" heatid="4149" lane="7" entrytime="00:04:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:05.67" />
                    <SPLIT distance="150" swimtime="00:01:40.70" />
                    <SPLIT distance="200" swimtime="00:02:15.15" />
                    <SPLIT distance="250" swimtime="00:02:49.16" />
                    <SPLIT distance="300" swimtime="00:03:23.20" />
                    <SPLIT distance="350" swimtime="00:03:57.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="618" reactiontime="+70" swimtime="00:17:02.05" resultid="2282" heatid="4159" lane="3" entrytime="00:17:13.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:06.88" />
                    <SPLIT distance="150" swimtime="00:01:42.11" />
                    <SPLIT distance="200" swimtime="00:02:17.42" />
                    <SPLIT distance="250" swimtime="00:02:52.69" />
                    <SPLIT distance="300" swimtime="00:03:27.80" />
                    <SPLIT distance="350" swimtime="00:04:02.84" />
                    <SPLIT distance="400" swimtime="00:04:37.84" />
                    <SPLIT distance="450" swimtime="00:05:12.46" />
                    <SPLIT distance="500" swimtime="00:05:46.97" />
                    <SPLIT distance="550" swimtime="00:06:21.41" />
                    <SPLIT distance="600" swimtime="00:06:55.76" />
                    <SPLIT distance="650" swimtime="00:07:30.26" />
                    <SPLIT distance="700" swimtime="00:08:04.55" />
                    <SPLIT distance="750" swimtime="00:08:38.71" />
                    <SPLIT distance="800" swimtime="00:09:12.55" />
                    <SPLIT distance="850" swimtime="00:09:46.64" />
                    <SPLIT distance="900" swimtime="00:10:20.45" />
                    <SPLIT distance="950" swimtime="00:10:54.51" />
                    <SPLIT distance="1000" swimtime="00:11:28.07" />
                    <SPLIT distance="1050" swimtime="00:12:02.28" />
                    <SPLIT distance="1100" swimtime="00:12:35.71" />
                    <SPLIT distance="1150" swimtime="00:13:09.39" />
                    <SPLIT distance="1200" swimtime="00:13:42.49" />
                    <SPLIT distance="1250" swimtime="00:14:16.39" />
                    <SPLIT distance="1300" swimtime="00:14:49.56" />
                    <SPLIT distance="1350" swimtime="00:15:23.44" />
                    <SPLIT distance="1400" swimtime="00:15:56.85" />
                    <SPLIT distance="1450" swimtime="00:16:29.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Sztendel" birthdate="2008-05-09" gender="M" nation="POL" license="101105700232" swrid="4976970" athleteid="2340">
              <RESULTS>
                <RESULT eventid="1120" points="284" reactiontime="+81" swimtime="00:00:31.80" resultid="2341" heatid="4025" lane="0" />
                <RESULT eventid="1166" points="283" reactiontime="+77" swimtime="00:00:39.50" resultid="2342" heatid="4041" lane="1" entrytime="00:00:40.85" entrycourse="LCM" />
                <RESULT eventid="1350" points="258" swimtime="00:01:29.30" resultid="2343" heatid="4079" lane="7" entrytime="00:01:30.50" entrycourse="LCM" />
                <RESULT eventid="1521" points="260" reactiontime="+85" swimtime="00:03:17.57" resultid="2344" heatid="4120" lane="4" entrytime="00:03:12.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:35.36" />
                    <SPLIT distance="150" swimtime="00:02:25.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Płoszka" birthdate="2005-12-17" gender="M" nation="POL" license="101105700239" swrid="5075843" athleteid="2376">
              <RESULTS>
                <RESULT eventid="1120" points="590" reactiontime="+73" swimtime="00:00:24.93" resultid="2377" heatid="4032" lane="1" entrytime="00:00:25.25" entrycourse="LCM" />
                <RESULT eventid="1212" points="639" reactiontime="+71" swimtime="00:00:57.44" resultid="2378" heatid="4050" lane="4" entrytime="00:00:56.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="705" reactiontime="+67" swimtime="00:01:54.59" resultid="2379" heatid="4072" lane="4" entrytime="00:01:53.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.12" />
                    <SPLIT distance="100" swimtime="00:00:56.24" />
                    <SPLIT distance="150" swimtime="00:01:26.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="590" reactiontime="+69" swimtime="00:00:26.55" resultid="2380" heatid="4094" lane="6" entrytime="00:00:26.23" entrycourse="LCM" />
                <RESULT eventid="1446" points="666" reactiontime="+69" swimtime="00:08:37.49" resultid="2381" heatid="4097" lane="5" entrytime="00:08:57.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:02.61" />
                    <SPLIT distance="150" swimtime="00:01:35.12" />
                    <SPLIT distance="200" swimtime="00:02:08.14" />
                    <SPLIT distance="250" swimtime="00:02:40.94" />
                    <SPLIT distance="300" swimtime="00:03:13.71" />
                    <SPLIT distance="350" swimtime="00:03:46.41" />
                    <SPLIT distance="400" swimtime="00:04:19.34" />
                    <SPLIT distance="450" swimtime="00:04:51.80" />
                    <SPLIT distance="500" swimtime="00:05:24.63" />
                    <SPLIT distance="550" swimtime="00:05:57.14" />
                    <SPLIT distance="600" swimtime="00:06:30.50" />
                    <SPLIT distance="650" swimtime="00:07:03.02" />
                    <SPLIT distance="700" swimtime="00:07:36.04" />
                    <SPLIT distance="750" swimtime="00:08:08.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="686" reactiontime="+70" swimtime="00:00:53.17" resultid="2382" heatid="4115" lane="8" entrytime="00:00:54.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="644" reactiontime="+69" swimtime="00:02:08.16" resultid="2383" heatid="4125" lane="4" entrytime="00:02:05.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                    <SPLIT distance="100" swimtime="00:01:01.73" />
                    <SPLIT distance="150" swimtime="00:01:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="707" reactiontime="+68" swimtime="00:04:06.97" resultid="2384" heatid="4149" lane="4" entrytime="00:04:07.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                    <SPLIT distance="100" swimtime="00:00:58.12" />
                    <SPLIT distance="150" swimtime="00:02:32.36" />
                    <SPLIT distance="200" swimtime="00:02:00.60" />
                    <SPLIT distance="250" swimtime="00:03:36.87" />
                    <SPLIT distance="300" swimtime="00:03:04.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="681" reactiontime="+70" swimtime="00:16:29.78" resultid="2385" heatid="4159" lane="5" entrytime="00:17:08.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:02.31" />
                    <SPLIT distance="150" swimtime="00:01:35.31" />
                    <SPLIT distance="200" swimtime="00:02:08.50" />
                    <SPLIT distance="250" swimtime="00:02:41.16" />
                    <SPLIT distance="300" swimtime="00:03:14.77" />
                    <SPLIT distance="350" swimtime="00:03:48.34" />
                    <SPLIT distance="400" swimtime="00:04:21.72" />
                    <SPLIT distance="450" swimtime="00:04:54.86" />
                    <SPLIT distance="500" swimtime="00:05:28.56" />
                    <SPLIT distance="550" swimtime="00:06:02.01" />
                    <SPLIT distance="600" swimtime="00:06:35.41" />
                    <SPLIT distance="650" swimtime="00:07:08.45" />
                    <SPLIT distance="700" swimtime="00:07:41.85" />
                    <SPLIT distance="750" swimtime="00:08:15.16" />
                    <SPLIT distance="800" swimtime="00:08:48.32" />
                    <SPLIT distance="850" swimtime="00:09:21.50" />
                    <SPLIT distance="900" swimtime="00:09:54.38" />
                    <SPLIT distance="950" swimtime="00:10:27.12" />
                    <SPLIT distance="1000" swimtime="00:11:00.46" />
                    <SPLIT distance="1050" swimtime="00:11:33.30" />
                    <SPLIT distance="1100" swimtime="00:12:07.20" />
                    <SPLIT distance="1150" swimtime="00:12:41.05" />
                    <SPLIT distance="1200" swimtime="00:13:14.40" />
                    <SPLIT distance="1250" swimtime="00:13:47.76" />
                    <SPLIT distance="1300" swimtime="00:15:27.02" />
                    <SPLIT distance="1350" swimtime="00:14:54.15" />
                    <SPLIT distance="1400" swimtime="00:16:29.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Banasiak" birthdate="2005-07-04" gender="M" nation="POL" license="101105700136" swrid="5118421" athleteid="2359">
              <RESULTS>
                <RESULT eventid="1120" points="518" reactiontime="+69" swimtime="00:00:26.02" resultid="2360" heatid="4032" lane="9" entrytime="00:00:25.52" entrycourse="LCM" />
                <RESULT eventid="1212" points="514" reactiontime="+76" swimtime="00:01:01.77" resultid="2361" heatid="4050" lane="6" entrytime="00:00:59.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="565" reactiontime="+68" swimtime="00:00:26.93" resultid="2362" heatid="4094" lane="7" entrytime="00:00:26.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Mochnal" birthdate="2005-09-11" gender="M" nation="POL" license="101105700240" swrid="4980423" athleteid="2397">
              <RESULTS>
                <RESULT eventid="1212" points="599" reactiontime="+68" swimtime="00:00:58.71" resultid="2398" heatid="4050" lane="2" entrytime="00:00:59.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="558" reactiontime="+66" swimtime="00:02:03.89" resultid="2399" heatid="4072" lane="2" entrytime="00:02:02.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                    <SPLIT distance="100" swimtime="00:00:59.91" />
                    <SPLIT distance="150" swimtime="00:01:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="531" reactiontime="+66" swimtime="00:00:27.50" resultid="2400" heatid="4089" lane="1" />
                <RESULT eventid="1446" points="581" reactiontime="+66" swimtime="00:09:01.70" resultid="2401" heatid="4096" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:40.41" />
                    <SPLIT distance="200" swimtime="00:02:15.17" />
                    <SPLIT distance="250" swimtime="00:02:49.24" />
                    <SPLIT distance="300" swimtime="00:03:23.01" />
                    <SPLIT distance="350" swimtime="00:03:57.22" />
                    <SPLIT distance="400" swimtime="00:04:31.04" />
                    <SPLIT distance="450" swimtime="00:05:05.52" />
                    <SPLIT distance="500" swimtime="00:05:38.86" />
                    <SPLIT distance="550" swimtime="00:06:13.56" />
                    <SPLIT distance="600" swimtime="00:06:47.49" />
                    <SPLIT distance="650" swimtime="00:07:21.99" />
                    <SPLIT distance="700" swimtime="00:07:55.95" />
                    <SPLIT distance="750" swimtime="00:08:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="641" reactiontime="+67" swimtime="00:02:08.37" resultid="2402" heatid="4125" lane="3" entrytime="00:02:07.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:02.27" />
                    <SPLIT distance="150" swimtime="00:01:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="614" reactiontime="+64" swimtime="00:04:18.84" resultid="2403" heatid="4149" lane="6" entrytime="00:04:17.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.20" />
                    <SPLIT distance="100" swimtime="00:01:01.31" />
                    <SPLIT distance="150" swimtime="00:02:41.15" />
                    <SPLIT distance="200" swimtime="00:02:08.26" />
                    <SPLIT distance="250" swimtime="00:03:47.86" />
                    <SPLIT distance="300" swimtime="00:03:15.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="620" reactiontime="+65" swimtime="00:17:01.03" resultid="2404" heatid="4159" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                    <SPLIT distance="100" swimtime="00:01:04.67" />
                    <SPLIT distance="150" swimtime="00:01:38.49" />
                    <SPLIT distance="200" swimtime="00:02:12.77" />
                    <SPLIT distance="250" swimtime="00:02:46.60" />
                    <SPLIT distance="300" swimtime="00:03:21.17" />
                    <SPLIT distance="350" swimtime="00:03:55.03" />
                    <SPLIT distance="400" swimtime="00:04:29.85" />
                    <SPLIT distance="450" swimtime="00:05:03.77" />
                    <SPLIT distance="500" swimtime="00:05:38.34" />
                    <SPLIT distance="550" swimtime="00:06:12.64" />
                    <SPLIT distance="600" swimtime="00:06:47.16" />
                    <SPLIT distance="650" swimtime="00:07:21.32" />
                    <SPLIT distance="700" swimtime="00:07:55.95" />
                    <SPLIT distance="750" swimtime="00:08:30.28" />
                    <SPLIT distance="800" swimtime="00:09:04.96" />
                    <SPLIT distance="850" swimtime="00:09:39.30" />
                    <SPLIT distance="900" swimtime="00:10:14.12" />
                    <SPLIT distance="950" swimtime="00:10:48.84" />
                    <SPLIT distance="1000" swimtime="00:11:23.42" />
                    <SPLIT distance="1050" swimtime="00:11:58.02" />
                    <SPLIT distance="1100" swimtime="00:12:33.08" />
                    <SPLIT distance="1150" swimtime="00:13:07.58" />
                    <SPLIT distance="1200" swimtime="00:13:41.47" />
                    <SPLIT distance="1250" swimtime="00:14:15.31" />
                    <SPLIT distance="1300" swimtime="00:14:50.12" />
                    <SPLIT distance="1350" swimtime="00:15:24.55" />
                    <SPLIT distance="1400" swimtime="00:15:59.41" />
                    <SPLIT distance="1450" swimtime="00:16:32.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Jasiński" birthdate="2003-01-07" gender="M" nation="POL" license="101105700219" swrid="4947532" athleteid="2317">
              <RESULTS>
                <RESULT eventid="1120" points="529" reactiontime="+74" swimtime="00:00:25.85" resultid="2318" heatid="4031" lane="8" entrytime="00:00:26.61" entrycourse="LCM" />
                <RESULT eventid="1166" points="542" reactiontime="+83" swimtime="00:00:31.82" resultid="2319" heatid="4043" lane="2" entrytime="00:00:31.93" entrycourse="LCM" />
                <RESULT eventid="1396" points="535" reactiontime="+76" swimtime="00:00:27.43" resultid="2320" heatid="4093" lane="2" entrytime="00:00:27.76" entrycourse="LCM" />
                <RESULT eventid="1475" points="537" reactiontime="+83" swimtime="00:00:57.70" resultid="2321" heatid="4108" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gerard" lastname="Napieraj" birthdate="2009-12-23" gender="M" nation="POL" license="101105700282" swrid="4976720" athleteid="2352">
              <RESULTS>
                <RESULT eventid="1120" points="192" reactiontime="+90" swimtime="00:00:36.20" resultid="2353" heatid="4027" lane="9" entrytime="00:00:35.87" entrycourse="LCM" />
                <RESULT eventid="1258" points="176" reactiontime="+72" swimtime="00:00:42.79" resultid="2354" heatid="4057" lane="3" entrytime="00:00:44.71" entrycourse="LCM" />
                <RESULT eventid="1304" points="183" reactiontime="+77" swimtime="00:02:59.43" resultid="2355" heatid="4066" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:24.31" />
                    <SPLIT distance="150" swimtime="00:02:12.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="193" reactiontime="+88" swimtime="00:01:21.13" resultid="2356" heatid="4110" lane="9" entrytime="00:01:23.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="181" reactiontime="+62" swimtime="00:01:31.65" resultid="2357" heatid="4134" lane="8" entrytime="00:01:35.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="193" reactiontime="+60" swimtime="00:03:13.47" resultid="2358" heatid="4153" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="150" swimtime="00:02:26.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Kurzawa" birthdate="2007-03-28" gender="M" nation="POL" license="101105700237" swrid="5259892" athleteid="2363">
              <RESULTS>
                <RESULT eventid="1120" points="323" reactiontime="+76" swimtime="00:00:30.46" resultid="2364" heatid="4029" lane="7" entrytime="00:00:30.37" entrycourse="LCM" />
                <RESULT eventid="1258" points="248" reactiontime="+75" swimtime="00:00:38.17" resultid="2365" heatid="4058" lane="2" entrytime="00:00:37.95" entrycourse="LCM" />
                <RESULT eventid="1304" points="287" reactiontime="+86" swimtime="00:02:34.53" resultid="2366" heatid="4069" lane="3" entrytime="00:02:30.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:01:57.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="321" reactiontime="+81" swimtime="00:01:08.48" resultid="2367" heatid="4111" lane="2" entrytime="00:01:08.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Tkacz" birthdate="2009-11-16" gender="M" nation="POL" license="101105700254" swrid="4977282" athleteid="2393">
              <RESULTS>
                <RESULT eventid="1166" points="228" reactiontime="+82" swimtime="00:00:42.43" resultid="2394" heatid="4040" lane="7" entrytime="00:00:44.13" entrycourse="LCM" />
                <RESULT eventid="1350" points="189" reactiontime="+61" swimtime="00:01:39.10" resultid="2395" heatid="4078" lane="5" entrytime="00:01:41.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="197" reactiontime="+91" swimtime="00:03:36.71" resultid="2396" heatid="4120" lane="2" entrytime="00:03:36.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.81" />
                    <SPLIT distance="100" swimtime="00:01:43.97" />
                    <SPLIT distance="150" swimtime="00:02:41.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Liśkiewicz" birthdate="2008-04-05" gender="F" nation="POL" license="101105600290" swrid="5456466" athleteid="2306">
              <RESULTS>
                <RESULT eventid="1070" points="263" reactiontime="+85" swimtime="00:00:36.90" resultid="2307" heatid="4017" lane="9" entrytime="00:00:37.44" entrycourse="LCM" />
                <RESULT eventid="1327" points="232" reactiontime="+87" swimtime="00:01:44.33" resultid="2308" heatid="4074" lane="9" entrytime="00:01:47.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="240" swimtime="00:03:43.74" resultid="2309" heatid="4116" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.33" />
                    <SPLIT distance="100" swimtime="00:01:50.47" />
                    <SPLIT distance="150" swimtime="00:02:48.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="239" reactiontime="+93" swimtime="00:06:20.55" resultid="2310" heatid="4144" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                    <SPLIT distance="100" swimtime="00:01:29.00" />
                    <SPLIT distance="150" swimtime="00:02:18.26" />
                    <SPLIT distance="200" swimtime="00:03:07.30" />
                    <SPLIT distance="250" swimtime="00:03:56.55" />
                    <SPLIT distance="300" swimtime="00:04:46.45" />
                    <SPLIT distance="350" swimtime="00:05:34.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwier" lastname="Inglik" birthdate="2009-09-09" gender="M" nation="POL" license="101105700255" swrid="4977109" athleteid="2328">
              <RESULTS>
                <RESULT eventid="1120" points="186" reactiontime="+61" swimtime="00:00:36.60" resultid="2329" heatid="4025" lane="3" />
                <RESULT eventid="1166" points="155" reactiontime="+74" swimtime="00:00:48.21" resultid="2330" heatid="4039" lane="6" entrytime="00:00:51.19" entrycourse="LCM" />
                <RESULT eventid="1258" status="DNS" swimtime="00:00:00.00" resultid="2331" heatid="4056" lane="9" />
                <RESULT eventid="1350" points="144" reactiontime="+67" swimtime="00:01:48.32" resultid="2332" heatid="4078" lane="8" entrytime="00:01:50.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="180" reactiontime="+84" swimtime="00:01:22.93" resultid="2333" heatid="4109" lane="4" entrytime="00:01:23.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Jurda" birthdate="2009-02-04" gender="M" nation="POL" license="101105700259" swrid="5254078" athleteid="2386">
              <RESULTS>
                <RESULT eventid="1166" points="365" reactiontime="+72" swimtime="00:00:36.31" resultid="2387" heatid="4041" lane="4" entrytime="00:00:36.77" entrycourse="LCM" />
                <RESULT eventid="1258" points="281" reactiontime="+72" swimtime="00:00:36.63" resultid="2388" heatid="4058" lane="5" entrytime="00:00:36.99" entrycourse="LCM" />
                <RESULT eventid="1350" points="348" reactiontime="+73" swimtime="00:01:20.81" resultid="2389" heatid="4080" lane="9" entrytime="00:01:22.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="369" reactiontime="+83" swimtime="00:02:55.75" resultid="2390" heatid="4121" lane="6" entrytime="00:02:58.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:01:29.17" />
                    <SPLIT distance="150" swimtime="00:02:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="333" reactiontime="+88" swimtime="00:02:44.33" resultid="2391" heatid="4141" lane="3" entrytime="00:02:45.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:22.05" />
                    <SPLIT distance="150" swimtime="00:02:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="299" reactiontime="+82" swimtime="00:02:47.23" resultid="2392" heatid="4153" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:01:23.55" />
                    <SPLIT distance="150" swimtime="00:02:07.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Jasiński" birthdate="2003-01-07" gender="M" nation="POL" license="101105700218" swrid="4947533" athleteid="2409">
              <RESULTS>
                <RESULT eventid="1304" points="534" reactiontime="+70" swimtime="00:02:05.68" resultid="2410" heatid="4072" lane="7" entrytime="00:02:03.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                    <SPLIT distance="100" swimtime="00:01:01.61" />
                    <SPLIT distance="150" swimtime="00:01:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="558" reactiontime="+76" swimtime="00:09:08.88" resultid="2411" heatid="4097" lane="2" entrytime="00:09:16.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:04.89" />
                    <SPLIT distance="150" swimtime="00:01:39.33" />
                    <SPLIT distance="200" swimtime="00:02:13.73" />
                    <SPLIT distance="250" swimtime="00:02:48.28" />
                    <SPLIT distance="300" swimtime="00:03:22.51" />
                    <SPLIT distance="350" swimtime="00:03:56.88" />
                    <SPLIT distance="400" swimtime="00:04:31.27" />
                    <SPLIT distance="450" swimtime="00:05:05.74" />
                    <SPLIT distance="500" swimtime="00:05:40.58" />
                    <SPLIT distance="550" swimtime="00:06:15.42" />
                    <SPLIT distance="600" swimtime="00:06:50.25" />
                    <SPLIT distance="650" swimtime="00:07:25.42" />
                    <SPLIT distance="700" swimtime="00:08:00.60" />
                    <SPLIT distance="750" swimtime="00:08:35.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="522" reactiontime="+74" swimtime="00:00:58.26" resultid="2412" heatid="4107" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="587" reactiontime="+78" swimtime="00:04:22.81" resultid="2413" heatid="4149" lane="0" entrytime="00:04:33.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                    <SPLIT distance="100" swimtime="00:01:03.27" />
                    <SPLIT distance="150" swimtime="00:01:36.40" />
                    <SPLIT distance="200" swimtime="00:02:10.31" />
                    <SPLIT distance="250" swimtime="00:02:43.39" />
                    <SPLIT distance="300" swimtime="00:03:17.09" />
                    <SPLIT distance="350" swimtime="00:03:50.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Grzebieluch" birthdate="2005-07-29" gender="F" nation="POL" license="101105600265" swrid="5118445" athleteid="2296">
              <RESULTS>
                <RESULT eventid="1070" points="562" reactiontime="+69" swimtime="00:00:28.68" resultid="2297" heatid="4022" lane="9" entrytime="00:00:29.04" entrycourse="LCM" />
                <RESULT eventid="1235" points="624" reactiontime="+64" swimtime="00:00:31.56" resultid="2298" heatid="4055" lane="3" entrytime="00:00:31.73" entrycourse="LCM" />
                <RESULT eventid="1373" points="469" reactiontime="+74" swimtime="00:00:31.44" resultid="2299" heatid="4083" lane="0" />
                <RESULT eventid="1451" points="544" reactiontime="+69" swimtime="00:01:03.33" resultid="2300" heatid="4104" lane="6" entrytime="00:01:04.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="602" reactiontime="+66" swimtime="00:01:08.17" resultid="2301" heatid="4130" lane="3" entrytime="00:01:08.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="560" reactiontime="+67" swimtime="00:02:29.64" resultid="2302" heatid="4152" lane="3" entrytime="00:02:29.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:12.58" />
                    <SPLIT distance="150" swimtime="00:01:51.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Kruzerowska" birthdate="2004-09-20" gender="F" nation="POL" license="101105600107" swrid="4941663" athleteid="2290">
              <RESULTS>
                <RESULT eventid="1070" points="480" reactiontime="+85" swimtime="00:00:30.21" resultid="2291" heatid="4021" lane="0" entrytime="00:00:29.73" entrycourse="LCM" />
                <RESULT eventid="1235" points="577" reactiontime="+55" swimtime="00:00:32.40" resultid="2292" heatid="4055" lane="6" entrytime="00:00:32.56" entrycourse="LCM" />
                <RESULT eventid="1373" points="483" reactiontime="+73" swimtime="00:00:31.13" resultid="2293" heatid="4083" lane="2" />
                <RESULT eventid="1590" points="588" reactiontime="+51" swimtime="00:01:08.71" resultid="2294" heatid="4130" lane="5" entrytime="00:01:08.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="593" reactiontime="+55" swimtime="00:02:26.75" resultid="2295" heatid="4152" lane="4" entrytime="00:02:25.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:48.81" />
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kowalewski" birthdate="2006-08-15" gender="M" nation="POL" license="101105700170" swrid="5195497" athleteid="2283">
              <RESULTS>
                <RESULT eventid="1065" points="458" reactiontime="+77" swimtime="00:05:16.22" resultid="2284" heatid="4012" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:09.18" />
                    <SPLIT distance="150" swimtime="00:03:20.47" />
                    <SPLIT distance="200" swimtime="00:02:36.60" />
                    <SPLIT distance="250" swimtime="00:04:42.09" />
                    <SPLIT distance="300" swimtime="00:04:05.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="455" reactiontime="+79" swimtime="00:00:33.73" resultid="2285" heatid="4042" lane="5" entrytime="00:00:34.12" entrycourse="LCM" />
                <RESULT eventid="1350" points="408" reactiontime="+82" swimtime="00:01:16.69" resultid="2286" heatid="4080" lane="6" entrytime="00:01:17.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="473" reactiontime="+79" swimtime="00:02:41.78" resultid="2287" heatid="4122" lane="9" entrytime="00:02:45.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:19.60" />
                    <SPLIT distance="150" swimtime="00:02:01.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="344" reactiontime="+81" swimtime="00:02:38.03" resultid="2288" heatid="4124" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:12.63" />
                    <SPLIT distance="150" swimtime="00:01:55.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="405" reactiontime="+88" swimtime="00:02:34.08" resultid="2289" heatid="4140" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:01:58.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksy" lastname="Kusiński" birthdate="2002-06-04" gender="M" nation="POL" license="101105700248" swrid="4793534" athleteid="2322">
              <RESULTS>
                <RESULT eventid="1120" points="638" reactiontime="+74" swimtime="00:00:24.28" resultid="2323" heatid="4032" lane="5" entrytime="00:00:24.14" entrycourse="LCM" />
                <RESULT eventid="1258" points="602" reactiontime="+73" swimtime="00:00:28.41" resultid="2324" heatid="4060" lane="5" entrytime="00:00:28.47" entrycourse="LCM" />
                <RESULT eventid="1396" points="655" reactiontime="+75" swimtime="00:00:25.64" resultid="2325" heatid="4094" lane="4" entrytime="00:00:25.95" entrycourse="LCM" />
                <RESULT eventid="1475" points="670" reactiontime="+77" swimtime="00:00:53.60" resultid="2326" heatid="4115" lane="6" entrytime="00:00:52.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="593" reactiontime="+71" swimtime="00:01:01.69" resultid="2327" heatid="4132" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Czernielewski" birthdate="2008-12-30" gender="M" nation="POL" license="101105700233" swrid="4977036" athleteid="2311">
              <RESULTS>
                <RESULT eventid="1120" points="159" reactiontime="+87" swimtime="00:00:38.56" resultid="2312" heatid="4026" lane="6" entrytime="00:00:37.59" entrycourse="LCM" />
                <RESULT eventid="1258" points="140" reactiontime="+89" swimtime="00:00:46.21" resultid="2313" heatid="4057" lane="2" entrytime="00:00:45.27" entrycourse="LCM" />
                <RESULT eventid="1396" points="83" reactiontime="+75" swimtime="00:00:51.03" resultid="2314" heatid="4090" lane="3" />
                <RESULT eventid="1475" points="132" reactiontime="+98" swimtime="00:01:32.05" resultid="2315" heatid="4107" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="161" reactiontime="+87" swimtime="00:03:25.69" resultid="2316" heatid="4153" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                    <SPLIT distance="100" swimtime="00:01:45.20" />
                    <SPLIT distance="150" swimtime="00:02:37.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Szewczyk" birthdate="2004-12-21" gender="M" nation="POL" license="101105700110" swrid="5034854" athleteid="2405">
              <RESULTS>
                <RESULT eventid="1258" points="560" reactiontime="+67" swimtime="00:00:29.11" resultid="2406" heatid="4060" lane="3" entrytime="00:00:28.83" entrycourse="LCM" />
                <RESULT eventid="1396" points="554" reactiontime="+74" swimtime="00:00:27.10" resultid="2407" heatid="4094" lane="8" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="1613" points="581" reactiontime="+64" swimtime="00:01:02.11" resultid="2408" heatid="4136" lane="5" entrytime="00:01:02.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Kamiński" birthdate="2008-12-04" gender="M" nation="POL" license="101105700249" swrid="5334767" athleteid="2334">
              <RESULTS>
                <RESULT eventid="1120" points="333" reactiontime="+64" swimtime="00:00:30.16" resultid="2335" heatid="4028" lane="3" entrytime="00:00:31.36" entrycourse="LCM" />
                <RESULT eventid="1166" points="242" reactiontime="+64" swimtime="00:00:41.59" resultid="2336" heatid="4040" lane="5" entrytime="00:00:42.97" entrycourse="LCM" />
                <RESULT eventid="1350" points="224" swimtime="00:01:33.65" resultid="2337" heatid="4079" lane="9" entrytime="00:01:35.40" entrycourse="LCM" />
                <RESULT eventid="1396" points="250" reactiontime="+69" swimtime="00:00:35.33" resultid="2338" heatid="4090" lane="6" />
                <RESULT eventid="1475" points="301" reactiontime="+67" swimtime="00:01:09.94" resultid="2339" heatid="4106" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Pogoda" birthdate="2005-01-23" gender="M" nation="POL" license="101105700242" swrid="5113366" athleteid="2267">
              <RESULTS>
                <RESULT eventid="1065" points="604" reactiontime="+71" swimtime="00:04:48.40" resultid="2268" heatid="4013" lane="5" entrytime="00:04:44.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="150" swimtime="00:01:41.77" />
                    <SPLIT distance="200" swimtime="00:02:17.47" />
                    <SPLIT distance="250" swimtime="00:02:58.13" />
                    <SPLIT distance="300" swimtime="00:03:39.39" />
                    <SPLIT distance="350" swimtime="00:04:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="517" reactiontime="+68" swimtime="00:00:29.90" resultid="2269" heatid="4060" lane="1" entrytime="00:00:29.40" entrycourse="LCM" />
                <RESULT eventid="1350" points="533" reactiontime="+73" swimtime="00:01:10.14" resultid="2270" heatid="4077" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="572" reactiontime="+75" swimtime="00:02:31.91" resultid="2271" heatid="4120" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:12.76" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="550" reactiontime="+64" swimtime="00:01:03.27" resultid="2272" heatid="4136" lane="7" entrytime="00:01:03.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="578" reactiontime="+72" swimtime="00:02:16.83" resultid="2273" heatid="4142" lane="5" entrytime="00:02:14.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:04.73" />
                    <SPLIT distance="150" swimtime="00:01:45.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="584" reactiontime="+64" swimtime="00:02:13.86" resultid="2274" heatid="4155" lane="4" entrytime="00:02:09.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:05.91" />
                    <SPLIT distance="150" swimtime="00:01:40.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="583" reactiontime="+80" swimtime="00:17:22.42" resultid="2275" heatid="4159" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:05.17" />
                    <SPLIT distance="150" swimtime="00:01:39.44" />
                    <SPLIT distance="200" swimtime="00:02:13.81" />
                    <SPLIT distance="250" swimtime="00:02:48.08" />
                    <SPLIT distance="300" swimtime="00:03:22.70" />
                    <SPLIT distance="350" swimtime="00:03:57.40" />
                    <SPLIT distance="400" swimtime="00:04:32.23" />
                    <SPLIT distance="450" swimtime="00:05:07.08" />
                    <SPLIT distance="500" swimtime="00:05:41.96" />
                    <SPLIT distance="550" swimtime="00:06:17.02" />
                    <SPLIT distance="600" swimtime="00:06:52.03" />
                    <SPLIT distance="650" swimtime="00:07:27.02" />
                    <SPLIT distance="700" swimtime="00:08:02.13" />
                    <SPLIT distance="750" swimtime="00:08:37.26" />
                    <SPLIT distance="800" swimtime="00:09:12.08" />
                    <SPLIT distance="850" swimtime="00:09:47.20" />
                    <SPLIT distance="900" swimtime="00:10:22.33" />
                    <SPLIT distance="950" swimtime="00:10:57.39" />
                    <SPLIT distance="1000" swimtime="00:11:32.52" />
                    <SPLIT distance="1050" swimtime="00:12:07.92" />
                    <SPLIT distance="1100" swimtime="00:12:43.34" />
                    <SPLIT distance="1150" swimtime="00:13:18.70" />
                    <SPLIT distance="1200" swimtime="00:13:53.82" />
                    <SPLIT distance="1250" swimtime="00:14:28.93" />
                    <SPLIT distance="1300" swimtime="00:15:04.08" />
                    <SPLIT distance="1350" swimtime="00:15:39.26" />
                    <SPLIT distance="1400" swimtime="00:16:14.13" />
                    <SPLIT distance="1450" swimtime="00:16:48.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08614" nation="POL" region="14" clubid="3029" name="Stowarzyszenie SIG NOVUM">
          <ATHLETES>
            <ATHLETE firstname="Filip" lastname="Kusztykiewicz" birthdate="2008-11-19" gender="M" nation="POL" license="108614700023" swrid="5200061" athleteid="3051">
              <RESULTS>
                <RESULT eventid="1166" points="368" reactiontime="+73" swimtime="00:00:36.20" resultid="3052" heatid="4039" lane="8" />
                <RESULT eventid="1350" points="353" reactiontime="+70" swimtime="00:01:20.45" resultid="3053" heatid="4080" lane="7" entrytime="00:01:19.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Grzybowska" birthdate="2006-09-09" gender="F" nation="POL" license="108614600028" swrid="5166605" athleteid="3030">
              <RESULTS>
                <RESULT eventid="1070" points="466" reactiontime="+84" swimtime="00:00:30.53" resultid="3031" heatid="4015" lane="6" />
                <RESULT eventid="1235" points="381" reactiontime="+81" swimtime="00:00:37.20" resultid="3032" heatid="4052" lane="7" />
                <RESULT eventid="1281" points="416" reactiontime="+81" swimtime="00:02:31.28" resultid="3033" heatid="4061" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                    <SPLIT distance="150" swimtime="00:01:52.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Luterek" birthdate="2004-01-19" gender="F" nation="POL" license="108614600027" swrid="5200064" athleteid="3034">
              <RESULTS>
                <RESULT eventid="1070" points="452" reactiontime="+74" swimtime="00:00:30.82" resultid="3035" heatid="4015" lane="1" />
                <RESULT eventid="1143" points="443" reactiontime="+74" swimtime="00:00:38.56" resultid="3036" heatid="4034" lane="1" />
                <RESULT eventid="1373" points="338" reactiontime="+74" swimtime="00:00:35.04" resultid="3037" heatid="4084" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Żółtowski" birthdate="1975-03-22" gender="M" nation="POL" license="508614700063" swrid="4302693" athleteid="3041">
              <RESULTS>
                <RESULT eventid="1120" points="384" reactiontime="+80" swimtime="00:00:28.76" resultid="3042" heatid="4025" lane="1" />
                <RESULT eventid="1304" points="314" reactiontime="+81" swimtime="00:02:30.01" resultid="3043" heatid="4066" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:11.37" />
                    <SPLIT distance="150" swimtime="00:01:50.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Werpachowski" birthdate="2005-12-21" gender="M" nation="POL" license="108614700033" swrid="5108790" athleteid="3044">
              <RESULTS>
                <RESULT eventid="1120" points="529" reactiontime="+72" swimtime="00:00:25.84" resultid="3045" heatid="4024" lane="6" />
                <RESULT eventid="1212" points="514" reactiontime="+73" swimtime="00:01:01.76" resultid="3046" heatid="4047" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="473" reactiontime="+79" swimtime="00:02:10.86" resultid="3047" heatid="4068" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:04.07" />
                    <SPLIT distance="150" swimtime="00:01:38.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Woźniak" birthdate="2008-10-27" gender="F" nation="POL" license="108614600022" swrid="5200082" athleteid="3048">
              <RESULTS>
                <RESULT eventid="1143" points="334" swimtime="00:00:42.34" resultid="3049" heatid="4033" lane="5" />
                <RESULT eventid="1327" points="307" swimtime="00:01:35.02" resultid="3050" heatid="4074" lane="3" entrytime="00:01:34.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Szpak" birthdate="2006-09-29" gender="M" nation="POL" license="108614700047" swrid="5456638" athleteid="3038">
              <RESULTS>
                <RESULT eventid="1120" points="303" reactiontime="+76" swimtime="00:00:31.10" resultid="3039" heatid="4028" lane="2" entrytime="00:00:31.61" entrycourse="LCM" />
                <RESULT eventid="1396" points="262" reactiontime="+74" swimtime="00:00:34.78" resultid="3040" heatid="4090" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="07311" nation="POL" region="11" clubid="3100" name="UKS &quot;Dwójeczka&quot; Częstochowa">
          <ATHLETES>
            <ATHLETE firstname="Ireneusz" lastname="Stachurski" birthdate="1969-07-22" gender="M" nation="POL" license="107311700001" athleteid="3101">
              <RESULTS>
                <RESULT eventid="1475" points="190" swimtime="00:01:21.48" resultid="3102" heatid="4108" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="155" reactiontime="+48" swimtime="00:06:49.49" resultid="3103" heatid="4148" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:30.76" />
                    <SPLIT distance="150" swimtime="00:02:25.38" />
                    <SPLIT distance="200" swimtime="00:03:19.68" />
                    <SPLIT distance="250" swimtime="00:04:13.69" />
                    <SPLIT distance="300" swimtime="00:05:07.77" />
                    <SPLIT distance="350" swimtime="00:06:01.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01305" nation="POL" region="05" clubid="3478" name="UKS Piątka Konstantynów Łódzki">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Ber" birthdate="2007-04-19" gender="F" nation="POL" license="101305600220" swrid="5198056" athleteid="3518">
              <RESULTS>
                <RESULT eventid="1070" status="DNS" swimtime="00:00:00.00" resultid="3519" heatid="4020" lane="2" entrytime="00:00:30.06" entrycourse="LCM" />
                <RESULT eventid="1281" status="DNS" swimtime="00:00:00.00" resultid="3520" heatid="4065" lane="9" entrytime="00:02:19.58" entrycourse="LCM" />
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="3521" heatid="4104" lane="0" entrytime="00:01:04.84" entrycourse="LCM" />
                <RESULT eventid="1590" status="DNS" swimtime="00:00:00.00" resultid="3522" heatid="4127" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Figiel" birthdate="2007-05-18" gender="M" nation="POL" license="101305700224" swrid="5198058" athleteid="3557">
              <RESULTS>
                <RESULT eventid="1120" points="389" reactiontime="+64" swimtime="00:00:28.64" resultid="3558" heatid="4030" lane="6" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1304" points="430" reactiontime="+70" swimtime="00:02:15.10" resultid="3559" heatid="4071" lane="2" entrytime="00:02:11.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                    <SPLIT distance="100" swimtime="00:01:05.23" />
                    <SPLIT distance="150" swimtime="00:01:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="455" reactiontime="+66" swimtime="00:01:00.98" resultid="3560" heatid="4113" lane="6" entrytime="00:01:00.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1797" points="442" reactiontime="+69" swimtime="00:19:02.92" resultid="3561" heatid="4159" lane="1" entrytime="00:18:26.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:41.12" />
                    <SPLIT distance="200" swimtime="00:02:16.83" />
                    <SPLIT distance="250" swimtime="00:02:52.89" />
                    <SPLIT distance="300" swimtime="00:03:28.79" />
                    <SPLIT distance="350" swimtime="00:04:05.61" />
                    <SPLIT distance="400" swimtime="00:04:42.87" />
                    <SPLIT distance="450" swimtime="00:05:20.27" />
                    <SPLIT distance="500" swimtime="00:05:57.51" />
                    <SPLIT distance="550" swimtime="00:06:34.80" />
                    <SPLIT distance="600" swimtime="00:07:13.42" />
                    <SPLIT distance="650" swimtime="00:07:52.73" />
                    <SPLIT distance="700" swimtime="00:08:32.51" />
                    <SPLIT distance="750" swimtime="00:09:12.39" />
                    <SPLIT distance="800" swimtime="00:09:52.42" />
                    <SPLIT distance="850" swimtime="00:10:32.77" />
                    <SPLIT distance="900" swimtime="00:11:12.59" />
                    <SPLIT distance="950" swimtime="00:11:53.14" />
                    <SPLIT distance="1000" swimtime="00:12:33.24" />
                    <SPLIT distance="1050" swimtime="00:13:13.79" />
                    <SPLIT distance="1100" swimtime="00:13:53.47" />
                    <SPLIT distance="1150" swimtime="00:14:33.56" />
                    <SPLIT distance="1200" swimtime="00:15:13.79" />
                    <SPLIT distance="1250" swimtime="00:15:53.30" />
                    <SPLIT distance="1300" swimtime="00:16:32.53" />
                    <SPLIT distance="1350" swimtime="00:17:11.05" />
                    <SPLIT distance="1400" swimtime="00:17:49.06" />
                    <SPLIT distance="1450" swimtime="00:18:26.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Krata" birthdate="2009-07-22" gender="M" nation="POL" license="101305700289" swrid="5356912" athleteid="3552">
              <RESULTS>
                <RESULT eventid="1120" points="258" reactiontime="+83" swimtime="00:00:32.82" resultid="3553" heatid="4027" lane="1" entrytime="00:00:34.10" entrycourse="LCM" />
                <RESULT eventid="1304" points="194" reactiontime="+81" swimtime="00:02:55.96" resultid="3554" heatid="4068" lane="3" entrytime="00:03:46.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:24.78" />
                    <SPLIT distance="150" swimtime="00:02:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="228" reactiontime="+71" swimtime="00:01:16.71" resultid="3555" heatid="4107" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="162" reactiontime="+80" swimtime="00:01:34.94" resultid="3556" heatid="4133" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Nuszczyński" birthdate="2007-06-14" gender="M" nation="POL" license="101305700222" swrid="5198048" athleteid="3562">
              <RESULTS>
                <RESULT eventid="1120" points="360" reactiontime="+74" swimtime="00:00:29.39" resultid="3563" heatid="4029" lane="4" entrytime="00:00:29.36" entrycourse="LCM" />
                <RESULT eventid="1258" points="396" reactiontime="+74" swimtime="00:00:32.68" resultid="3564" heatid="4059" lane="2" entrytime="00:00:33.40" entrycourse="LCM" />
                <RESULT eventid="1304" points="339" reactiontime="+75" swimtime="00:02:26.20" resultid="3565" heatid="4067" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:47.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonina" lastname="Sulak" birthdate="2006-04-09" gender="F" nation="POL" license="101305600208" swrid="5075908" athleteid="3485">
              <RESULTS>
                <RESULT eventid="1060" points="595" reactiontime="+79" swimtime="00:05:16.54" resultid="3486" heatid="4011" lane="2" entrytime="00:05:18.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                    <SPLIT distance="150" swimtime="00:01:52.21" />
                    <SPLIT distance="200" swimtime="00:02:32.41" />
                    <SPLIT distance="250" swimtime="00:03:17.97" />
                    <SPLIT distance="300" swimtime="00:04:02.68" />
                    <SPLIT distance="350" swimtime="00:04:40.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="571" reactiontime="+75" swimtime="00:02:16.11" resultid="3487" heatid="4065" lane="2" entrytime="00:02:16.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                    <SPLIT distance="150" swimtime="00:01:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="550" reactiontime="+72" swimtime="00:01:03.11" resultid="3488" heatid="4105" lane="8" entrytime="00:01:03.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="553" reactiontime="+76" swimtime="00:02:33.65" resultid="3489" heatid="4138" lane="2" entrytime="00:02:31.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:12.87" />
                    <SPLIT distance="150" swimtime="00:01:58.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="544" reactiontime="+78" swimtime="00:09:53.75" resultid="3490" heatid="4156" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:10.79" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                    <SPLIT distance="200" swimtime="00:02:26.06" />
                    <SPLIT distance="250" swimtime="00:03:03.81" />
                    <SPLIT distance="300" swimtime="00:03:41.33" />
                    <SPLIT distance="350" swimtime="00:04:19.20" />
                    <SPLIT distance="400" swimtime="00:04:56.89" />
                    <SPLIT distance="450" swimtime="00:05:33.99" />
                    <SPLIT distance="500" swimtime="00:06:11.59" />
                    <SPLIT distance="550" swimtime="00:06:49.46" />
                    <SPLIT distance="600" swimtime="00:07:27.02" />
                    <SPLIT distance="650" swimtime="00:08:04.39" />
                    <SPLIT distance="700" swimtime="00:08:41.92" />
                    <SPLIT distance="750" swimtime="00:09:18.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Stankiewicz" birthdate="2005-07-26" gender="M" nation="POL" license="101305700173" swrid="5075901" athleteid="3582">
              <RESULTS>
                <RESULT comment="G1 - Pływak nie złamał powierzchni wody głową przed lub na linii 15 m po starcie lub nawrocie." eventid="1258" reactiontime="+62" status="DSQ" swimtime="00:00:31.78" resultid="3583" heatid="4059" lane="5" entrytime="00:00:31.36" entrycourse="LCM" />
                <RESULT eventid="1475" points="469" reactiontime="+66" swimtime="00:01:00.37" resultid="3584" heatid="4112" lane="3" entrytime="00:01:02.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="442" reactiontime="+66" swimtime="00:01:08.03" resultid="3585" heatid="4135" lane="5" entrytime="00:01:07.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="407" reactiontime="+70" swimtime="00:02:30.91" resultid="3586" heatid="4155" lane="0" entrytime="00:02:26.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:14.89" />
                    <SPLIT distance="150" swimtime="00:01:54.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Wawrzyniak" birthdate="2009-07-22" gender="F" nation="POL" license="101305600254" swrid="5288810" athleteid="3496">
              <RESULTS>
                <RESULT eventid="1070" points="328" reactiontime="+83" swimtime="00:00:34.31" resultid="3497" heatid="4017" lane="8" entrytime="00:00:36.78" entrycourse="LCM" />
                <RESULT eventid="1281" points="314" reactiontime="+91" swimtime="00:02:46.11" resultid="3498" heatid="4062" lane="3" entrytime="00:02:59.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:21.04" />
                    <SPLIT distance="150" swimtime="00:02:06.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="264" reactiontime="+88" swimtime="00:00:38.08" resultid="3499" heatid="4084" lane="3" entrytime="00:00:47.74" entrycourse="LCM" />
                <RESULT eventid="1451" points="342" reactiontime="+92" swimtime="00:01:13.92" resultid="3500" heatid="4100" lane="5" entrytime="00:01:22.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="240" swimtime="00:01:32.53" resultid="3501" heatid="4127" lane="5" entrytime="00:01:36.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karina" lastname="Łysakowska" birthdate="2006-03-22" gender="F" nation="POL" license="101305600215" swrid="5159128" athleteid="3513">
              <RESULTS>
                <RESULT eventid="1070" points="589" reactiontime="+76" swimtime="00:00:28.23" resultid="3514" heatid="4022" lane="5" entrytime="00:00:28.46" entrycourse="LCM" />
                <RESULT eventid="1373" points="550" reactiontime="+74" swimtime="00:00:29.80" resultid="3515" heatid="4088" lane="5" entrytime="00:00:29.75" entrycourse="LCM" />
                <RESULT eventid="1451" points="591" reactiontime="+77" swimtime="00:01:01.60" resultid="3516" heatid="4105" lane="4" entrytime="00:01:01.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="567" reactiontime="+78" swimtime="00:04:45.64" resultid="3517" heatid="4145" lane="3" entrytime="00:04:45.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                    <SPLIT distance="150" swimtime="00:01:43.32" />
                    <SPLIT distance="200" swimtime="00:02:19.96" />
                    <SPLIT distance="250" swimtime="00:02:56.40" />
                    <SPLIT distance="300" swimtime="00:03:33.33" />
                    <SPLIT distance="350" swimtime="00:04:10.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Sterniczuk" birthdate="2003-06-16" gender="F" nation="POL" license="101305600144" swrid="4947560" athleteid="3479">
              <RESULTS>
                <RESULT eventid="1060" points="523" reactiontime="+81" swimtime="00:05:30.54" resultid="3480" heatid="4011" lane="1" entrytime="00:05:32.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:57.91" />
                    <SPLIT distance="200" swimtime="00:02:40.75" />
                    <SPLIT distance="250" swimtime="00:03:27.17" />
                    <SPLIT distance="300" swimtime="00:04:14.37" />
                    <SPLIT distance="350" swimtime="00:04:52.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="458" reactiontime="+76" swimtime="00:00:38.12" resultid="3481" heatid="4037" lane="9" entrytime="00:00:38.36" entrycourse="LCM" />
                <RESULT eventid="1327" points="482" reactiontime="+76" swimtime="00:01:21.79" resultid="3482" heatid="4075" lane="5" entrytime="00:01:23.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="427" reactiontime="+79" swimtime="00:00:32.42" resultid="3483" heatid="4087" lane="3" entrytime="00:00:31.83" entrycourse="LCM" />
                <RESULT eventid="1498" points="476" reactiontime="+84" swimtime="00:02:58.15" resultid="3484" heatid="4118" lane="0" entrytime="00:02:58.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                    <SPLIT distance="150" swimtime="00:02:12.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Laudańska" birthdate="2009-09-21" gender="F" nation="POL" license="101305600279" swrid="4977075" athleteid="3502">
              <RESULTS>
                <RESULT eventid="1070" points="212" reactiontime="+84" swimtime="00:00:39.69" resultid="3503" heatid="4016" lane="6" entrytime="00:00:41.82" entrycourse="LCM" />
                <RESULT eventid="1327" points="127" reactiontime="+89" swimtime="00:02:07.42" resultid="3504" heatid="4073" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="186" reactiontime="+84" swimtime="00:01:30.47" resultid="3505" heatid="4100" lane="8" entrytime="00:01:37.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="161" reactiontime="+78" swimtime="00:01:45.68" resultid="3506" heatid="4127" lane="6" entrytime="00:01:48.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Kaczmarek" birthdate="2007-10-31" gender="F" nation="POL" license="101305600219" swrid="5198054" athleteid="3507">
              <RESULTS>
                <RESULT eventid="1070" points="534" reactiontime="+84" swimtime="00:00:29.16" resultid="3508" heatid="4022" lane="1" entrytime="00:00:28.86" entrycourse="LCM" />
                <RESULT eventid="1143" points="543" reactiontime="+81" swimtime="00:00:36.02" resultid="3509" heatid="4036" lane="3" entrytime="00:00:38.93" entrycourse="LCM" />
                <RESULT eventid="1327" points="524" reactiontime="+82" swimtime="00:01:19.50" resultid="3510" heatid="4075" lane="7" entrytime="00:01:27.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="502" reactiontime="+87" swimtime="00:01:05.03" resultid="3511" heatid="4105" lane="1" entrytime="00:01:03.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="516" reactiontime="+78" swimtime="00:02:37.18" resultid="3512" heatid="4138" lane="9" entrytime="00:02:38.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:02:00.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Kowalczyk" birthdate="2005-10-14" gender="F" nation="POL" license="101305600168" swrid="5075895" athleteid="3523">
              <RESULTS>
                <RESULT eventid="1070" points="466" reactiontime="+80" swimtime="00:00:30.51" resultid="3524" heatid="4020" lane="8" entrytime="00:00:30.78" entrycourse="LCM" />
                <RESULT eventid="1281" points="465" reactiontime="+85" swimtime="00:02:25.81" resultid="3525" heatid="4063" lane="3" entrytime="00:02:29.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:49.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="489" reactiontime="+90" swimtime="00:01:05.63" resultid="3526" heatid="4103" lane="3" entrytime="00:01:05.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="370" reactiontime="+82" swimtime="00:01:20.16" resultid="3527" heatid="4126" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Romanowski" birthdate="2003-06-16" gender="M" nation="POL" license="101305700141" swrid="4947551" athleteid="3544">
              <RESULTS>
                <RESULT eventid="1120" points="674" reactiontime="+66" swimtime="00:00:23.84" resultid="3545" heatid="4032" lane="4" entrytime="00:00:24.04" entrycourse="LCM" />
                <RESULT eventid="1396" points="608" reactiontime="+66" swimtime="00:00:26.28" resultid="3546" heatid="4094" lane="1" entrytime="00:00:26.37" entrycourse="LCM" />
                <RESULT eventid="1475" points="706" reactiontime="+65" swimtime="00:00:52.68" resultid="3547" heatid="4115" lane="4" entrytime="00:00:52.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Misztal" birthdate="2006-04-12" gender="M" nation="POL" license="101305700191" swrid="5138252" athleteid="3855">
              <RESULTS>
                <RESULT eventid="1120" points="456" reactiontime="+79" swimtime="00:00:27.16" resultid="3856" heatid="4031" lane="9" entrytime="00:00:26.96" entrycourse="LCM" />
                <RESULT eventid="1396" points="435" reactiontime="+80" swimtime="00:00:29.39" resultid="3857" heatid="4093" lane="9" entrytime="00:00:28.87" entrycourse="LCM" />
                <RESULT eventid="1166" points="374" reactiontime="+80" swimtime="00:00:36.01" resultid="3858" heatid="4042" lane="7" entrytime="00:00:35.76" entrycourse="LCM" />
                <RESULT eventid="1475" points="492" reactiontime="+80" swimtime="00:00:59.41" resultid="3859" heatid="4113" lane="7" entrytime="00:01:00.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="392" reactiontime="+77" swimtime="00:02:35.66" resultid="3860" heatid="4140" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:12.81" />
                    <SPLIT distance="150" swimtime="00:02:00.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Klaudia" lastname="Bujnowicz" birthdate="2007-09-26" gender="F" nation="POL" license="101305600223" swrid="5198051" athleteid="3533">
              <RESULTS>
                <RESULT eventid="1070" points="339" reactiontime="+83" swimtime="00:00:33.92" resultid="3534" heatid="4018" lane="0" entrytime="00:00:34.45" entrycourse="LCM" />
                <RESULT eventid="1235" points="295" reactiontime="+81" swimtime="00:00:40.50" resultid="3535" heatid="4053" lane="2" entrytime="00:00:39.96" entrycourse="LCM" />
                <RESULT eventid="1281" points="297" reactiontime="+81" swimtime="00:02:49.23" resultid="3536" heatid="4062" lane="4" entrytime="00:02:50.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:20.52" />
                    <SPLIT distance="150" swimtime="00:02:05.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="303" reactiontime="+80" swimtime="00:01:25.65" resultid="3537" heatid="4128" lane="2" entrytime="00:01:25.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="307" reactiontime="+86" swimtime="00:03:02.72" resultid="3538" heatid="4150" lane="4" entrytime="00:03:03.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:01:29.43" />
                    <SPLIT distance="150" swimtime="00:02:17.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Leśniewski" birthdate="2003-11-15" gender="M" nation="POL" license="101305700236" swrid="4947520" athleteid="3539">
              <RESULTS>
                <RESULT eventid="1120" points="521" reactiontime="+69" swimtime="00:00:25.97" resultid="3540" heatid="4031" lane="5" entrytime="00:00:25.80" entrycourse="LCM" />
                <RESULT eventid="1258" points="603" reactiontime="+65" swimtime="00:00:28.40" resultid="3541" heatid="4060" lane="6" entrytime="00:00:28.93" entrycourse="LCM" />
                <RESULT eventid="1475" points="531" reactiontime="+71" swimtime="00:00:57.90" resultid="3542" heatid="4114" lane="7" entrytime="00:00:56.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G1 - Pływak nie złamał powierzchni wody głową przed lub na linii 15 m po starcie lub nawrocie." eventid="1613" reactiontime="+65" status="DSQ" swimtime="00:01:07.18" resultid="3543" heatid="4135" lane="4" entrytime="00:01:06.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Skóra" birthdate="2003-08-05" gender="M" nation="POL" license="101305700143" swrid="5033406" athleteid="3577">
              <RESULTS>
                <RESULT eventid="1166" points="774" reactiontime="+72" swimtime="00:00:28.26" resultid="3578" heatid="4043" lane="4" entrytime="00:00:28.31" entrycourse="LCM" />
                <RESULT eventid="1350" points="700" reactiontime="+74" swimtime="00:01:04.06" resultid="3579" heatid="4081" lane="4" entrytime="00:01:02.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="612" reactiontime="+72" swimtime="00:00:26.22" resultid="3580" heatid="4089" lane="2" />
                <RESULT eventid="1521" points="638" reactiontime="+71" swimtime="00:02:26.50" resultid="3581" heatid="4122" lane="5" entrytime="00:02:24.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                    <SPLIT distance="150" swimtime="00:01:48.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Kowalczyk" birthdate="2009-04-27" gender="F" nation="POL" license="101305600272" swrid="5288817" athleteid="3491">
              <RESULTS>
                <RESULT eventid="1070" points="346" swimtime="00:00:33.69" resultid="3492" heatid="4015" lane="0" />
                <RESULT eventid="1189" points="246" reactiontime="+85" swimtime="00:01:28.52" resultid="3493" heatid="4044" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="275" reactiontime="+71" swimtime="00:00:37.53" resultid="3494" heatid="4084" lane="8" />
                <RESULT eventid="1451" points="305" swimtime="00:01:16.74" resultid="3495" heatid="4099" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Kaczanowska" birthdate="2005-03-14" gender="F" nation="POL" license="101305600321" swrid="5113368" athleteid="3528">
              <RESULTS>
                <RESULT eventid="1070" points="452" reactiontime="+74" swimtime="00:00:30.84" resultid="3529" heatid="4019" lane="4" entrytime="00:00:31.09" entrycourse="LCM" />
                <RESULT eventid="1281" points="442" reactiontime="+79" swimtime="00:02:28.28" resultid="3530" heatid="4063" lane="4" entrytime="00:02:27.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="150" swimtime="00:01:49.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="456" reactiontime="+78" swimtime="00:01:07.16" resultid="3531" heatid="4102" lane="4" entrytime="00:01:07.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="370" swimtime="00:01:20.14" resultid="3532" heatid="4129" lane="1" entrytime="00:01:19.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Pawlak" birthdate="2003-12-29" gender="M" nation="POL" license="101305700320" swrid="4947522" athleteid="3549">
              <RESULTS>
                <RESULT eventid="1120" points="521" reactiontime="+81" swimtime="00:00:25.97" resultid="3550" heatid="4031" lane="6" entrytime="00:00:26.15" entrycourse="LCM" />
                <RESULT eventid="1304" points="462" reactiontime="+87" swimtime="00:02:11.85" resultid="3551" heatid="4071" lane="1" entrytime="00:02:12.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="100" swimtime="00:01:03.70" />
                    <SPLIT distance="150" swimtime="00:01:38.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Rucińska" birthdate="2006-02-07" gender="F" nation="POL" license="101305600206" swrid="5075909" athleteid="3571">
              <RESULTS>
                <RESULT eventid="1143" points="499" reactiontime="+78" swimtime="00:00:37.05" resultid="3572" heatid="4036" lane="4" entrytime="00:00:38.42" entrycourse="LCM" />
                <RESULT eventid="1327" points="473" reactiontime="+82" swimtime="00:01:22.29" resultid="3573" heatid="4076" lane="0" entrytime="00:01:22.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="465" reactiontime="+68" swimtime="00:02:59.44" resultid="3574" heatid="4118" lane="7" entrytime="00:02:56.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="100" swimtime="00:01:26.29" />
                    <SPLIT distance="150" swimtime="00:02:13.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" status="DNS" swimtime="00:00:00.00" resultid="3575" heatid="4137" lane="6" entrytime="00:02:41.94" entrycourse="LCM" />
                <RESULT eventid="1728" points="423" reactiontime="+76" swimtime="00:02:44.23" resultid="3576" heatid="4152" lane="9" entrytime="00:02:38.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:21.47" />
                    <SPLIT distance="150" swimtime="00:02:03.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08114" nation="POL" region="14" clubid="2003" name="AZS  KU Uniwersytetu Warszawskiego">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Rębas" birthdate="1989-12-11" gender="M" nation="POL" license="508114700069" swrid="4251117" athleteid="2012">
              <RESULTS>
                <RESULT eventid="1212" points="572" reactiontime="+75" swimtime="00:00:59.63" resultid="2013" heatid="4047" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="550" reactiontime="+71" swimtime="00:00:27.18" resultid="2014" heatid="4090" lane="8" />
                <RESULT eventid="1475" status="DNS" swimtime="00:00:00.00" resultid="2015" heatid="4115" lane="9" entrytime="00:00:55.04" entrycourse="LCM" />
                <RESULT eventid="1659" status="DNS" swimtime="00:00:00.00" resultid="2016" heatid="4140" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Micorek" birthdate="1993-08-25" gender="M" nation="POL" license="108114700041" swrid="4086676" athleteid="2004">
              <RESULTS>
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="2005" heatid="4023" lane="4" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="2006" heatid="4047" lane="5" />
                <RESULT eventid="1396" points="557" reactiontime="+76" swimtime="00:00:27.06" resultid="2007" heatid="4094" lane="0" entrytime="00:00:27.25" entrycourse="LCM" />
                <RESULT eventid="1475" status="DNS" swimtime="00:00:00.00" resultid="2008" heatid="4106" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Godlewski" birthdate="1996-05-26" gender="M" nation="POL" license="108114700059" swrid="4285522" athleteid="2009">
              <RESULTS>
                <RESULT eventid="1166" points="551" reactiontime="+73" swimtime="00:00:31.65" resultid="2010" heatid="4043" lane="7" entrytime="00:00:32.18" entrycourse="LCM" />
                <RESULT eventid="1350" points="496" reactiontime="+80" swimtime="00:01:11.81" resultid="2011" heatid="4077" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03605" nation="POL" region="05" clubid="2177" name="KS ,,Masters&apos;&apos; Łódź">
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Adamska" birthdate="1984-09-25" gender="F" nation="POL" license="503605600036" athleteid="2188">
              <RESULTS>
                <RESULT eventid="1235" points="265" reactiontime="+72" swimtime="00:00:41.99" resultid="2189" heatid="4052" lane="9" />
                <RESULT eventid="1373" points="245" swimtime="00:00:39.03" resultid="2190" heatid="4084" lane="0" />
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="2191" heatid="4098" lane="8" />
                <RESULT eventid="1590" status="DNS" swimtime="00:00:00.00" resultid="2192" heatid="4127" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Olejarczyk" birthdate="1979-06-12" gender="M" nation="POL" license="503605700007" swrid="4992959" athleteid="2178">
              <RESULTS>
                <RESULT eventid="1120" points="481" reactiontime="+83" swimtime="00:00:26.67" resultid="2179" heatid="4024" lane="4" />
                <RESULT eventid="1212" points="425" reactiontime="+84" swimtime="00:01:05.82" resultid="2180" heatid="4048" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1475" points="455" reactiontime="+82" swimtime="00:01:00.97" resultid="2181" heatid="4107" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1567" points="287" reactiontime="+91" swimtime="00:02:47.86" resultid="2182" heatid="4124" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:59.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="503605600029" athleteid="2183">
              <RESULTS>
                <RESULT eventid="1189" points="114" reactiontime="+99" swimtime="00:01:54.17" resultid="2184" heatid="4044" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="130" reactiontime="+53" swimtime="00:03:42.46" resultid="2185" heatid="4061" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                    <SPLIT distance="100" swimtime="00:01:48.05" />
                    <SPLIT distance="150" swimtime="00:02:46.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="105" reactiontime="+88" swimtime="00:04:17.59" resultid="2186" heatid="4123" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.34" />
                    <SPLIT distance="100" swimtime="00:02:01.73" />
                    <SPLIT distance="150" swimtime="00:03:11.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="132" reactiontime="+90" swimtime="00:07:44.11" resultid="2187" heatid="4144" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.59" />
                    <SPLIT distance="100" swimtime="00:01:45.84" />
                    <SPLIT distance="150" swimtime="00:02:45.65" />
                    <SPLIT distance="200" swimtime="00:03:45.45" />
                    <SPLIT distance="250" swimtime="00:04:46.30" />
                    <SPLIT distance="300" swimtime="00:05:46.18" />
                    <SPLIT distance="350" swimtime="00:06:47.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08414" nation="POL" region="14" clubid="3689" name="UKS WAWER Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Maja" lastname="Wesołek" birthdate="2006-04-07" gender="F" nation="POL" license="108414600049" swrid="5462077" athleteid="3690">
              <RESULTS>
                <RESULT eventid="1070" status="DNS" swimtime="00:00:00.00" resultid="3691" heatid="4015" lane="5" />
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="3692" heatid="4051" lane="5" />
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="3693" heatid="4099" lane="3" />
                <RESULT eventid="1590" status="DNS" swimtime="00:00:00.00" resultid="3694" heatid="4126" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05415" nation="POL" region="15" clubid="2073" name="Kaliski Klub Sportowy  ,,Włókniarz&apos;&apos; 1925 Kalisz">
          <ATHLETES>
            <ATHLETE firstname="Miłosz" lastname="Żurawski" birthdate="2007-11-10" gender="M" nation="POL" license="105415700154" swrid="4998230" athleteid="2106">
              <RESULTS>
                <RESULT eventid="1521" points="304" reactiontime="+75" swimtime="00:03:07.48" resultid="2107" heatid="4121" lane="9" entrytime="00:03:08.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                    <SPLIT distance="100" swimtime="00:01:32.59" />
                    <SPLIT distance="150" swimtime="00:02:22.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="299" reactiontime="+72" swimtime="00:05:29.00" resultid="2108" heatid="4148" lane="7" entrytime="00:05:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:19.00" />
                    <SPLIT distance="150" swimtime="00:02:00.97" />
                    <SPLIT distance="200" swimtime="00:02:42.88" />
                    <SPLIT distance="250" swimtime="00:03:25.22" />
                    <SPLIT distance="300" swimtime="00:04:07.15" />
                    <SPLIT distance="350" swimtime="00:04:50.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Tyc" birthdate="2005-02-11" gender="M" nation="POL" license="105415700234" swrid="5202216" athleteid="2096">
              <RESULTS>
                <RESULT eventid="1475" points="259" reactiontime="+83" swimtime="00:01:13.57" resultid="2097" heatid="4108" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="258" reactiontime="+92" swimtime="00:03:17.98" resultid="2098" heatid="4119" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="100" swimtime="00:01:38.78" />
                    <SPLIT distance="150" swimtime="00:02:29.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Szymański" birthdate="2005-05-06" gender="M" nation="POL" license="105415700007" swrid="4945641" athleteid="2086">
              <RESULTS>
                <RESULT eventid="1475" points="532" reactiontime="+67" swimtime="00:00:57.86" resultid="2087" heatid="4106" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="537" reactiontime="+66" swimtime="00:01:03.78" resultid="2088" heatid="4136" lane="2" entrytime="00:01:03.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="534" reactiontime="+64" swimtime="00:02:17.93" resultid="2089" heatid="4155" lane="7" entrytime="00:02:17.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="150" swimtime="00:01:43.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Krupka" birthdate="2007-08-25" gender="F" nation="POL" license="105415600130" swrid="4901159" athleteid="2082">
              <RESULTS>
                <RESULT eventid="1451" points="424" reactiontime="+73" swimtime="00:01:08.81" resultid="2083" heatid="4102" lane="7" entrytime="00:01:09.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="339" reactiontime="+60" swimtime="00:01:22.50" resultid="2084" heatid="4127" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1682" points="313" reactiontime="+73" swimtime="00:05:48.03" resultid="2085" heatid="4144" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:18.82" />
                    <SPLIT distance="150" swimtime="00:02:03.40" />
                    <SPLIT distance="200" swimtime="00:02:49.23" />
                    <SPLIT distance="250" swimtime="00:03:34.89" />
                    <SPLIT distance="300" swimtime="00:04:21.08" />
                    <SPLIT distance="350" swimtime="00:05:05.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kacprzyk" birthdate="2005-03-28" gender="M" nation="POL" license="105415700233" swrid="5164754" athleteid="2099">
              <RESULTS>
                <RESULT eventid="1475" points="341" reactiontime="+73" swimtime="00:01:07.09" resultid="2100" heatid="4112" lane="9" entrytime="00:01:07.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="173" reactiontime="+77" swimtime="00:01:32.95" resultid="2101" heatid="4133" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Jarzycka" birthdate="2006-01-19" gender="F" nation="POL" license="105415600153" swrid="5153513" athleteid="2074">
              <RESULTS>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="2075" heatid="4102" lane="2" entrytime="00:01:08.99" entrycourse="LCM" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2076" heatid="4116" lane="1" />
                <RESULT eventid="1682" status="DNS" swimtime="00:00:00.00" resultid="2077" heatid="4143" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Stodzież" birthdate="2007-02-09" gender="M" nation="POL" license="105415700149" swrid="4997813" athleteid="2102">
              <RESULTS>
                <RESULT eventid="1521" points="272" reactiontime="+83" swimtime="00:03:14.63" resultid="2103" heatid="4119" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                    <SPLIT distance="100" swimtime="00:01:35.63" />
                    <SPLIT distance="150" swimtime="00:02:27.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="341" reactiontime="+73" swimtime="00:01:14.17" resultid="2104" heatid="4135" lane="6" entrytime="00:01:11.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="329" reactiontime="+82" swimtime="00:02:42.12" resultid="2105" heatid="4154" lane="2" entrytime="00:02:42.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:21.70" />
                    <SPLIT distance="150" swimtime="00:02:03.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Harabasz" birthdate="2007-07-01" gender="M" nation="POL" license="105415700066" swrid="5197753" athleteid="2093">
              <RESULTS>
                <RESULT eventid="1475" points="317" reactiontime="+80" swimtime="00:01:08.79" resultid="2094" heatid="4108" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="303" reactiontime="+78" swimtime="00:05:27.54" resultid="2095" heatid="4147" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:59.18" />
                    <SPLIT distance="200" swimtime="00:02:41.44" />
                    <SPLIT distance="250" swimtime="00:03:24.22" />
                    <SPLIT distance="300" swimtime="00:04:07.63" />
                    <SPLIT distance="350" swimtime="00:04:50.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Spychalski" birthdate="2007-01-07" gender="M" nation="POL" license="105415700161" swrid="5249561" athleteid="2090">
              <RESULTS>
                <RESULT eventid="1475" points="268" reactiontime="+88" swimtime="00:01:12.72" resultid="2091" heatid="4110" lane="5" entrytime="00:01:12.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="222" reactiontime="+89" swimtime="00:01:25.59" resultid="2092" heatid="4132" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Juszczak" birthdate="2007-03-28" gender="F" nation="POL" license="105415600046" swrid="5197762" athleteid="2078">
              <RESULTS>
                <RESULT eventid="1451" points="301" reactiontime="+80" swimtime="00:01:17.15" resultid="2079" heatid="4098" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="342" reactiontime="+77" swimtime="00:01:22.27" resultid="2080" heatid="4129" lane="9" entrytime="00:01:20.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="315" reactiontime="+65" swimtime="00:03:01.10" resultid="2081" heatid="4151" lane="8" entrytime="00:02:56.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                    <SPLIT distance="100" swimtime="00:01:28.58" />
                    <SPLIT distance="150" swimtime="00:02:15.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03015" nation="POL" region="15" clubid="3299" name="UKS Fala Swarzędz">
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Wermiński" birthdate="2004-09-26" gender="M" nation="POL" license="103015700016" swrid="5096951" athleteid="3304">
              <RESULTS>
                <RESULT eventid="1120" points="550" reactiontime="+70" swimtime="00:00:25.51" resultid="3305" heatid="4023" lane="3" />
                <RESULT eventid="1258" points="481" reactiontime="+89" swimtime="00:00:30.63" resultid="3306" heatid="4056" lane="8" />
                <RESULT eventid="1350" points="540" reactiontime="+68" swimtime="00:01:09.84" resultid="3307" heatid="4081" lane="6" entrytime="00:01:08.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Szmyt" birthdate="2003-04-16" gender="M" nation="POL" license="103015700022" swrid="4920334" athleteid="3300">
              <RESULTS>
                <RESULT eventid="1120" points="576" reactiontime="+78" swimtime="00:00:25.12" resultid="3301" heatid="4024" lane="1" />
                <RESULT comment="G1 - Pływak nie złamał powierzchni wody głową przed lub na linii 15 m po starcie lub nawrocie." eventid="1258" reactiontime="+71" status="DSQ" swimtime="00:00:28.50" resultid="3302" heatid="4060" lane="4" entrytime="00:00:28.43" entrycourse="LCM" />
                <RESULT eventid="1396" points="550" reactiontime="+71" swimtime="00:00:27.18" resultid="3303" heatid="4089" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00805" nation="POL" region="05" clubid="2872" name="Sekcja Pływacka Meduza Pajęczno">
          <ATHLETES>
            <ATHLETE firstname="Mikołaj" lastname="Popiel" birthdate="2006-01-01" gender="M" nation="POL" license="100805700087" swrid="5191084" athleteid="2873">
              <RESULTS>
                <RESULT eventid="1613" points="603" reactiontime="+67" swimtime="00:01:01.37" resultid="2874" heatid="4136" lane="6" entrytime="00:01:02.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1751" points="593" reactiontime="+62" swimtime="00:02:13.19" resultid="2875" heatid="4155" lane="5" entrytime="00:02:12.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:05.89" />
                    <SPLIT distance="150" swimtime="00:01:40.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02105" nation="POL" region="05" clubid="2216" name="LKS ,,Opocznianka&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Filip" lastname="Bielecki" birthdate="2008-12-17" gender="M" nation="POL" license="102105700035" swrid="5356910" athleteid="2245">
              <RESULTS>
                <RESULT eventid="1120" points="196" reactiontime="+83" swimtime="00:00:35.95" resultid="2246" heatid="4027" lane="8" entrytime="00:00:34.97" entrycourse="LCM" />
                <RESULT eventid="1258" points="130" reactiontime="+81" swimtime="00:00:47.29" resultid="2247" heatid="4057" lane="7" entrytime="00:00:45.34" entrycourse="LCM" />
                <RESULT eventid="1475" points="213" swimtime="00:01:18.47" resultid="2248" heatid="4108" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="141" reactiontime="+91" swimtime="00:01:39.43" resultid="2249" heatid="4133" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Bogusławska" birthdate="2008-01-03" gender="F" nation="POL" license="102105600020" swrid="5213997" athleteid="2233">
              <RESULTS>
                <RESULT eventid="1070" points="373" reactiontime="+67" swimtime="00:00:32.86" resultid="2234" heatid="4018" lane="5" entrytime="00:00:33.48" entrycourse="LCM" />
                <RESULT eventid="1327" points="320" reactiontime="+57" swimtime="00:01:33.69" resultid="2235" heatid="4074" lane="7" entrytime="00:01:35.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Bogatek" birthdate="2008-06-03" gender="F" nation="POL" license="102105600010" swrid="5203912" athleteid="2217">
              <RESULTS>
                <RESULT eventid="1070" points="440" reactiontime="+69" swimtime="00:00:31.12" resultid="2218" heatid="4019" lane="3" entrytime="00:00:31.25" entrycourse="LCM" />
                <RESULT eventid="1373" points="287" reactiontime="+72" swimtime="00:00:37.00" resultid="2219" heatid="4086" lane="1" entrytime="00:00:35.36" entrycourse="LCM" />
                <RESULT eventid="1451" points="417" reactiontime="+68" swimtime="00:01:09.17" resultid="2220" heatid="4102" lane="3" entrytime="00:01:07.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="343" reactiontime="+83" swimtime="00:01:22.17" resultid="2221" heatid="4126" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Pęczek" birthdate="2007-08-27" gender="M" nation="POL" license="102105700026" swrid="4951738" athleteid="2250">
              <RESULTS>
                <RESULT eventid="1120" points="336" reactiontime="+89" swimtime="00:00:30.07" resultid="2251" heatid="4029" lane="1" entrytime="00:00:30.66" entrycourse="LCM" />
                <RESULT eventid="1258" points="262" reactiontime="+79" swimtime="00:00:37.46" resultid="2252" heatid="4056" lane="2" />
                <RESULT eventid="1475" points="336" swimtime="00:01:07.41" resultid="2253" heatid="4107" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="300" reactiontime="+73" swimtime="00:01:17.37" resultid="2254" heatid="4135" lane="8" entrytime="00:01:18.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Melka" birthdate="2009-06-30" gender="F" nation="POL" license="102105600030" swrid="5214052" athleteid="2222">
              <RESULTS>
                <RESULT eventid="1070" points="384" reactiontime="+79" swimtime="00:00:32.55" resultid="2223" heatid="4018" lane="4" entrytime="00:00:33.27" entrycourse="LCM" />
                <RESULT eventid="1143" points="317" reactiontime="+74" swimtime="00:00:43.09" resultid="2224" heatid="4034" lane="8" />
                <RESULT eventid="1373" points="271" swimtime="00:00:37.73" resultid="2225" heatid="4085" lane="3" entrytime="00:00:37.13" entrycourse="LCM" />
                <RESULT eventid="1451" points="354" reactiontime="+75" swimtime="00:01:13.03" resultid="2226" heatid="4099" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="324" reactiontime="+81" swimtime="00:01:23.81" resultid="2227" heatid="4128" lane="0" entrytime="00:01:30.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Bogatek" birthdate="2007-04-11" gender="M" nation="POL" license="102105700011" swrid="4951550" athleteid="2239">
              <RESULTS>
                <RESULT eventid="1120" points="422" reactiontime="+67" swimtime="00:00:27.86" resultid="2240" heatid="4030" lane="7" entrytime="00:00:28.20" entrycourse="LCM" />
                <RESULT eventid="1258" points="401" reactiontime="+77" swimtime="00:00:32.52" resultid="2241" heatid="4059" lane="1" entrytime="00:00:35.04" entrycourse="LCM" />
                <RESULT eventid="1475" points="455" reactiontime="+66" swimtime="00:01:00.97" resultid="2242" heatid="4112" lane="4" entrytime="00:01:01.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="409" reactiontime="+79" swimtime="00:01:09.80" resultid="2243" heatid="4135" lane="3" entrytime="00:01:10.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="387" reactiontime="+68" swimtime="00:05:01.77" resultid="2244" heatid="4147" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                    <SPLIT distance="150" swimtime="00:01:53.46" />
                    <SPLIT distance="200" swimtime="00:02:31.36" />
                    <SPLIT distance="250" swimtime="00:03:10.23" />
                    <SPLIT distance="300" swimtime="00:03:49.37" />
                    <SPLIT distance="350" swimtime="00:04:26.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kalina" lastname="Kęska" birthdate="2008-05-16" gender="F" nation="POL" license="102105600021" swrid="5214053" athleteid="2236">
              <RESULTS>
                <RESULT eventid="1070" points="321" reactiontime="+95" swimtime="00:00:34.55" resultid="2237" heatid="4018" lane="8" entrytime="00:00:34.31" entrycourse="LCM" />
                <RESULT eventid="1327" points="267" reactiontime="+87" swimtime="00:01:39.58" resultid="2238" heatid="4074" lane="2" entrytime="00:01:35.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Stańczyk" birthdate="2009-12-05" gender="F" nation="POL" license="102105600029" swrid="5225174" athleteid="2228">
              <RESULTS>
                <RESULT eventid="1070" points="217" swimtime="00:00:39.33" resultid="2229" heatid="4016" lane="3" entrytime="00:00:39.45" entrycourse="LCM" />
                <RESULT eventid="1235" points="177" reactiontime="+74" swimtime="00:00:48.01" resultid="2230" heatid="4052" lane="5" entrytime="00:00:45.45" entrycourse="LCM" />
                <RESULT eventid="1451" points="204" reactiontime="+72" swimtime="00:01:27.83" resultid="2231" heatid="4100" lane="1" entrytime="00:01:27.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="181" reactiontime="+85" swimtime="00:01:41.72" resultid="2232" heatid="4127" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Faustyna" lastname="Karbownik" birthdate="2008-01-01" gender="F" nation="POL" license="102105600023" swrid="5203932" athleteid="2255">
              <RESULTS>
                <RESULT eventid="1189" points="164" reactiontime="+90" swimtime="00:01:41.20" resultid="2256" heatid="4045" lane="9" entrytime="00:01:24.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="161" reactiontime="+85" swimtime="00:00:44.85" resultid="2257" heatid="4083" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04005" nation="POL" region="05" clubid="2115" name="KP Raw-Swim">
          <ATHLETES>
            <ATHLETE firstname="Oliwia" lastname="Kłos" birthdate="2007-02-03" gender="F" nation="POL" license="104005600001" swrid="5198067" athleteid="2121">
              <RESULTS>
                <RESULT eventid="1070" points="526" reactiontime="+73" swimtime="00:00:29.31" resultid="2122" heatid="4021" lane="4" entrytime="00:00:29.33" entrycourse="LCM" />
                <RESULT eventid="1143" points="505" reactiontime="+81" swimtime="00:00:36.90" resultid="2123" heatid="4037" lane="1" entrytime="00:00:36.55" entrycourse="LCM" />
                <RESULT eventid="1451" points="450" reactiontime="+82" swimtime="00:01:07.46" resultid="2124" heatid="4098" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1774" points="356" reactiontime="+79" swimtime="00:11:23.80" resultid="2125" heatid="4156" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:01:58.17" />
                    <SPLIT distance="200" swimtime="00:02:41.12" />
                    <SPLIT distance="250" swimtime="00:03:24.62" />
                    <SPLIT distance="300" swimtime="00:04:08.05" />
                    <SPLIT distance="350" swimtime="00:04:52.67" />
                    <SPLIT distance="400" swimtime="00:05:36.33" />
                    <SPLIT distance="450" swimtime="00:06:20.86" />
                    <SPLIT distance="500" swimtime="00:07:04.70" />
                    <SPLIT distance="550" swimtime="00:07:48.90" />
                    <SPLIT distance="600" swimtime="00:08:32.90" />
                    <SPLIT distance="650" swimtime="00:09:16.88" />
                    <SPLIT distance="700" swimtime="00:09:59.98" />
                    <SPLIT distance="750" swimtime="00:10:43.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Majewski" birthdate="2008-06-02" gender="M" nation="POL" license="104005700004" swrid="5096067" athleteid="2138">
              <RESULTS>
                <RESULT eventid="1120" points="264" reactiontime="+68" swimtime="00:00:32.58" resultid="2139" heatid="4028" lane="6" entrytime="00:00:31.59" entrycourse="LCM" />
                <RESULT eventid="1166" points="300" reactiontime="+79" swimtime="00:00:38.74" resultid="2140" heatid="4041" lane="0" entrytime="00:00:40.99" entrycourse="LCM" />
                <RESULT eventid="1396" points="236" reactiontime="+70" swimtime="00:00:35.99" resultid="2141" heatid="4091" lane="3" entrytime="00:00:36.72" entrycourse="LCM" />
                <RESULT eventid="1475" points="273" reactiontime="+72" swimtime="00:01:12.31" resultid="2142" heatid="4110" lane="2" entrytime="00:01:12.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1521" points="258" reactiontime="+71" swimtime="00:03:18.03" resultid="2143" heatid="4119" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                    <SPLIT distance="100" swimtime="00:01:35.54" />
                    <SPLIT distance="150" swimtime="00:02:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1659" points="260" reactiontime="+70" swimtime="00:02:58.51" resultid="2144" heatid="4140" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:25.90" />
                    <SPLIT distance="150" swimtime="00:02:17.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Galińska" birthdate="2008-10-21" gender="F" nation="POL" license="104005600006" swrid="5096186" athleteid="2132">
              <RESULTS>
                <RESULT eventid="1070" points="372" reactiontime="+82" swimtime="00:00:32.90" resultid="2133" heatid="4019" lane="8" entrytime="00:00:32.29" entrycourse="LCM" />
                <RESULT eventid="1235" points="344" reactiontime="+76" swimtime="00:00:38.49" resultid="2134" heatid="4053" lane="3" entrytime="00:00:38.68" entrycourse="LCM" />
                <RESULT eventid="1373" points="289" reactiontime="+79" swimtime="00:00:36.95" resultid="2135" heatid="4082" lane="5" />
                <RESULT eventid="1451" points="354" reactiontime="+80" swimtime="00:01:13.07" resultid="2136" heatid="4102" lane="8" entrytime="00:01:11.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="320" reactiontime="+82" swimtime="00:01:24.16" resultid="2137" heatid="4128" lane="6" entrytime="00:01:24.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julita" lastname="Niewczas" birthdate="2008-05-15" gender="F" nation="POL" license="104005600008" swrid="5198068" athleteid="2116">
              <RESULTS>
                <RESULT eventid="1070" points="529" reactiontime="+83" swimtime="00:00:29.25" resultid="2117" heatid="4021" lane="2" entrytime="00:00:29.51" entrycourse="LCM" />
                <RESULT eventid="1327" points="489" reactiontime="+91" swimtime="00:01:21.37" resultid="2118" heatid="4076" lane="1" entrytime="00:01:20.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="516" reactiontime="+80" swimtime="00:01:04.46" resultid="2119" heatid="4103" lane="5" entrytime="00:01:05.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1728" points="431" reactiontime="+84" swimtime="00:02:43.21" resultid="2120" heatid="4150" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                    <SPLIT distance="150" swimtime="00:02:04.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roxana" lastname="Mydłowska" birthdate="2010-07-29" gender="F" nation="POL" license="104005600024" swrid="5277455" athleteid="3699">
              <RESULTS>
                <RESULT eventid="1070" points="350" reactiontime="+72" status="EXH" swimtime="00:00:33.57" resultid="3700" heatid="4015" lane="7" />
                <RESULT eventid="1451" points="342" reactiontime="+60" status="EXH" swimtime="00:01:13.89" resultid="3701" heatid="4101" lane="3" entrytime="00:01:13.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="315" reactiontime="+78" status="EXH" swimtime="00:02:46.01" resultid="3702" heatid="4061" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:04.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Szcześniak" birthdate="2009-07-10" gender="F" nation="POL" license="104005600015" swrid="5254099" athleteid="2126">
              <RESULTS>
                <RESULT eventid="1070" points="439" reactiontime="+87" swimtime="00:00:31.13" resultid="2127" heatid="4019" lane="0" entrytime="00:00:32.59" entrycourse="LCM" />
                <RESULT eventid="1143" points="310" reactiontime="+68" swimtime="00:00:43.40" resultid="2128" heatid="4035" lane="7" entrytime="00:00:43.87" entrycourse="LCM" />
                <RESULT eventid="1327" points="302" reactiontime="+86" swimtime="00:01:35.57" resultid="2129" heatid="4074" lane="1" entrytime="00:01:35.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="330" reactiontime="+76" swimtime="00:00:35.32" resultid="2130" heatid="4085" lane="5" entrytime="00:00:36.91" entrycourse="LCM" />
                <RESULT eventid="1451" points="398" reactiontime="+79" swimtime="00:01:10.25" resultid="2131" heatid="4101" lane="4" entrytime="00:01:12.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kumanowski" birthdate="2008-10-20" gender="M" nation="POL" license="104005700005" swrid="5096065" athleteid="2151">
              <RESULTS>
                <RESULT eventid="1120" points="406" reactiontime="+77" swimtime="00:00:28.22" resultid="2152" heatid="4030" lane="8" entrytime="00:00:28.40" entrycourse="LCM" />
                <RESULT eventid="1212" points="351" reactiontime="+72" swimtime="00:01:10.16" resultid="2153" heatid="4049" lane="9" entrytime="00:01:10.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="388" reactiontime="+79" swimtime="00:00:30.51" resultid="2154" heatid="4092" lane="8" entrytime="00:00:32.13" entrycourse="LCM" />
                <RESULT eventid="1475" points="387" reactiontime="+75" swimtime="00:01:04.33" resultid="2155" heatid="4112" lane="6" entrytime="00:01:03.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Szubert-Olszacki" birthdate="2009-01-13" gender="M" nation="POL" license="104005700014" swrid="5269103" athleteid="2145">
              <RESULTS>
                <RESULT eventid="1120" points="308" reactiontime="+72" swimtime="00:00:30.93" resultid="2146" heatid="4028" lane="5" entrytime="00:00:31.26" entrycourse="LCM" />
                <RESULT eventid="1166" points="238" reactiontime="+78" swimtime="00:00:41.87" resultid="2147" heatid="4040" lane="6" entrytime="00:00:43.12" entrycourse="LCM" />
                <RESULT eventid="1396" points="211" reactiontime="+76" swimtime="00:00:37.37" resultid="2148" heatid="4091" lane="8" entrytime="00:00:37.85" entrycourse="LCM" />
                <RESULT eventid="1475" points="304" reactiontime="+64" swimtime="00:01:09.76" resultid="2149" heatid="4111" lane="7" entrytime="00:01:08.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1705" points="312" reactiontime="+69" swimtime="00:05:24.30" resultid="2150" heatid="4147" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:16.87" />
                    <SPLIT distance="150" swimtime="00:01:58.26" />
                    <SPLIT distance="200" swimtime="00:02:39.11" />
                    <SPLIT distance="250" swimtime="00:03:21.14" />
                    <SPLIT distance="300" swimtime="00:04:04.00" />
                    <SPLIT distance="350" swimtime="00:04:45.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00405" nation="POL" region="05" clubid="2049" name="EKS Skra Bełchatów">
          <ATHLETES>
            <ATHLETE firstname="Maja" lastname="Górny" birthdate="2007-06-28" gender="F" nation="POL" license="100405600129" swrid="5196295" athleteid="2050">
              <RESULTS>
                <RESULT eventid="1070" points="456" reactiontime="+81" swimtime="00:00:30.73" resultid="2051" heatid="4020" lane="1" entrytime="00:00:30.48" entrycourse="LCM" />
                <RESULT eventid="1281" points="434" reactiontime="+80" swimtime="00:02:29.13" resultid="2052" heatid="4063" lane="6" entrytime="00:02:30.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:12.27" />
                    <SPLIT distance="150" swimtime="00:01:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="299" reactiontime="+87" swimtime="00:00:36.50" resultid="2053" heatid="4086" lane="0" entrytime="00:00:35.74" entrycourse="LCM" />
                <RESULT eventid="1451" points="468" reactiontime="+76" swimtime="00:01:06.58" resultid="2054" heatid="4103" lane="9" entrytime="00:01:06.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="355" reactiontime="+67" swimtime="00:01:21.28" resultid="2055" heatid="4129" lane="8" entrytime="00:01:19.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Sokołowska" birthdate="2007-03-18" gender="F" nation="POL" license="100405600136" swrid="5219474" athleteid="2056">
              <RESULTS>
                <RESULT eventid="1070" points="410" reactiontime="+88" swimtime="00:00:31.85" resultid="2057" heatid="4019" lane="1" entrytime="00:00:32.06" entrycourse="LCM" />
                <RESULT eventid="1189" points="297" reactiontime="+77" swimtime="00:01:23.09" resultid="2058" heatid="4045" lane="8" entrytime="00:01:21.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="313" reactiontime="+87" swimtime="00:00:35.98" resultid="2059" heatid="4086" lane="8" entrytime="00:00:35.58" entrycourse="LCM" />
                <RESULT eventid="1451" points="389" reactiontime="+87" swimtime="00:01:10.81" resultid="2060" heatid="4102" lane="1" entrytime="00:01:09.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1636" points="368" reactiontime="+86" swimtime="00:02:55.95" resultid="2061" heatid="4137" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:24.24" />
                    <SPLIT distance="150" swimtime="00:02:16.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Kowalczyk" birthdate="2007-03-11" gender="M" nation="POL" license="100405700146" swrid="5400118" athleteid="2062">
              <RESULTS>
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="2063" heatid="4027" lane="5" entrytime="00:00:32.74" entrycourse="LCM" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="2064" heatid="4069" lane="6" entrytime="00:02:33.18" entrycourse="LCM" />
                <RESULT eventid="1475" status="DNS" swimtime="00:00:00.00" resultid="2065" heatid="4107" lane="4" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="2066" heatid="4132" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

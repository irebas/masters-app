<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="MTP Delfin Cieszyn" version="Build 23880">
    <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Katowice" name="Zimowe Otwarte Mistrzostwa Polski Masters" course="SCM" hostclub="UKS Wodnik 29 Katowice" hostclub.url="http://www.wodnik29.pl" nation="POL" organizer="UKS Wodnik 29 Katowice" organizer.url="http://www.wodnik29.pl" timing="AUTOMATIC">
      <AGEDATE value="2014-11-16" type="YEAR" />
      <POOL name="AZS AWF KATOWICE" lanemin="1" lanemax="6" />
      <POINTTABLE pointtableid="3005" name="FINA Point Scoring" version="2012" />
      <CONTACT city="Katowice" email="kontakt@delfincieszyn.pl" name="Łukasz Widzik" phone="660749175" street="Mikołowska 72" />
      <SESSIONS>
        <SESSION date="2014-11-14" daytime="11:00" name="I Blok (Piątek)" number="1" warmupfrom="10:00">
          <EVENTS>
            <EVENT eventid="1058" daytime="11:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1060" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2661" />
                    <RANKING order="2" place="2" resultid="7253" />
                    <RANKING order="3" place="3" resultid="7215" />
                    <RANKING order="4" place="4" resultid="6457" />
                    <RANKING order="5" place="5" resultid="7189" />
                    <RANKING order="6" place="6" resultid="5074" />
                    <RANKING order="7" place="7" resultid="6181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1061" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7134" />
                    <RANKING order="2" place="2" resultid="5812" />
                    <RANKING order="3" place="3" resultid="2361" />
                    <RANKING order="4" place="4" resultid="4216" />
                    <RANKING order="5" place="5" resultid="5969" />
                    <RANKING order="6" place="6" resultid="6383" />
                    <RANKING order="7" place="7" resultid="2781" />
                    <RANKING order="8" place="8" resultid="4985" />
                    <RANKING order="9" place="-1" resultid="3251" />
                    <RANKING order="10" place="-1" resultid="3927" />
                    <RANKING order="11" place="-1" resultid="5585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3148" />
                    <RANKING order="2" place="2" resultid="4111" />
                    <RANKING order="3" place="3" resultid="4719" />
                    <RANKING order="4" place="4" resultid="5527" />
                    <RANKING order="5" place="5" resultid="6376" />
                    <RANKING order="6" place="6" resultid="6371" />
                    <RANKING order="7" place="7" resultid="6036" />
                    <RANKING order="8" place="-1" resultid="5834" />
                    <RANKING order="9" place="-1" resultid="6360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3716" />
                    <RANKING order="2" place="2" resultid="6052" />
                    <RANKING order="3" place="3" resultid="3732" />
                    <RANKING order="4" place="4" resultid="4264" />
                    <RANKING order="5" place="5" resultid="3908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5746" />
                    <RANKING order="2" place="2" resultid="5502" />
                    <RANKING order="3" place="3" resultid="4411" />
                    <RANKING order="4" place="4" resultid="5125" />
                    <RANKING order="5" place="5" resultid="6206" />
                    <RANKING order="6" place="6" resultid="4426" />
                    <RANKING order="7" place="7" resultid="6365" />
                    <RANKING order="8" place="8" resultid="5579" />
                    <RANKING order="9" place="9" resultid="5604" />
                    <RANKING order="10" place="10" resultid="5801" />
                    <RANKING order="11" place="11" resultid="5707" />
                    <RANKING order="12" place="-1" resultid="5390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4395" />
                    <RANKING order="2" place="2" resultid="3469" />
                    <RANKING order="3" place="3" resultid="2828" />
                    <RANKING order="4" place="4" resultid="4848" />
                    <RANKING order="5" place="5" resultid="3808" />
                    <RANKING order="6" place="-1" resultid="6379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5483" />
                    <RANKING order="2" place="2" resultid="5434" />
                    <RANKING order="3" place="3" resultid="6201" />
                    <RANKING order="4" place="4" resultid="6196" />
                    <RANKING order="5" place="5" resultid="5662" />
                    <RANKING order="6" place="6" resultid="5596" />
                    <RANKING order="7" place="7" resultid="6083" />
                    <RANKING order="8" place="-1" resultid="5343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6186" />
                    <RANKING order="2" place="2" resultid="4893" />
                    <RANKING order="3" place="3" resultid="4540" />
                    <RANKING order="4" place="4" resultid="2837" />
                    <RANKING order="5" place="5" resultid="4462" />
                    <RANKING order="6" place="6" resultid="3670" />
                    <RANKING order="7" place="7" resultid="6076" />
                    <RANKING order="8" place="-1" resultid="5322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4901" />
                    <RANKING order="2" place="2" resultid="4744" />
                    <RANKING order="3" place="3" resultid="3538" />
                    <RANKING order="4" place="4" resultid="3572" />
                    <RANKING order="5" place="-1" resultid="3403" />
                    <RANKING order="6" place="-1" resultid="3560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6097" />
                    <RANKING order="2" place="2" resultid="5346" />
                    <RANKING order="3" place="3" resultid="4702" />
                    <RANKING order="4" place="4" resultid="5058" />
                    <RANKING order="5" place="5" resultid="4489" />
                    <RANKING order="6" place="6" resultid="3553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4726" />
                    <RANKING order="2" place="2" resultid="3566" />
                    <RANKING order="3" place="3" resultid="2472" />
                    <RANKING order="4" place="4" resultid="3547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1073" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1059" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1074" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7331" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7332" daytime="11:01" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7333" daytime="11:03" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7334" daytime="11:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7335" daytime="11:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7336" daytime="11:07" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7337" daytime="11:08" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7338" daytime="11:09" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7339" daytime="11:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7340" daytime="11:11" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7341" daytime="11:12" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7342" daytime="11:13" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7343" daytime="11:14" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7344" daytime="11:15" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" daytime="11:17" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1076" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2479" />
                    <RANKING order="2" place="2" resultid="2503" />
                    <RANKING order="3" place="3" resultid="7206" />
                    <RANKING order="4" place="4" resultid="2599" />
                    <RANKING order="5" place="5" resultid="6476" />
                    <RANKING order="6" place="6" resultid="3429" />
                    <RANKING order="7" place="7" resultid="7226" />
                    <RANKING order="8" place="8" resultid="6354" />
                    <RANKING order="9" place="9" resultid="4003" />
                    <RANKING order="10" place="10" resultid="4134" />
                    <RANKING order="11" place="-1" resultid="7197" />
                    <RANKING order="12" place="-1" resultid="2455" />
                    <RANKING order="13" place="-1" resultid="6484" />
                    <RANKING order="14" place="-1" resultid="7150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7222" />
                    <RANKING order="2" place="2" resultid="5788" />
                    <RANKING order="3" place="3" resultid="5104" />
                    <RANKING order="4" place="4" resultid="4456" />
                    <RANKING order="5" place="5" resultid="3441" />
                    <RANKING order="6" place="6" resultid="2761" />
                    <RANKING order="7" place="7" resultid="2788" />
                    <RANKING order="8" place="8" resultid="2736" />
                    <RANKING order="9" place="9" resultid="2747" />
                    <RANKING order="10" place="10" resultid="5118" />
                    <RANKING order="11" place="11" resultid="5179" />
                    <RANKING order="12" place="12" resultid="3229" />
                    <RANKING order="13" place="13" resultid="2973" />
                    <RANKING order="14" place="-1" resultid="2752" />
                    <RANKING order="15" place="-1" resultid="4223" />
                    <RANKING order="16" place="-1" resultid="4379" />
                    <RANKING order="17" place="-1" resultid="5184" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2962" />
                    <RANKING order="2" place="2" resultid="4121" />
                    <RANKING order="3" place="3" resultid="2796" />
                    <RANKING order="4" place="4" resultid="6451" />
                    <RANKING order="5" place="5" resultid="2722" />
                    <RANKING order="6" place="6" resultid="6464" />
                    <RANKING order="7" place="7" resultid="3876" />
                    <RANKING order="8" place="8" resultid="2562" />
                    <RANKING order="9" place="9" resultid="2952" />
                    <RANKING order="10" place="10" resultid="3955" />
                    <RANKING order="11" place="11" resultid="2901" />
                    <RANKING order="12" place="12" resultid="6318" />
                    <RANKING order="13" place="13" resultid="6332" />
                    <RANKING order="14" place="14" resultid="2906" />
                    <RANKING order="15" place="15" resultid="3443" />
                    <RANKING order="16" place="16" resultid="5026" />
                    <RANKING order="17" place="17" resultid="5860" />
                    <RANKING order="18" place="18" resultid="4140" />
                    <RANKING order="19" place="19" resultid="3246" />
                    <RANKING order="20" place="20" resultid="2741" />
                    <RANKING order="21" place="21" resultid="2977" />
                    <RANKING order="22" place="21" resultid="3241" />
                    <RANKING order="23" place="23" resultid="2943" />
                    <RANKING order="24" place="24" resultid="2896" />
                    <RANKING order="25" place="25" resultid="2887" />
                    <RANKING order="26" place="26" resultid="2968" />
                    <RANKING order="27" place="27" resultid="2756" />
                    <RANKING order="28" place="28" resultid="6327" />
                    <RANKING order="29" place="29" resultid="4971" />
                    <RANKING order="30" place="30" resultid="4753" />
                    <RANKING order="31" place="-1" resultid="4317" />
                    <RANKING order="32" place="-1" resultid="5197" />
                    <RANKING order="33" place="-1" resultid="5898" />
                    <RANKING order="34" place="-1" resultid="5907" />
                    <RANKING order="35" place="-1" resultid="5945" />
                    <RANKING order="36" place="-1" resultid="6061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5978" />
                    <RANKING order="2" place="2" resultid="6311" />
                    <RANKING order="3" place="3" resultid="5474" />
                    <RANKING order="4" place="4" resultid="4785" />
                    <RANKING order="5" place="5" resultid="2912" />
                    <RANKING order="6" place="6" resultid="6292" />
                    <RANKING order="7" place="7" resultid="6300" />
                    <RANKING order="8" place="8" resultid="5515" />
                    <RANKING order="9" place="9" resultid="4938" />
                    <RANKING order="10" place="10" resultid="5866" />
                    <RANKING order="11" place="11" resultid="4092" />
                    <RANKING order="12" place="12" resultid="7127" />
                    <RANKING order="13" place="13" resultid="2929" />
                    <RANKING order="14" place="14" resultid="2981" />
                    <RANKING order="15" place="15" resultid="2883" />
                    <RANKING order="16" place="16" resultid="3748" />
                    <RANKING order="17" place="17" resultid="2918" />
                    <RANKING order="18" place="18" resultid="4671" />
                    <RANKING order="19" place="19" resultid="6029" />
                    <RANKING order="20" place="20" resultid="6322" />
                    <RANKING order="21" place="-1" resultid="3775" />
                    <RANKING order="22" place="-1" resultid="5952" />
                    <RANKING order="23" place="-1" resultid="6149" />
                    <RANKING order="24" place="-1" resultid="6420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5369" />
                    <RANKING order="2" place="2" resultid="4794" />
                    <RANKING order="3" place="3" resultid="4293" />
                    <RANKING order="4" place="4" resultid="3235" />
                    <RANKING order="5" place="5" resultid="5571" />
                    <RANKING order="6" place="6" resultid="3760" />
                    <RANKING order="7" place="7" resultid="3157" />
                    <RANKING order="8" place="8" resultid="3740" />
                    <RANKING order="9" place="9" resultid="5609" />
                    <RANKING order="10" place="10" resultid="3177" />
                    <RANKING order="11" place="11" resultid="4311" />
                    <RANKING order="12" place="12" resultid="5590" />
                    <RANKING order="13" place="13" resultid="4821" />
                    <RANKING order="14" place="14" resultid="3768" />
                    <RANKING order="15" place="15" resultid="3224" />
                    <RANKING order="16" place="16" resultid="3172" />
                    <RANKING order="17" place="17" resultid="5820" />
                    <RANKING order="18" place="18" resultid="4338" />
                    <RANKING order="19" place="19" resultid="3692" />
                    <RANKING order="20" place="20" resultid="5767" />
                    <RANKING order="21" place="21" resultid="3695" />
                    <RANKING order="22" place="22" resultid="6351" />
                    <RANKING order="23" place="-1" resultid="2807" />
                    <RANKING order="24" place="-1" resultid="3445" />
                    <RANKING order="25" place="-1" resultid="3686" />
                    <RANKING order="26" place="-1" resultid="3754" />
                    <RANKING order="27" place="-1" resultid="4065" />
                    <RANKING order="28" place="-1" resultid="6469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3039" />
                    <RANKING order="2" place="2" resultid="5132" />
                    <RANKING order="3" place="3" resultid="3489" />
                    <RANKING order="4" place="4" resultid="2646" />
                    <RANKING order="5" place="5" resultid="2488" />
                    <RANKING order="6" place="6" resultid="3260" />
                    <RANKING order="7" place="7" resultid="6258" />
                    <RANKING order="8" place="8" resultid="4857" />
                    <RANKING order="9" place="9" resultid="4075" />
                    <RANKING order="10" place="10" resultid="5760" />
                    <RANKING order="11" place="11" resultid="4635" />
                    <RANKING order="12" place="12" resultid="3635" />
                    <RANKING order="13" place="13" resultid="4803" />
                    <RANKING order="14" place="14" resultid="4102" />
                    <RANKING order="15" place="15" resultid="4044" />
                    <RANKING order="16" place="16" resultid="5652" />
                    <RANKING order="17" place="17" resultid="6252" />
                    <RANKING order="18" place="18" resultid="3885" />
                    <RANKING order="19" place="19" resultid="4344" />
                    <RANKING order="20" place="20" resultid="3189" />
                    <RANKING order="21" place="21" resultid="4546" />
                    <RANKING order="22" place="22" resultid="4554" />
                    <RANKING order="23" place="-1" resultid="3934" />
                    <RANKING order="24" place="-1" resultid="2414" />
                    <RANKING order="25" place="-1" resultid="3047" />
                    <RANKING order="26" place="-1" resultid="3216" />
                    <RANKING order="27" place="-1" resultid="4964" />
                    <RANKING order="28" place="-1" resultid="5332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6432" />
                    <RANKING order="2" place="2" resultid="4620" />
                    <RANKING order="3" place="3" resultid="2532" />
                    <RANKING order="4" place="4" resultid="2593" />
                    <RANKING order="5" place="5" resultid="3056" />
                    <RANKING order="6" place="6" resultid="6246" />
                    <RANKING order="7" place="7" resultid="4505" />
                    <RANKING order="8" place="8" resultid="3805" />
                    <RANKING order="9" place="9" resultid="4830" />
                    <RANKING order="10" place="10" resultid="3679" />
                    <RANKING order="11" place="11" resultid="6239" />
                    <RANKING order="12" place="12" resultid="2435" />
                    <RANKING order="13" place="13" resultid="5522" />
                    <RANKING order="14" place="14" resultid="2572" />
                    <RANKING order="15" place="-1" resultid="4151" />
                    <RANKING order="16" place="-1" resultid="5304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4302" />
                    <RANKING order="2" place="2" resultid="2445" />
                    <RANKING order="3" place="3" resultid="5772" />
                    <RANKING order="4" place="4" resultid="5336" />
                    <RANKING order="5" place="5" resultid="4647" />
                    <RANKING order="6" place="6" resultid="4748" />
                    <RANKING order="7" place="7" resultid="6068" />
                    <RANKING order="8" place="8" resultid="6443" />
                    <RANKING order="9" place="9" resultid="6220" />
                    <RANKING order="10" place="10" resultid="2844" />
                    <RANKING order="11" place="11" resultid="3941" />
                    <RANKING order="12" place="12" resultid="4689" />
                    <RANKING order="13" place="13" resultid="2551" />
                    <RANKING order="14" place="14" resultid="5450" />
                    <RANKING order="15" place="15" resultid="5252" />
                    <RANKING order="16" place="16" resultid="6225" />
                    <RANKING order="17" place="-1" resultid="3132" />
                    <RANKING order="18" place="-1" resultid="4449" />
                    <RANKING order="19" place="-1" resultid="5533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2466" />
                    <RANKING order="2" place="2" resultid="2391" />
                    <RANKING order="3" place="3" resultid="5936" />
                    <RANKING order="4" place="4" resultid="5752" />
                    <RANKING order="5" place="5" resultid="3394" />
                    <RANKING order="6" place="6" resultid="3368" />
                    <RANKING order="7" place="-1" resultid="7236" />
                    <RANKING order="8" place="-1" resultid="2426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2404" />
                    <RANKING order="2" place="2" resultid="4740" />
                    <RANKING order="3" place="3" resultid="4812" />
                    <RANKING order="4" place="4" resultid="5491" />
                    <RANKING order="5" place="5" resultid="4480" />
                    <RANKING order="6" place="6" resultid="5464" />
                    <RANKING order="7" place="7" resultid="2853" />
                    <RANKING order="8" place="8" resultid="4760" />
                    <RANKING order="9" place="9" resultid="4444" />
                    <RANKING order="10" place="10" resultid="3592" />
                    <RANKING order="11" place="-1" resultid="4207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4914" />
                    <RANKING order="2" place="2" resultid="6131" />
                    <RANKING order="3" place="3" resultid="4526" />
                    <RANKING order="4" place="4" resultid="4566" />
                    <RANKING order="5" place="5" resultid="3611" />
                    <RANKING order="6" place="6" resultid="3584" />
                    <RANKING order="7" place="7" resultid="4023" />
                    <RANKING order="8" place="8" resultid="3624" />
                    <RANKING order="9" place="9" resultid="3628" />
                    <RANKING order="10" place="-1" resultid="5005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4638" />
                    <RANKING order="2" place="2" resultid="2382" />
                    <RANKING order="3" place="3" resultid="5794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3867" />
                    <RANKING order="2" place="2" resultid="4402" />
                    <RANKING order="3" place="-1" resultid="5327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1090" agemax="94" agemin="90" name="N: 90 - 94 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7345" daytime="11:17" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7346" daytime="11:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7347" daytime="11:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7348" daytime="11:27" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7349" daytime="11:29" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7350" daytime="11:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7351" daytime="11:31" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7352" daytime="11:32" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7353" daytime="11:33" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7354" daytime="11:34" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7355" daytime="11:35" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7356" daytime="11:37" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7357" daytime="11:38" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7358" daytime="11:39" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7359" daytime="11:40" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7360" daytime="11:41" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7361" daytime="11:42" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7362" daytime="11:43" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7363" daytime="11:44" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7364" daytime="11:45" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="7365" daytime="11:46" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="7366" daytime="11:47" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="7367" daytime="11:48" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="7368" daytime="11:49" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="7369" daytime="11:50" number="25" order="25" status="OFFICIAL" />
                <HEAT heatid="7370" daytime="11:51" number="26" order="26" status="OFFICIAL" />
                <HEAT heatid="7371" daytime="11:52" number="27" order="27" status="OFFICIAL" />
                <HEAT heatid="7372" daytime="11:53" number="28" order="28" status="OFFICIAL" />
                <HEAT heatid="7373" daytime="11:54" number="29" order="29" status="OFFICIAL" />
                <HEAT heatid="7374" daytime="11:54" number="30" order="30" status="OFFICIAL" />
                <HEAT heatid="7375" daytime="11:55" number="31" order="31" status="OFFICIAL" />
                <HEAT heatid="7376" daytime="11:56" number="32" order="32" status="OFFICIAL" />
                <HEAT heatid="7377" daytime="11:57" number="33" order="33" status="OFFICIAL" />
                <HEAT heatid="7378" daytime="11:58" number="34" order="34" status="OFFICIAL" />
                <HEAT heatid="7379" daytime="11:59" number="35" order="35" status="OFFICIAL" />
                <HEAT heatid="7380" daytime="12:00" number="36" order="36" status="OFFICIAL" />
                <HEAT heatid="7381" daytime="12:01" number="37" order="37" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="12:02" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2662" />
                    <RANKING order="2" place="2" resultid="5173" />
                    <RANKING order="3" place="3" resultid="3519" />
                    <RANKING order="4" place="-1" resultid="5851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4498" />
                    <RANKING order="2" place="2" resultid="5970" />
                    <RANKING order="3" place="3" resultid="4256" />
                    <RANKING order="4" place="4" resultid="2715" />
                    <RANKING order="5" place="5" resultid="2705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3149" />
                    <RANKING order="2" place="2" resultid="4112" />
                    <RANKING order="3" place="3" resultid="6037" />
                    <RANKING order="4" place="-1" resultid="6140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5509" />
                    <RANKING order="2" place="2" resultid="5503" />
                    <RANKING order="3" place="3" resultid="3526" />
                    <RANKING order="4" place="4" resultid="6366" />
                    <RANKING order="5" place="5" resultid="7244" />
                    <RANKING order="6" place="6" resultid="5580" />
                    <RANKING order="7" place="7" resultid="2671" />
                    <RANKING order="8" place="-1" resultid="3723" />
                    <RANKING order="9" place="-1" resultid="4712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4534" />
                    <RANKING order="2" place="2" resultid="2829" />
                    <RANKING order="3" place="3" resultid="4275" />
                    <RANKING order="4" place="4" resultid="4849" />
                    <RANKING order="5" place="5" resultid="6044" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4908" />
                    <RANKING order="2" place="2" resultid="5484" />
                    <RANKING order="3" place="3" resultid="6090" />
                    <RANKING order="4" place="4" resultid="4471" />
                    <RANKING order="5" place="5" resultid="6084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4680" />
                    <RANKING order="2" place="2" resultid="4894" />
                    <RANKING order="3" place="3" resultid="4463" />
                    <RANKING order="4" place="4" resultid="3671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3404" />
                    <RANKING order="2" place="2" resultid="4438" />
                    <RANKING order="3" place="3" resultid="3386" />
                    <RANKING order="4" place="4" resultid="3978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6022" />
                    <RANKING order="2" place="2" resultid="4490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1104" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1105" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1106" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1107" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1108" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7382" daytime="12:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7383" daytime="12:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7384" daytime="12:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7385" daytime="12:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7386" daytime="12:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7387" daytime="12:27" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7388" daytime="12:31" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7389" daytime="12:35" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="12:38" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7198" />
                    <RANKING order="2" place="2" resultid="2600" />
                    <RANKING order="3" place="3" resultid="2504" />
                    <RANKING order="4" place="4" resultid="6338" />
                    <RANKING order="5" place="5" resultid="7227" />
                    <RANKING order="6" place="-1" resultid="6477" />
                    <RANKING order="7" place="-1" resultid="6485" />
                    <RANKING order="8" place="-1" resultid="7151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7142" />
                    <RANKING order="2" place="2" resultid="5105" />
                    <RANKING order="3" place="3" resultid="5166" />
                    <RANKING order="4" place="4" resultid="2762" />
                    <RANKING order="5" place="5" resultid="4417" />
                    <RANKING order="6" place="-1" resultid="4222" />
                    <RANKING order="7" place="-1" resultid="4380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4626" />
                    <RANKING order="2" place="2" resultid="3996" />
                    <RANKING order="3" place="3" resultid="2723" />
                    <RANKING order="4" place="4" resultid="2585" />
                    <RANKING order="5" place="5" resultid="2542" />
                    <RANKING order="6" place="6" resultid="4325" />
                    <RANKING order="7" place="7" resultid="3877" />
                    <RANKING order="8" place="8" resultid="2953" />
                    <RANKING order="9" place="9" resultid="6346" />
                    <RANKING order="10" place="10" resultid="2888" />
                    <RANKING order="11" place="11" resultid="2944" />
                    <RANKING order="12" place="-1" resultid="2936" />
                    <RANKING order="13" place="-1" resultid="5899" />
                    <RANKING order="14" place="-1" resultid="5908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5979" />
                    <RANKING order="2" place="2" resultid="3206" />
                    <RANKING order="3" place="3" resultid="4786" />
                    <RANKING order="4" place="4" resultid="5475" />
                    <RANKING order="5" place="5" resultid="5141" />
                    <RANKING order="6" place="6" resultid="6150" />
                    <RANKING order="7" place="7" resultid="3988" />
                    <RANKING order="8" place="8" resultid="4839" />
                    <RANKING order="9" place="9" resultid="5313" />
                    <RANKING order="10" place="10" resultid="5825" />
                    <RANKING order="11" place="-1" resultid="5953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4795" />
                    <RANKING order="2" place="2" resultid="4294" />
                    <RANKING order="3" place="3" resultid="4605" />
                    <RANKING order="4" place="4" resultid="5572" />
                    <RANKING order="5" place="5" resultid="3741" />
                    <RANKING order="6" place="6" resultid="4822" />
                    <RANKING order="7" place="-1" resultid="2808" />
                    <RANKING order="8" place="-1" resultid="3900" />
                    <RANKING order="9" place="-1" resultid="4066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3490" />
                    <RANKING order="2" place="2" resultid="3040" />
                    <RANKING order="3" place="3" resultid="5133" />
                    <RANKING order="4" place="4" resultid="2489" />
                    <RANKING order="5" place="5" resultid="2372" />
                    <RANKING order="6" place="6" resultid="2655" />
                    <RANKING order="7" place="7" resultid="3935" />
                    <RANKING order="8" place="8" resultid="4930" />
                    <RANKING order="9" place="9" resultid="3800" />
                    <RANKING order="10" place="10" resultid="4858" />
                    <RANKING order="11" place="11" resultid="5653" />
                    <RANKING order="12" place="12" resultid="5381" />
                    <RANKING order="13" place="13" resultid="4675" />
                    <RANKING order="14" place="-1" resultid="3217" />
                    <RANKING order="15" place="-1" resultid="3636" />
                    <RANKING order="16" place="-1" resultid="4965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6017" />
                    <RANKING order="2" place="2" resultid="2533" />
                    <RANKING order="3" place="3" resultid="4831" />
                    <RANKING order="4" place="4" resultid="2608" />
                    <RANKING order="5" place="5" resultid="2436" />
                    <RANKING order="6" place="6" resultid="2496" />
                    <RANKING order="7" place="-1" resultid="5442" />
                    <RANKING order="8" place="-1" resultid="4011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4303" />
                    <RANKING order="2" place="2" resultid="5534" />
                    <RANKING order="3" place="3" resultid="5777" />
                    <RANKING order="4" place="4" resultid="3133" />
                    <RANKING order="5" place="5" resultid="4923" />
                    <RANKING order="6" place="6" resultid="5451" />
                    <RANKING order="7" place="7" resultid="2682" />
                    <RANKING order="8" place="8" resultid="3164" />
                    <RANKING order="9" place="-1" resultid="6069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4954" />
                    <RANKING order="2" place="2" resultid="3458" />
                    <RANKING order="3" place="3" resultid="3644" />
                    <RANKING order="4" place="4" resultid="5937" />
                    <RANKING order="5" place="5" resultid="5929" />
                    <RANKING order="6" place="6" resultid="2689" />
                    <RANKING order="7" place="7" resultid="5961" />
                    <RANKING order="8" place="8" resultid="3378" />
                    <RANKING order="9" place="9" resultid="3602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2405" />
                    <RANKING order="2" place="2" resultid="4813" />
                    <RANKING order="3" place="3" resultid="5492" />
                    <RANKING order="4" place="4" resultid="3593" />
                    <RANKING order="5" place="-1" resultid="4208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4915" />
                    <RANKING order="2" place="2" resultid="3612" />
                    <RANKING order="3" place="-1" resultid="3585" />
                    <RANKING order="4" place="-1" resultid="4246" />
                    <RANKING order="5" place="-1" resultid="4567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3412" />
                    <RANKING order="2" place="2" resultid="4639" />
                    <RANKING order="3" place="3" resultid="4977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1124" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1125" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7390" daytime="12:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7391" daytime="12:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7392" daytime="12:49" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7393" daytime="12:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7394" daytime="12:59" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7395" daytime="13:03" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7396" daytime="13:07" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7397" daytime="13:11" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7398" daytime="13:14" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7399" daytime="13:18" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7400" daytime="13:21" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7401" daytime="13:24" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7402" daytime="13:28" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7403" daytime="13:31" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7404" daytime="13:34" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7405" daytime="13:37" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7406" daytime="13:40" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7407" daytime="13:43" number="18" order="18" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1126" daytime="13:46" gender="X" number="5" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1143" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5261" />
                    <RANKING order="2" place="2" resultid="4356" />
                    <RANKING order="3" place="3" resultid="6389" />
                    <RANKING order="4" place="4" resultid="3781" />
                    <RANKING order="5" place="5" resultid="5395" />
                    <RANKING order="6" place="6" resultid="6391" />
                    <RANKING order="7" place="-1" resultid="5842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5541" />
                    <RANKING order="2" place="2" resultid="4944" />
                    <RANKING order="3" place="3" resultid="3782" />
                    <RANKING order="4" place="4" resultid="4349" />
                    <RANKING order="5" place="5" resultid="5624" />
                    <RANKING order="6" place="-1" resultid="6279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4574" />
                    <RANKING order="2" place="2" resultid="5543" />
                    <RANKING order="3" place="3" resultid="6278" />
                    <RANKING order="4" place="4" resultid="3698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4576" />
                    <RANKING order="2" place="-1" resultid="3419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2323" agemax="319" agemin="280" name="F: 280 - 319 lat " calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="359" agemin="320" name="G: 320 - 359 lat " calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7408" daytime="13:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7409" daytime="13:49" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7410" daytime="13:53" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7411" daytime="13:55" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="13:58" gender="F" number="6" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2698" />
                    <RANKING order="2" place="2" resultid="5075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5813" />
                    <RANKING order="2" place="2" resultid="5586" />
                    <RANKING order="3" place="3" resultid="4217" />
                    <RANKING order="4" place="4" resultid="4128" />
                    <RANKING order="5" place="-1" resultid="4081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5352" />
                    <RANKING order="2" place="2" resultid="4332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2814" />
                    <RANKING order="2" place="2" resultid="3708" />
                    <RANKING order="3" place="3" resultid="6053" />
                    <RANKING order="4" place="4" resultid="4265" />
                    <RANKING order="5" place="5" resultid="7069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4713" />
                    <RANKING order="2" place="2" resultid="3724" />
                    <RANKING order="3" place="3" resultid="7245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3470" />
                    <RANKING order="2" place="2" resultid="4276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4472" />
                    <RANKING order="2" place="2" resultid="5597" />
                    <RANKING order="3" place="3" resultid="4086" />
                    <RANKING order="4" place="4" resultid="5663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5059" />
                    <RANKING order="2" place="-1" resultid="3620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1161" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1162" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1163" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1164" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7902" daytime="13:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7903" daytime="14:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7904" daytime="14:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7905" daytime="14:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7906" daytime="15:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="15:11" gender="M" number="7" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1166" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7193" />
                    <RANKING order="2" place="2" resultid="3430" />
                    <RANKING order="3" place="3" resultid="7945" />
                    <RANKING order="4" place="-1" resultid="6065" />
                    <RANKING order="5" place="-1" resultid="7927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3478" />
                    <RANKING order="2" place="2" resultid="6176" />
                    <RANKING order="3" place="-1" resultid="3181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4627" />
                    <RANKING order="2" place="2" resultid="2543" />
                    <RANKING order="3" place="3" resultid="4122" />
                    <RANKING order="4" place="4" resultid="2556" />
                    <RANKING order="5" place="5" resultid="5027" />
                    <RANKING order="6" place="-1" resultid="4972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3207" />
                    <RANKING order="2" place="2" resultid="4421" />
                    <RANKING order="3" place="3" resultid="5314" />
                    <RANKING order="4" place="4" resultid="2804" />
                    <RANKING order="5" place="5" resultid="5142" />
                    <RANKING order="6" place="6" resultid="2731" />
                    <RANKING order="7" place="7" resultid="2930" />
                    <RANKING order="8" place="8" resultid="5826" />
                    <RANKING order="9" place="9" resultid="5867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3452" />
                    <RANKING order="2" place="2" resultid="2451" />
                    <RANKING order="3" place="3" resultid="3769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7158" />
                    <RANKING order="2" place="2" resultid="3048" />
                    <RANKING order="3" place="3" resultid="2580" />
                    <RANKING order="4" place="4" resultid="3801" />
                    <RANKING order="5" place="5" resultid="5761" />
                    <RANKING order="6" place="6" resultid="4103" />
                    <RANKING order="7" place="7" resultid="4804" />
                    <RANKING order="8" place="8" resultid="4045" />
                    <RANKING order="9" place="9" resultid="4547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6231" />
                    <RANKING order="2" place="2" resultid="2497" />
                    <RANKING order="3" place="3" resultid="3510" />
                    <RANKING order="4" place="4" resultid="4405" />
                    <RANKING order="5" place="5" resultid="2573" />
                    <RANKING order="6" place="6" resultid="4558" />
                    <RANKING order="7" place="7" resultid="4152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4690" />
                    <RANKING order="2" place="2" resultid="3942" />
                    <RANKING order="3" place="3" resultid="2683" />
                    <RANKING order="4" place="4" resultid="6442" />
                    <RANKING order="5" place="5" resultid="2677" />
                    <RANKING order="6" place="6" resultid="6226" />
                    <RANKING order="7" place="7" resultid="5044" />
                    <RANKING order="8" place="8" resultid="5253" />
                    <RANKING order="9" place="-1" resultid="2845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6114" />
                    <RANKING order="2" place="2" resultid="3395" />
                    <RANKING order="3" place="3" resultid="3645" />
                    <RANKING order="4" place="4" resultid="2427" />
                    <RANKING order="5" place="5" resultid="7237" />
                    <RANKING order="6" place="-1" resultid="2392" />
                    <RANKING order="7" place="-1" resultid="3603" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2854" />
                    <RANKING order="2" place="2" resultid="6027" />
                    <RANKING order="3" place="-1" resultid="4481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6132" />
                    <RANKING order="2" place="2" resultid="7936" />
                    <RANKING order="3" place="-1" resultid="4527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1180" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1181" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7907" daytime="15:11" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7908" daytime="15:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7909" daytime="16:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7910" daytime="17:01" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7911" daytime="17:27" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7912" daytime="17:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7913" daytime="18:16" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7914" daytime="18:39" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7915" daytime="19:02" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7916" daytime="19:23" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7917" daytime="19:44" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2014-11-15" daytime="08:00" name="II Blok (Sobota)" number="2" warmupfrom="07:00">
          <EVENTS>
            <EVENT eventid="1183" daytime="08:00" gender="F" number="8" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1184" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7216" />
                    <RANKING order="2" place="2" resultid="2699" />
                    <RANKING order="3" place="3" resultid="3881" />
                    <RANKING order="4" place="4" resultid="3948" />
                    <RANKING order="5" place="5" resultid="7325" />
                    <RANKING order="6" place="-1" resultid="7318" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2362" />
                    <RANKING order="2" place="2" resultid="7135" />
                    <RANKING order="3" place="3" resultid="5814" />
                    <RANKING order="4" place="4" resultid="4499" />
                    <RANKING order="5" place="5" resultid="4129" />
                    <RANKING order="6" place="6" resultid="2525" />
                    <RANKING order="7" place="7" resultid="4257" />
                    <RANKING order="8" place="8" resultid="2782" />
                    <RANKING order="9" place="-1" resultid="2711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7175" />
                    <RANKING order="2" place="2" resultid="3161" />
                    <RANKING order="3" place="3" resultid="5013" />
                    <RANKING order="4" place="4" resultid="4286" />
                    <RANKING order="5" place="5" resultid="6361" />
                    <RANKING order="6" place="6" resultid="5528" />
                    <RANKING order="7" place="7" resultid="2823" />
                    <RANKING order="8" place="-1" resultid="5835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3709" />
                    <RANKING order="2" place="2" resultid="3733" />
                    <RANKING order="3" place="3" resultid="5017" />
                    <RANKING order="4" place="4" resultid="3909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5504" />
                    <RANKING order="2" place="2" resultid="5510" />
                    <RANKING order="3" place="3" resultid="3835" />
                    <RANKING order="4" place="4" resultid="6207" />
                    <RANKING order="5" place="5" resultid="4427" />
                    <RANKING order="6" place="6" resultid="3527" />
                    <RANKING order="7" place="7" resultid="3725" />
                    <RANKING order="8" place="8" resultid="5708" />
                    <RANKING order="9" place="9" resultid="7246" />
                    <RANKING order="10" place="10" resultid="5581" />
                    <RANKING order="11" place="-1" resultid="6367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4396" />
                    <RANKING order="2" place="2" resultid="2830" />
                    <RANKING order="3" place="3" resultid="3840" />
                    <RANKING order="4" place="4" resultid="6045" />
                    <RANKING order="5" place="5" resultid="3893" />
                    <RANKING order="6" place="6" resultid="6380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5435" />
                    <RANKING order="2" place="2" resultid="6091" />
                    <RANKING order="3" place="3" resultid="7849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5323" />
                    <RANKING order="2" place="2" resultid="4682" />
                    <RANKING order="3" place="3" resultid="3504" />
                    <RANKING order="4" place="-1" resultid="4464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4902" />
                    <RANKING order="2" place="2" resultid="3387" />
                    <RANKING order="3" place="3" resultid="3573" />
                    <RANKING order="4" place="-1" resultid="3561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6098" />
                    <RANKING order="2" place="2" resultid="4703" />
                    <RANKING order="3" place="3" resultid="5347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4727" />
                    <RANKING order="2" place="2" resultid="5784" />
                    <RANKING order="3" place="3" resultid="2473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1197" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1198" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1199" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7431" daytime="08:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7432" daytime="08:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7433" daytime="08:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7434" daytime="08:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7435" daytime="08:07" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7436" daytime="08:08" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7437" daytime="08:09" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7438" daytime="08:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7439" daytime="08:11" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7440" daytime="08:12" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7441" daytime="08:14" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1200" daytime="08:15" gender="M" number="9" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1201" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7183" />
                    <RANKING order="2" place="2" resultid="7199" />
                    <RANKING order="3" place="3" resultid="3431" />
                    <RANKING order="4" place="4" resultid="2481" />
                    <RANKING order="5" place="5" resultid="2505" />
                    <RANKING order="6" place="6" resultid="7208" />
                    <RANKING order="7" place="7" resultid="6165" />
                    <RANKING order="8" place="8" resultid="7063" />
                    <RANKING order="9" place="9" resultid="4866" />
                    <RANKING order="10" place="-1" resultid="2638" />
                    <RANKING order="11" place="-1" resultid="6355" />
                    <RANKING order="12" place="-1" resultid="6478" />
                    <RANKING order="13" place="-1" resultid="7152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5789" />
                    <RANKING order="2" place="2" resultid="6158" />
                    <RANKING order="3" place="3" resultid="6427" />
                    <RANKING order="4" place="4" resultid="5702" />
                    <RANKING order="5" place="5" resultid="5087" />
                    <RANKING order="6" place="6" resultid="7143" />
                    <RANKING order="7" place="7" resultid="5716" />
                    <RANKING order="8" place="8" resultid="5185" />
                    <RANKING order="9" place="9" resultid="2737" />
                    <RANKING order="10" place="-1" resultid="2974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3027" />
                    <RANKING order="2" place="2" resultid="2563" />
                    <RANKING order="3" place="3" resultid="2586" />
                    <RANKING order="4" place="4" resultid="5909" />
                    <RANKING order="5" place="5" resultid="5861" />
                    <RANKING order="6" place="6" resultid="6347" />
                    <RANKING order="7" place="7" resultid="6333" />
                    <RANKING order="8" place="8" resultid="5946" />
                    <RANKING order="9" place="9" resultid="2978" />
                    <RANKING order="10" place="-1" resultid="2937" />
                    <RANKING order="11" place="-1" resultid="2945" />
                    <RANKING order="12" place="-1" resultid="2969" />
                    <RANKING order="13" place="-1" resultid="5198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3435" />
                    <RANKING order="2" place="2" resultid="4787" />
                    <RANKING order="3" place="3" resultid="5476" />
                    <RANKING order="4" place="4" resultid="3142" />
                    <RANKING order="5" place="5" resultid="5954" />
                    <RANKING order="6" place="6" resultid="4268" />
                    <RANKING order="7" place="7" resultid="6151" />
                    <RANKING order="8" place="8" resultid="6301" />
                    <RANKING order="9" place="9" resultid="5868" />
                    <RANKING order="10" place="10" resultid="3776" />
                    <RANKING order="11" place="11" resultid="4513" />
                    <RANKING order="12" place="-1" resultid="2398" />
                    <RANKING order="13" place="-1" resultid="2922" />
                    <RANKING order="14" place="-1" resultid="3989" />
                    <RANKING order="15" place="-1" resultid="5827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5615" />
                    <RANKING order="2" place="2" resultid="3829" />
                    <RANKING order="3" place="3" resultid="3178" />
                    <RANKING order="4" place="4" resultid="5246" />
                    <RANKING order="5" place="5" resultid="5821" />
                    <RANKING order="6" place="-1" resultid="3173" />
                    <RANKING order="7" place="-1" resultid="4067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5134" />
                    <RANKING order="2" place="2" resultid="5680" />
                    <RANKING order="3" place="3" resultid="4966" />
                    <RANKING order="4" place="4" resultid="2581" />
                    <RANKING order="5" place="5" resultid="4096" />
                    <RANKING order="6" place="6" resultid="4859" />
                    <RANKING order="7" place="7" resultid="5762" />
                    <RANKING order="8" place="8" resultid="5654" />
                    <RANKING order="9" place="9" resultid="5382" />
                    <RANKING order="10" place="10" resultid="3190" />
                    <RANKING order="11" place="-1" resultid="3049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6018" />
                    <RANKING order="2" place="2" resultid="6433" />
                    <RANKING order="3" place="3" resultid="4621" />
                    <RANKING order="4" place="4" resultid="6424" />
                    <RANKING order="5" place="5" resultid="4506" />
                    <RANKING order="6" place="6" resultid="2437" />
                    <RANKING order="7" place="7" resultid="3821" />
                    <RANKING order="8" place="8" resultid="3680" />
                    <RANKING order="9" place="9" resultid="6247" />
                    <RANKING order="10" place="10" resultid="4238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6104" />
                    <RANKING order="2" place="2" resultid="4304" />
                    <RANKING order="3" place="3" resultid="4664" />
                    <RANKING order="4" place="4" resultid="2864" />
                    <RANKING order="5" place="5" resultid="4749" />
                    <RANKING order="6" place="6" resultid="2684" />
                    <RANKING order="7" place="7" resultid="6219" />
                    <RANKING order="8" place="8" resultid="4924" />
                    <RANKING order="9" place="9" resultid="5045" />
                    <RANKING order="10" place="-1" resultid="5254" />
                    <RANKING order="11" place="-1" resultid="4450" />
                    <RANKING order="12" place="-1" resultid="4691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4955" />
                    <RANKING order="2" place="2" resultid="5307" />
                    <RANKING order="3" place="3" resultid="2393" />
                    <RANKING order="4" place="4" resultid="3646" />
                    <RANKING order="5" place="5" resultid="2428" />
                    <RANKING order="6" place="6" resultid="5962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4708" />
                    <RANKING order="2" place="2" resultid="4814" />
                    <RANKING order="3" place="3" resultid="4761" />
                    <RANKING order="4" place="4" resultid="5875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4916" />
                    <RANKING order="2" place="2" resultid="3613" />
                    <RANKING order="3" place="3" resultid="5892" />
                    <RANKING order="4" place="4" resultid="4024" />
                    <RANKING order="5" place="5" resultid="4528" />
                    <RANKING order="6" place="6" resultid="3629" />
                    <RANKING order="7" place="-1" resultid="5006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4640" />
                    <RANKING order="2" place="-1" resultid="5795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3869" />
                    <RANKING order="2" place="-1" resultid="3373" />
                    <RANKING order="3" place="-1" resultid="4403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1215" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1216" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7442" daytime="08:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7443" daytime="08:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7444" daytime="08:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7445" daytime="08:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7446" daytime="08:21" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7447" daytime="08:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7448" daytime="08:23" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7449" daytime="08:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7450" daytime="08:26" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7451" daytime="08:27" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7452" daytime="08:28" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7453" daytime="08:29" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7454" daytime="08:30" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7455" daytime="08:31" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7456" daytime="08:32" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7457" daytime="08:33" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7458" daytime="08:34" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7459" daytime="08:35" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7460" daytime="08:36" number="19" order="19" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1217" daytime="08:37" gender="F" number="10" order="13" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1218" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7190" />
                    <RANKING order="2" place="2" resultid="2663" />
                    <RANKING order="3" place="3" resultid="5853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5068" />
                    <RANKING order="2" place="2" resultid="5971" />
                    <RANKING order="3" place="3" resultid="2716" />
                    <RANKING order="4" place="4" resultid="5159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5922" />
                    <RANKING order="2" place="2" resultid="4146" />
                    <RANKING order="3" place="3" resultid="4113" />
                    <RANKING order="4" place="4" resultid="4333" />
                    <RANKING order="5" place="5" resultid="6038" />
                    <RANKING order="6" place="-1" resultid="5697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5916" />
                    <RANKING order="2" place="2" resultid="7070" />
                    <RANKING order="3" place="3" resultid="3910" />
                    <RANKING order="4" place="-1" resultid="5420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4714" />
                    <RANKING order="2" place="2" resultid="5126" />
                    <RANKING order="3" place="3" resultid="5809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4850" />
                    <RANKING order="2" place="2" resultid="4277" />
                    <RANKING order="3" place="3" resultid="3498" />
                    <RANKING order="4" place="4" resultid="3812" />
                    <RANKING order="5" place="5" resultid="3894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4909" />
                    <RANKING order="2" place="2" resultid="5094" />
                    <RANKING order="3" place="3" resultid="6092" />
                    <RANKING order="4" place="4" resultid="2517" />
                    <RANKING order="5" place="5" resultid="5385" />
                    <RANKING order="6" place="6" resultid="5598" />
                    <RANKING order="7" place="7" resultid="4020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4541" />
                    <RANKING order="2" place="2" resultid="4895" />
                    <RANKING order="3" place="3" resultid="3672" />
                    <RANKING order="4" place="4" resultid="3663" />
                    <RANKING order="5" place="5" resultid="2568" />
                    <RANKING order="6" place="6" resultid="6077" />
                    <RANKING order="7" place="7" resultid="2871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3405" />
                    <RANKING order="2" place="2" resultid="4037" />
                    <RANKING order="3" place="3" resultid="4439" />
                    <RANKING order="4" place="4" resultid="4016" />
                    <RANKING order="5" place="5" resultid="3979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4491" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4736" />
                    <RANKING order="2" place="2" resultid="3567" />
                    <RANKING order="3" place="3" resultid="3548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1231" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1232" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1233" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7461" daytime="08:37" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7462" daytime="08:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7463" daytime="08:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7464" daytime="08:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7465" daytime="09:01" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7466" daytime="09:06" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7467" daytime="09:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7468" daytime="09:14" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7469" daytime="09:17" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1234" daytime="09:21" gender="M" number="11" order="14" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1235" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6339" />
                    <RANKING order="2" place="2" resultid="7228" />
                    <RANKING order="3" place="3" resultid="4241" />
                    <RANKING order="4" place="-1" resultid="2639" />
                    <RANKING order="5" place="-1" resultid="6486" />
                    <RANKING order="6" place="-1" resultid="7153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4381" />
                    <RANKING order="2" place="2" resultid="5689" />
                    <RANKING order="3" place="3" resultid="5180" />
                    <RANKING order="4" place="4" resultid="2789" />
                    <RANKING order="5" place="5" resultid="5167" />
                    <RANKING order="6" place="6" resultid="5152" />
                    <RANKING order="7" place="7" resultid="2748" />
                    <RANKING order="8" place="8" resultid="4418" />
                    <RANKING order="9" place="-1" resultid="4614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3997" />
                    <RANKING order="2" place="2" resultid="4326" />
                    <RANKING order="3" place="3" resultid="2907" />
                    <RANKING order="4" place="4" resultid="2954" />
                    <RANKING order="5" place="5" resultid="5064" />
                    <RANKING order="6" place="6" resultid="5028" />
                    <RANKING order="7" place="7" resultid="3961" />
                    <RANKING order="8" place="8" resultid="2742" />
                    <RANKING order="9" place="9" resultid="3242" />
                    <RANKING order="10" place="10" resultid="2889" />
                    <RANKING order="11" place="-1" resultid="2544" />
                    <RANKING order="12" place="-1" resultid="5900" />
                    <RANKING order="13" place="-1" resultid="5910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5980" />
                    <RANKING order="2" place="2" resultid="3208" />
                    <RANKING order="3" place="3" resultid="5516" />
                    <RANKING order="4" place="4" resultid="5300" />
                    <RANKING order="5" place="5" resultid="5143" />
                    <RANKING order="6" place="6" resultid="4841" />
                    <RANKING order="7" place="7" resultid="3966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3031" />
                    <RANKING order="2" place="2" resultid="3236" />
                    <RANKING order="3" place="3" resultid="4606" />
                    <RANKING order="4" place="4" resultid="3742" />
                    <RANKING order="5" place="5" resultid="2879" />
                    <RANKING order="6" place="6" resultid="6120" />
                    <RANKING order="7" place="7" resultid="3816" />
                    <RANKING order="8" place="8" resultid="3225" />
                    <RANKING order="9" place="9" resultid="5712" />
                    <RANKING order="10" place="10" resultid="5768" />
                    <RANKING order="11" place="11" resultid="5000" />
                    <RANKING order="12" place="-1" resultid="2809" />
                    <RANKING order="13" place="-1" resultid="3901" />
                    <RANKING order="14" place="-1" resultid="5592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3825" />
                    <RANKING order="2" place="2" resultid="2373" />
                    <RANKING order="3" place="3" resultid="4931" />
                    <RANKING order="4" place="4" resultid="3972" />
                    <RANKING order="5" place="5" resultid="5498" />
                    <RANKING order="6" place="6" resultid="3579" />
                    <RANKING order="7" place="7" resultid="6253" />
                    <RANKING order="8" place="8" resultid="4104" />
                    <RANKING order="9" place="9" resultid="4993" />
                    <RANKING order="10" place="10" resultid="4676" />
                    <RANKING order="11" place="11" resultid="4555" />
                    <RANKING order="12" place="-1" resultid="3886" />
                    <RANKING order="13" place="-1" resultid="5099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5376" />
                    <RANKING order="2" place="2" resultid="2609" />
                    <RANKING order="3" place="3" resultid="6240" />
                    <RANKING order="4" place="4" resultid="4559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5778" />
                    <RANKING order="2" place="2" resultid="3134" />
                    <RANKING order="3" place="3" resultid="7059" />
                    <RANKING order="4" place="4" resultid="5452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4630" />
                    <RANKING order="2" place="2" resultid="3459" />
                    <RANKING order="3" place="3" resultid="3369" />
                    <RANKING order="4" place="4" resultid="2690" />
                    <RANKING order="5" place="5" resultid="5930" />
                    <RANKING order="6" place="6" resultid="3604" />
                    <RANKING order="7" place="-1" resultid="3862" />
                    <RANKING order="8" place="-1" resultid="6112" />
                    <RANKING order="9" place="-1" resultid="7238" />
                    <RANKING order="10" place="-1" resultid="3379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5424" />
                    <RANKING order="2" place="2" resultid="5465" />
                    <RANKING order="3" place="3" resultid="3594" />
                    <RANKING order="4" place="4" resultid="5876" />
                    <RANKING order="5" place="5" resultid="4209" />
                    <RANKING order="6" place="6" resultid="5881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4731" />
                    <RANKING order="2" place="2" resultid="4025" />
                    <RANKING order="3" place="3" resultid="3586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3413" />
                    <RANKING order="2" place="2" resultid="4978" />
                    <RANKING order="3" place="3" resultid="5796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3374" />
                    <RANKING order="2" place="2" resultid="7179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1249" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1250" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7470" daytime="09:21" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7471" daytime="09:27" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7472" daytime="09:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7473" daytime="09:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7474" daytime="09:43" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7475" daytime="09:47" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7476" daytime="09:51" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7477" daytime="09:55" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7478" daytime="09:59" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7479" daytime="10:02" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7480" daytime="10:06" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7481" daytime="10:09" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7482" daytime="10:13" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7483" daytime="10:16" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7484" daytime="10:19" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7485" daytime="10:23" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1251" daytime="10:26" gender="F" number="12" order="15" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1252" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2700" />
                    <RANKING order="2" place="2" resultid="7217" />
                    <RANKING order="3" place="3" resultid="5076" />
                    <RANKING order="4" place="4" resultid="6447" />
                    <RANKING order="5" place="-1" resultid="6287" />
                    <RANKING order="6" place="-1" resultid="6458" />
                    <RANKING order="7" place="-1" resultid="7319" />
                    <RANKING order="8" place="-1" resultid="7326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7136" />
                    <RANKING order="2" place="2" resultid="5815" />
                    <RANKING order="3" place="3" resultid="4218" />
                    <RANKING order="4" place="4" resultid="5069" />
                    <RANKING order="5" place="5" resultid="2528" />
                    <RANKING order="6" place="6" resultid="3928" />
                    <RANKING order="7" place="7" resultid="6384" />
                    <RANKING order="8" place="8" resultid="3252" />
                    <RANKING order="9" place="9" resultid="2783" />
                    <RANKING order="10" place="10" resultid="4986" />
                    <RANKING order="11" place="11" resultid="2801" />
                    <RANKING order="12" place="12" resultid="5051" />
                    <RANKING order="13" place="13" resultid="4082" />
                    <RANKING order="14" place="-1" resultid="2712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4948" />
                    <RANKING order="2" place="2" resultid="3150" />
                    <RANKING order="3" place="3" resultid="5353" />
                    <RANKING order="4" place="4" resultid="2824" />
                    <RANKING order="5" place="5" resultid="4720" />
                    <RANKING order="6" place="6" resultid="5035" />
                    <RANKING order="7" place="7" resultid="6125" />
                    <RANKING order="8" place="8" resultid="5529" />
                    <RANKING order="9" place="9" resultid="6039" />
                    <RANKING order="10" place="10" resultid="6377" />
                    <RANKING order="11" place="11" resultid="6372" />
                    <RANKING order="12" place="12" resultid="4434" />
                    <RANKING order="13" place="-1" resultid="5836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2815" />
                    <RANKING order="2" place="2" resultid="3717" />
                    <RANKING order="3" place="3" resultid="3734" />
                    <RANKING order="4" place="4" resultid="6054" />
                    <RANKING order="5" place="5" resultid="7071" />
                    <RANKING order="6" place="6" resultid="5018" />
                    <RANKING order="7" place="7" resultid="3658" />
                    <RANKING order="8" place="8" resultid="4520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4412" />
                    <RANKING order="2" place="2" resultid="7247" />
                    <RANKING order="3" place="3" resultid="5605" />
                    <RANKING order="4" place="4" resultid="5802" />
                    <RANKING order="5" place="5" resultid="2672" />
                    <RANKING order="6" place="-1" resultid="5391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3471" />
                    <RANKING order="2" place="2" resultid="4278" />
                    <RANKING order="3" place="3" resultid="2831" />
                    <RANKING order="4" place="4" resultid="3841" />
                    <RANKING order="5" place="-1" resultid="3809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5485" />
                    <RANKING order="2" place="2" resultid="6197" />
                    <RANKING order="3" place="3" resultid="5664" />
                    <RANKING order="4" place="4" resultid="6085" />
                    <RANKING order="5" place="-1" resultid="4021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4683" />
                    <RANKING order="2" place="2" resultid="6188" />
                    <RANKING order="3" place="3" resultid="3505" />
                    <RANKING order="4" place="4" resultid="2838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4903" />
                    <RANKING order="2" place="2" resultid="4745" />
                    <RANKING order="3" place="3" resultid="5457" />
                    <RANKING order="4" place="4" resultid="3540" />
                    <RANKING order="5" place="-1" resultid="3562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6099" />
                    <RANKING order="2" place="2" resultid="5348" />
                    <RANKING order="3" place="3" resultid="5060" />
                    <RANKING order="4" place="4" resultid="4492" />
                    <RANKING order="5" place="5" resultid="3554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4728" />
                    <RANKING order="2" place="2" resultid="3568" />
                    <RANKING order="3" place="3" resultid="3549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1265" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1266" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1267" agemax="-1" agemin="95" name="O: 95 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5675" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7486" daytime="10:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7487" daytime="10:29" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7488" daytime="10:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7489" daytime="10:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7490" daytime="10:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7491" daytime="10:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7492" daytime="10:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7493" daytime="10:42" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7494" daytime="10:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7495" daytime="10:45" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7496" daytime="10:47" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7497" daytime="10:49" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7498" daytime="10:50" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1268" daytime="10:52" gender="M" number="13" order="16" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1269" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7184" />
                    <RANKING order="2" place="2" resultid="2506" />
                    <RANKING order="3" place="3" resultid="2480" />
                    <RANKING order="4" place="4" resultid="2601" />
                    <RANKING order="5" place="5" resultid="5659" />
                    <RANKING order="6" place="6" resultid="6356" />
                    <RANKING order="7" place="7" resultid="4136" />
                    <RANKING order="8" place="-1" resultid="2456" />
                    <RANKING order="9" place="-1" resultid="6479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1270" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7223" />
                    <RANKING order="2" place="2" resultid="5790" />
                    <RANKING order="3" place="3" resultid="5671" />
                    <RANKING order="4" place="4" resultid="5106" />
                    <RANKING order="5" place="5" resultid="4457" />
                    <RANKING order="6" place="6" resultid="2790" />
                    <RANKING order="7" place="7" resultid="2738" />
                    <RANKING order="8" place="8" resultid="2763" />
                    <RANKING order="9" place="9" resultid="5119" />
                    <RANKING order="10" place="10" resultid="3230" />
                    <RANKING order="11" place="-1" resultid="2975" />
                    <RANKING order="12" place="-1" resultid="4224" />
                    <RANKING order="13" place="-1" resultid="5186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2963" />
                    <RANKING order="2" place="2" resultid="2724" />
                    <RANKING order="3" place="3" resultid="6465" />
                    <RANKING order="4" place="4" resultid="3878" />
                    <RANKING order="5" place="5" resultid="6334" />
                    <RANKING order="6" place="6" resultid="3956" />
                    <RANKING order="7" place="7" resultid="6319" />
                    <RANKING order="8" place="8" resultid="2902" />
                    <RANKING order="9" place="9" resultid="6460" />
                    <RANKING order="10" place="10" resultid="5862" />
                    <RANKING order="11" place="11" resultid="3247" />
                    <RANKING order="12" place="12" resultid="4318" />
                    <RANKING order="13" place="13" resultid="5190" />
                    <RANKING order="14" place="14" resultid="4973" />
                    <RANKING order="15" place="15" resultid="6328" />
                    <RANKING order="16" place="16" resultid="2970" />
                    <RANKING order="17" place="17" resultid="2757" />
                    <RANKING order="18" place="18" resultid="4754" />
                    <RANKING order="19" place="-1" resultid="6062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6312" />
                    <RANKING order="2" place="2" resultid="5955" />
                    <RANKING order="3" place="3" resultid="4788" />
                    <RANKING order="4" place="4" resultid="2913" />
                    <RANKING order="5" place="5" resultid="5080" />
                    <RANKING order="6" place="6" resultid="4939" />
                    <RANKING order="7" place="7" resultid="7128" />
                    <RANKING order="8" place="8" resultid="4093" />
                    <RANKING order="9" place="8" resultid="5315" />
                    <RANKING order="10" place="10" resultid="4422" />
                    <RANKING order="11" place="11" resultid="2982" />
                    <RANKING order="12" place="12" resultid="2931" />
                    <RANKING order="13" place="13" resultid="2732" />
                    <RANKING order="14" place="14" resultid="5149" />
                    <RANKING order="15" place="15" resultid="5022" />
                    <RANKING order="16" place="16" resultid="3777" />
                    <RANKING order="17" place="17" resultid="2884" />
                    <RANKING order="18" place="18" resultid="4672" />
                    <RANKING order="19" place="19" resultid="4550" />
                    <RANKING order="20" place="20" resultid="6030" />
                    <RANKING order="21" place="21" resultid="6323" />
                    <RANKING order="22" place="-1" resultid="6294" />
                    <RANKING order="23" place="-1" resultid="6421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4796" />
                    <RANKING order="2" place="2" resultid="5370" />
                    <RANKING order="3" place="3" resultid="4295" />
                    <RANKING order="4" place="4" resultid="3761" />
                    <RANKING order="5" place="5" resultid="4389" />
                    <RANKING order="6" place="6" resultid="3453" />
                    <RANKING order="7" place="7" resultid="5247" />
                    <RANKING order="8" place="8" resultid="5039" />
                    <RANKING order="9" place="9" resultid="4312" />
                    <RANKING order="10" place="10" resultid="5610" />
                    <RANKING order="11" place="11" resultid="4322" />
                    <RANKING order="12" place="12" resultid="6121" />
                    <RANKING order="13" place="13" resultid="3923" />
                    <RANKING order="14" place="14" resultid="3770" />
                    <RANKING order="15" place="15" resultid="4823" />
                    <RANKING order="16" place="16" resultid="4339" />
                    <RANKING order="17" place="17" resultid="3687" />
                    <RANKING order="18" place="18" resultid="3693" />
                    <RANKING order="19" place="19" resultid="5822" />
                    <RANKING order="20" place="20" resultid="5001" />
                    <RANKING order="21" place="21" resultid="6305" />
                    <RANKING order="22" place="-1" resultid="7314" />
                    <RANKING order="23" place="-1" resultid="3174" />
                    <RANKING order="24" place="-1" resultid="3755" />
                    <RANKING order="25" place="-1" resultid="4068" />
                    <RANKING order="26" place="-1" resultid="5360" />
                    <RANKING order="27" place="-1" resultid="5573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3041" />
                    <RANKING order="2" place="2" resultid="3491" />
                    <RANKING order="3" place="3" resultid="3515" />
                    <RANKING order="4" place="4" resultid="2490" />
                    <RANKING order="5" place="5" resultid="6259" />
                    <RANKING order="6" place="6" resultid="2647" />
                    <RANKING order="7" place="7" resultid="3846" />
                    <RANKING order="8" place="8" resultid="3936" />
                    <RANKING order="9" place="9" resultid="4860" />
                    <RANKING order="10" place="10" resultid="5763" />
                    <RANKING order="11" place="11" resultid="2656" />
                    <RANKING order="12" place="12" resultid="2374" />
                    <RANKING order="13" place="13" resultid="4105" />
                    <RANKING order="14" place="14" resultid="4046" />
                    <RANKING order="15" place="15" resultid="4636" />
                    <RANKING order="16" place="16" resultid="3637" />
                    <RANKING order="17" place="17" resultid="4805" />
                    <RANKING order="18" place="18" resultid="4516" />
                    <RANKING order="19" place="19" resultid="3191" />
                    <RANKING order="20" place="-1" resultid="3050" />
                    <RANKING order="21" place="-1" resultid="3218" />
                    <RANKING order="22" place="-1" resultid="5100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2594" />
                    <RANKING order="2" place="2" resultid="2534" />
                    <RANKING order="3" place="3" resultid="6248" />
                    <RANKING order="4" place="4" resultid="4832" />
                    <RANKING order="5" place="5" resultid="3806" />
                    <RANKING order="6" place="6" resultid="3681" />
                    <RANKING order="7" place="7" resultid="5523" />
                    <RANKING order="8" place="8" resultid="4153" />
                    <RANKING order="9" place="9" resultid="4009" />
                    <RANKING order="10" place="-1" resultid="4622" />
                    <RANKING order="11" place="-1" resultid="5113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4665" />
                    <RANKING order="2" place="2" resultid="2446" />
                    <RANKING order="3" place="3" resultid="4648" />
                    <RANKING order="4" place="4" resultid="6070" />
                    <RANKING order="5" place="5" resultid="2484" />
                    <RANKING order="6" place="6" resultid="5046" />
                    <RANKING order="7" place="7" resultid="6227" />
                    <RANKING order="8" place="8" resultid="3165" />
                    <RANKING order="9" place="9" resultid="5255" />
                    <RANKING order="10" place="-1" resultid="2846" />
                    <RANKING order="11" place="-1" resultid="3943" />
                    <RANKING order="12" place="-1" resultid="4451" />
                    <RANKING order="13" place="-1" resultid="5535" />
                    <RANKING order="14" place="-1" resultid="5773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2467" />
                    <RANKING order="2" place="2" resultid="2394" />
                    <RANKING order="3" place="3" resultid="5938" />
                    <RANKING order="4" place="4" resultid="5753" />
                    <RANKING order="5" place="5" resultid="3396" />
                    <RANKING order="6" place="-1" resultid="2429" />
                    <RANKING order="7" place="-1" resultid="6275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4482" />
                    <RANKING order="2" place="2" resultid="5493" />
                    <RANKING order="3" place="3" resultid="2855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5007" />
                    <RANKING order="2" place="2" resultid="6133" />
                    <RANKING order="3" place="3" resultid="5893" />
                    <RANKING order="4" place="4" resultid="4529" />
                    <RANKING order="5" place="5" resultid="4568" />
                    <RANKING order="6" place="6" resultid="3625" />
                    <RANKING order="7" place="-1" resultid="3630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4641" />
                    <RANKING order="2" place="2" resultid="5888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1283" agemax="94" agemin="90" name="N: 90 - 94 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7499" daytime="10:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7500" daytime="10:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7501" daytime="10:59" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7502" daytime="11:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7503" daytime="11:04" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7504" daytime="11:06" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7505" daytime="11:08" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7506" daytime="11:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7507" daytime="11:12" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7508" daytime="11:13" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7509" daytime="11:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7510" daytime="11:17" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7511" daytime="11:18" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7512" daytime="11:20" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7513" daytime="11:22" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7514" daytime="11:23" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7515" daytime="11:25" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7516" daytime="11:26" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7517" daytime="11:28" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7518" daytime="11:30" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="7519" daytime="11:31" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="7520" daytime="11:33" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="7521" daytime="11:34" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="7522" daytime="11:36" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="7523" daytime="11:37" number="25" order="25" status="OFFICIAL" />
                <HEAT heatid="7524" daytime="11:39" number="26" order="26" status="OFFICIAL" />
                <HEAT heatid="7525" daytime="11:40" number="27" order="27" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1285" daytime="11:42" gender="F" number="14" order="17" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1286" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7254" />
                    <RANKING order="2" place="2" resultid="2664" />
                    <RANKING order="3" place="3" resultid="7191" />
                    <RANKING order="4" place="4" resultid="5174" />
                    <RANKING order="5" place="5" resultid="3520" />
                    <RANKING order="6" place="6" resultid="3949" />
                    <RANKING order="7" place="7" resultid="7327" />
                    <RANKING order="8" place="-1" resultid="7320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2363" />
                    <RANKING order="2" place="2" resultid="4500" />
                    <RANKING order="3" place="3" resultid="5972" />
                    <RANKING order="4" place="4" resultid="4130" />
                    <RANKING order="5" place="5" resultid="3929" />
                    <RANKING order="6" place="6" resultid="5587" />
                    <RANKING order="7" place="7" resultid="2717" />
                    <RANKING order="8" place="8" resultid="5160" />
                    <RANKING order="9" place="9" resultid="2706" />
                    <RANKING order="10" place="-1" resultid="5052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4949" />
                    <RANKING order="2" place="2" resultid="3151" />
                    <RANKING order="3" place="3" resultid="5923" />
                    <RANKING order="4" place="4" resultid="5354" />
                    <RANKING order="5" place="5" resultid="4287" />
                    <RANKING order="6" place="6" resultid="6387" />
                    <RANKING order="7" place="7" resultid="6142" />
                    <RANKING order="8" place="8" resultid="5036" />
                    <RANKING order="9" place="9" resultid="6362" />
                    <RANKING order="10" place="-1" resultid="5530" />
                    <RANKING order="11" place="-1" resultid="6174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3710" />
                    <RANKING order="2" place="2" resultid="3718" />
                    <RANKING order="3" place="3" resultid="5917" />
                    <RANKING order="4" place="4" resultid="6055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5511" />
                    <RANKING order="2" place="2" resultid="5505" />
                    <RANKING order="3" place="3" resultid="5747" />
                    <RANKING order="4" place="4" resultid="5127" />
                    <RANKING order="5" place="5" resultid="3528" />
                    <RANKING order="6" place="6" resultid="3726" />
                    <RANKING order="7" place="7" resultid="6368" />
                    <RANKING order="8" place="8" resultid="5709" />
                    <RANKING order="9" place="9" resultid="5582" />
                    <RANKING order="10" place="10" resultid="2673" />
                    <RANKING order="11" place="-1" resultid="4413" />
                    <RANKING order="12" place="-1" resultid="4428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4397" />
                    <RANKING order="2" place="2" resultid="4535" />
                    <RANKING order="3" place="3" resultid="3472" />
                    <RANKING order="4" place="4" resultid="3499" />
                    <RANKING order="5" place="5" resultid="6046" />
                    <RANKING order="6" place="-1" resultid="4231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5486" />
                    <RANKING order="2" place="2" resultid="6202" />
                    <RANKING order="3" place="3" resultid="4473" />
                    <RANKING order="4" place="4" resultid="5599" />
                    <RANKING order="5" place="5" resultid="5665" />
                    <RANKING order="6" place="6" resultid="6086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4896" />
                    <RANKING order="2" place="2" resultid="6189" />
                    <RANKING order="3" place="3" resultid="5324" />
                    <RANKING order="4" place="4" resultid="3673" />
                    <RANKING order="5" place="-1" resultid="2839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3406" />
                    <RANKING order="2" place="2" resultid="5458" />
                    <RANKING order="3" place="3" resultid="3541" />
                    <RANKING order="4" place="4" resultid="4440" />
                    <RANKING order="5" place="5" resultid="3574" />
                    <RANKING order="6" place="6" resultid="3980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6023" />
                    <RANKING order="2" place="2" resultid="3555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1298" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1299" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1300" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1301" agemax="-1" agemin="95" name="O: 95 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5676" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7526" daytime="11:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7527" daytime="11:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7528" daytime="11:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7529" daytime="11:51" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7530" daytime="11:53" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7531" daytime="11:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7532" daytime="11:57" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7533" daytime="11:58" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7534" daytime="12:00" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7535" daytime="12:02" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7536" daytime="12:04" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7537" daytime="12:06" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="12:08" gender="M" number="15" order="18" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1303" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7200" />
                    <RANKING order="2" place="2" resultid="6340" />
                    <RANKING order="3" place="3" resultid="7209" />
                    <RANKING order="4" place="4" resultid="6166" />
                    <RANKING order="5" place="5" resultid="7064" />
                    <RANKING order="6" place="-1" resultid="3432" />
                    <RANKING order="7" place="-1" resultid="4004" />
                    <RANKING order="8" place="-1" resultid="6488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6428" />
                    <RANKING order="2" place="2" resultid="7144" />
                    <RANKING order="3" place="3" resultid="4382" />
                    <RANKING order="4" place="4" resultid="5703" />
                    <RANKING order="5" place="5" resultid="5168" />
                    <RANKING order="6" place="6" resultid="5088" />
                    <RANKING order="7" place="7" resultid="6159" />
                    <RANKING order="8" place="8" resultid="5717" />
                    <RANKING order="9" place="9" resultid="5153" />
                    <RANKING order="10" place="10" resultid="5649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3998" />
                    <RANKING order="2" place="2" resultid="4123" />
                    <RANKING order="3" place="3" resultid="6452" />
                    <RANKING order="4" place="4" resultid="2725" />
                    <RANKING order="5" place="5" resultid="2797" />
                    <RANKING order="6" place="6" resultid="2587" />
                    <RANKING order="7" place="7" resultid="5693" />
                    <RANKING order="8" place="8" resultid="4327" />
                    <RANKING order="9" place="9" resultid="2545" />
                    <RANKING order="10" place="10" resultid="3962" />
                    <RANKING order="11" place="11" resultid="3957" />
                    <RANKING order="12" place="12" resultid="5029" />
                    <RANKING order="13" place="13" resultid="5947" />
                    <RANKING order="14" place="14" resultid="5191" />
                    <RANKING order="15" place="15" resultid="2890" />
                    <RANKING order="16" place="16" resultid="2946" />
                    <RANKING order="17" place="17" resultid="2938" />
                    <RANKING order="18" place="-1" resultid="2897" />
                    <RANKING order="19" place="-1" resultid="2955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5981" />
                    <RANKING order="2" place="2" resultid="6152" />
                    <RANKING order="3" place="3" resultid="3143" />
                    <RANKING order="4" place="4" resultid="5477" />
                    <RANKING order="5" place="5" resultid="6313" />
                    <RANKING order="6" place="6" resultid="4269" />
                    <RANKING order="7" place="7" resultid="3990" />
                    <RANKING order="8" place="8" resultid="5081" />
                    <RANKING order="9" place="9" resultid="4940" />
                    <RANKING order="10" place="10" resultid="5316" />
                    <RANKING order="11" place="11" resultid="2923" />
                    <RANKING order="12" place="12" resultid="2983" />
                    <RANKING order="13" place="13" resultid="3749" />
                    <RANKING order="14" place="14" resultid="7129" />
                    <RANKING order="15" place="15" resultid="2919" />
                    <RANKING order="16" place="16" resultid="6031" />
                    <RANKING order="17" place="17" resultid="3967" />
                    <RANKING order="18" place="-1" resultid="5517" />
                    <RANKING order="19" place="-1" resultid="5828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4797" />
                    <RANKING order="2" place="2" resultid="4296" />
                    <RANKING order="3" place="3" resultid="5574" />
                    <RANKING order="4" place="4" resultid="3762" />
                    <RANKING order="5" place="5" resultid="3830" />
                    <RANKING order="6" place="6" resultid="5616" />
                    <RANKING order="7" place="7" resultid="5040" />
                    <RANKING order="8" place="8" resultid="4824" />
                    <RANKING order="9" place="9" resultid="5593" />
                    <RANKING order="10" place="10" resultid="2651" />
                    <RANKING order="11" place="11" resultid="6306" />
                    <RANKING order="12" place="-1" resultid="3743" />
                    <RANKING order="13" place="-1" resultid="3032" />
                    <RANKING order="14" place="-1" resultid="3237" />
                    <RANKING order="15" place="-1" resultid="3902" />
                    <RANKING order="16" place="-1" resultid="6470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5135" />
                    <RANKING order="2" place="2" resultid="3492" />
                    <RANKING order="3" place="2" resultid="5681" />
                    <RANKING order="4" place="4" resultid="4967" />
                    <RANKING order="5" place="5" resultid="3042" />
                    <RANKING order="6" place="6" resultid="3847" />
                    <RANKING order="7" place="7" resultid="2657" />
                    <RANKING order="8" place="8" resultid="2491" />
                    <RANKING order="9" place="9" resultid="4932" />
                    <RANKING order="10" place="10" resultid="5655" />
                    <RANKING order="11" place="11" resultid="5383" />
                    <RANKING order="12" place="12" resultid="4806" />
                    <RANKING order="13" place="13" resultid="4047" />
                    <RANKING order="14" place="14" resultid="3638" />
                    <RANKING order="15" place="-1" resultid="2648" />
                    <RANKING order="16" place="-1" resultid="3219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6434" />
                    <RANKING order="2" place="2" resultid="6019" />
                    <RANKING order="3" place="3" resultid="2535" />
                    <RANKING order="4" place="4" resultid="6232" />
                    <RANKING order="5" place="5" resultid="3058" />
                    <RANKING order="6" place="6" resultid="2438" />
                    <RANKING order="7" place="7" resultid="2610" />
                    <RANKING order="8" place="8" resultid="4406" />
                    <RANKING order="9" place="9" resultid="4560" />
                    <RANKING order="10" place="10" resultid="4008" />
                    <RANKING order="11" place="-1" resultid="4507" />
                    <RANKING order="12" place="-1" resultid="5114" />
                    <RANKING order="13" place="-1" resultid="5443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6105" />
                    <RANKING order="2" place="2" resultid="4305" />
                    <RANKING order="3" place="3" resultid="2865" />
                    <RANKING order="4" place="4" resultid="5779" />
                    <RANKING order="5" place="5" resultid="4649" />
                    <RANKING order="6" place="6" resultid="6221" />
                    <RANKING order="7" place="7" resultid="4925" />
                    <RANKING order="8" place="8" resultid="5453" />
                    <RANKING order="9" place="9" resultid="6071" />
                    <RANKING order="10" place="10" resultid="2552" />
                    <RANKING order="11" place="11" resultid="3166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2468" />
                    <RANKING order="2" place="2" resultid="4956" />
                    <RANKING order="3" place="3" resultid="5308" />
                    <RANKING order="4" place="4" resultid="6115" />
                    <RANKING order="5" place="5" resultid="5939" />
                    <RANKING order="6" place="6" resultid="3397" />
                    <RANKING order="7" place="7" resultid="2691" />
                    <RANKING order="8" place="8" resultid="5963" />
                    <RANKING order="9" place="-1" resultid="7239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2406" />
                    <RANKING order="2" place="2" resultid="4815" />
                    <RANKING order="3" place="3" resultid="4741" />
                    <RANKING order="4" place="4" resultid="4445" />
                    <RANKING order="5" place="5" resultid="4762" />
                    <RANKING order="6" place="6" resultid="3595" />
                    <RANKING order="7" place="-1" resultid="5425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4917" />
                    <RANKING order="2" place="2" resultid="6134" />
                    <RANKING order="3" place="3" resultid="4248" />
                    <RANKING order="4" place="4" resultid="4569" />
                    <RANKING order="5" place="5" resultid="3587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3414" />
                    <RANKING order="2" place="2" resultid="2384" />
                    <RANKING order="3" place="3" resultid="4979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1316" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1317" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1318" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7538" daytime="12:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7539" daytime="12:11" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7540" daytime="12:13" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7541" daytime="12:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7542" daytime="12:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7543" daytime="12:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7544" daytime="12:22" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7545" daytime="12:24" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7546" daytime="12:26" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7547" daytime="12:28" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7548" daytime="12:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7549" daytime="12:31" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7550" daytime="12:33" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7551" daytime="12:35" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7552" daytime="12:37" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7553" daytime="12:38" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7554" daytime="12:40" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7555" daytime="12:42" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7556" daytime="12:43" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7557" daytime="12:45" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="7558" daytime="12:47" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="7559" daytime="12:48" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="7560" daytime="12:50" number="23" order="23" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1319" daytime="12:52" gender="F" number="16" order="19" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1320" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1321" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4258" />
                    <RANKING order="2" place="2" resultid="4219" />
                    <RANKING order="3" place="3" resultid="4987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1322" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4114" />
                    <RANKING order="2" place="2" resultid="6143" />
                    <RANKING order="3" place="3" resultid="6126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1323" agemax="39" agemin="35" name="C: 35 - 39 lat" />
                <AGEGROUP agegroupid="1324" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1325" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4851" />
                    <RANKING order="2" place="-1" resultid="4232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1326" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2520" />
                    <RANKING order="2" place="2" resultid="5436" />
                    <RANKING order="3" place="3" resultid="4474" />
                    <RANKING order="4" place="4" resultid="4087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4465" />
                    <RANKING order="2" place="2" resultid="3664" />
                    <RANKING order="3" place="3" resultid="2872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1328" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1329" agemax="69" agemin="65" name="I: 65 - 69 lat" />
                <AGEGROUP agegroupid="1330" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1331" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1332" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1333" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1334" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1335" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7561" daytime="12:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7562" daytime="12:59" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7563" daytime="13:03" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1336" daytime="13:07" gender="M" number="17" order="20" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1337" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2602" />
                    <RANKING order="2" place="2" resultid="7229" />
                    <RANKING order="3" place="3" resultid="4867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1338" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5107" />
                    <RANKING order="2" place="2" resultid="3479" />
                    <RANKING order="3" place="3" resultid="2764" />
                    <RANKING order="4" place="-1" resultid="3534" />
                    <RANKING order="5" place="-1" resultid="4225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1339" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2557" />
                    <RANKING order="2" place="2" resultid="2819" />
                    <RANKING order="3" place="-1" resultid="5901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1340" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3209" />
                    <RANKING order="2" place="2" resultid="5144" />
                    <RANKING order="3" place="3" resultid="5869" />
                    <RANKING order="4" place="4" resultid="4842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1341" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4390" />
                    <RANKING order="2" place="2" resultid="4607" />
                    <RANKING order="3" place="3" resultid="4756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1342" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4076" />
                    <RANKING order="2" place="2" resultid="4345" />
                    <RANKING order="3" place="3" resultid="3887" />
                    <RANKING order="4" place="4" resultid="4994" />
                    <RANKING order="5" place="-1" resultid="2375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6233" />
                    <RANKING order="2" place="2" resultid="4833" />
                    <RANKING order="3" place="3" resultid="2574" />
                    <RANKING order="4" place="4" resultid="5444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5536" />
                    <RANKING order="2" place="2" resultid="3135" />
                    <RANKING order="3" place="3" resultid="4692" />
                    <RANKING order="4" place="4" resultid="2678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4631" />
                    <RANKING order="2" place="2" resultid="5931" />
                    <RANKING order="3" place="3" resultid="3647" />
                    <RANKING order="4" place="4" resultid="5754" />
                    <RANKING order="5" place="5" resultid="3605" />
                    <RANKING order="6" place="-1" resultid="3380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2407" />
                    <RANKING order="2" place="2" resultid="5494" />
                    <RANKING order="3" place="3" resultid="4483" />
                    <RANKING order="4" place="4" resultid="4210" />
                    <RANKING order="5" place="-1" resultid="7937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3614" />
                    <RANKING order="2" place="2" resultid="4249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1349" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1350" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1351" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1352" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7564" daytime="12:47" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7565" daytime="13:07" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7566" daytime="13:13" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7567" daytime="13:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7568" daytime="13:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7569" daytime="13:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7570" daytime="13:29" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7571" daytime="13:32" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1370" daytime="13:36" gender="F" number="18" order="22" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2324" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5201" />
                    <RANKING order="2" place="-1" resultid="2773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2325" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5200" />
                    <RANKING order="2" place="2" resultid="4350" />
                    <RANKING order="3" place="3" resultid="3779" />
                    <RANKING order="4" place="4" resultid="6393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2326" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5545" />
                    <RANKING order="2" place="2" resultid="5622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2327" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4580" />
                    <RANKING order="2" place="2" resultid="6280" />
                    <RANKING order="3" place="-1" resultid="5722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2328" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2329" agemax="319" agemin="280" name="F: 280 - 319 lat " calculate="TOTAL" />
                <AGEGROUP agegroupid="2330" agemax="359" agemin="320" name="G: 320 - 359 lat " calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7572" daytime="13:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7573" daytime="13:39" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1377" daytime="13:42" gender="M" number="19" order="23" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2331" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5203" />
                    <RANKING order="2" place="2" resultid="5720" />
                    <RANKING order="3" place="3" resultid="2775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2332" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2990" />
                    <RANKING order="2" place="2" resultid="2616" />
                    <RANKING order="3" place="3" resultid="6395" />
                    <RANKING order="4" place="4" resultid="2777" />
                    <RANKING order="5" place="5" resultid="2991" />
                    <RANKING order="6" place="6" resultid="3254" />
                    <RANKING order="7" place="7" resultid="2992" />
                    <RANKING order="8" place="8" resultid="5991" />
                    <RANKING order="9" place="9" resultid="2993" />
                    <RANKING order="10" place="10" resultid="4352" />
                    <RANKING order="11" place="-1" resultid="6397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2333" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5205" />
                    <RANKING order="2" place="2" resultid="4872" />
                    <RANKING order="3" place="3" resultid="4353" />
                    <RANKING order="4" place="4" resultid="3851" />
                    <RANKING order="5" place="5" resultid="5989" />
                    <RANKING order="6" place="6" resultid="5625" />
                    <RANKING order="7" place="7" resultid="3784" />
                    <RANKING order="8" place="8" resultid="5721" />
                    <RANKING order="9" place="9" resultid="3196" />
                    <RANKING order="10" place="10" resultid="7162" />
                    <RANKING order="11" place="11" resultid="3699" />
                    <RANKING order="12" place="-1" resultid="5397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2334" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5399" />
                    <RANKING order="2" place="2" resultid="6281" />
                    <RANKING order="3" place="3" resultid="5547" />
                    <RANKING order="4" place="4" resultid="5840" />
                    <RANKING order="5" place="5" resultid="2615" />
                    <RANKING order="6" place="6" resultid="4873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2335" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4653" />
                    <RANKING order="2" place="2" resultid="4767" />
                    <RANKING order="3" place="3" resultid="5549" />
                    <RANKING order="4" place="4" resultid="4582" />
                    <RANKING order="5" place="5" resultid="3652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2336" agemax="319" agemin="280" name="F: 280 - 319 lat " calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5986" />
                    <RANKING order="2" place="-1" resultid="3421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2337" agemax="359" agemin="320" name="G: 320 - 359 lat " calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7928" daytime="13:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7929" daytime="13:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7930" daytime="13:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7931" daytime="13:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7932" daytime="13:57" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7933" daytime="13:59" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7934" daytime="14:02" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2014-11-15" daytime="16:15" name="III Blok (Sobota)" number="3" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="1385" daytime="16:15" gender="F" number="20" order="22" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1386" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7255" />
                    <RANKING order="2" place="2" resultid="2665" />
                    <RANKING order="3" place="3" resultid="5175" />
                    <RANKING order="4" place="-1" resultid="5855" />
                    <RANKING order="5" place="-1" resultid="6473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1387" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5070" />
                    <RANKING order="2" place="2" resultid="3930" />
                    <RANKING order="3" place="3" resultid="5973" />
                    <RANKING order="4" place="4" resultid="2718" />
                    <RANKING order="5" place="5" resultid="5161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1388" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5924" />
                    <RANKING order="2" place="2" resultid="4147" />
                    <RANKING order="3" place="3" resultid="4115" />
                    <RANKING order="4" place="4" resultid="4334" />
                    <RANKING order="5" place="5" resultid="6127" />
                    <RANKING order="6" place="6" resultid="6040" />
                    <RANKING order="7" place="7" resultid="6373" />
                    <RANKING order="8" place="-1" resultid="5698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1389" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3711" />
                    <RANKING order="2" place="2" resultid="5918" />
                    <RANKING order="3" place="2" resultid="7072" />
                    <RANKING order="4" place="4" resultid="3911" />
                    <RANKING order="5" place="5" resultid="3659" />
                    <RANKING order="6" place="6" resultid="4041" />
                    <RANKING order="7" place="-1" resultid="5421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1390" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4715" />
                    <RANKING order="2" place="2" resultid="5128" />
                    <RANKING order="3" place="3" resultid="5810" />
                    <RANKING order="4" place="4" resultid="5583" />
                    <RANKING order="5" place="-1" resultid="5606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4398" />
                    <RANKING order="2" place="2" resultid="3842" />
                    <RANKING order="3" place="3" resultid="3500" />
                    <RANKING order="4" place="4" resultid="4852" />
                    <RANKING order="5" place="5" resultid="3813" />
                    <RANKING order="6" place="6" resultid="6047" />
                    <RANKING order="7" place="7" resultid="3895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1392" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4910" />
                    <RANKING order="2" place="2" resultid="5487" />
                    <RANKING order="3" place="3" resultid="5095" />
                    <RANKING order="4" place="4" resultid="6093" />
                    <RANKING order="5" place="5" resultid="2516" />
                    <RANKING order="6" place="6" resultid="5386" />
                    <RANKING order="7" place="-1" resultid="5600" />
                    <RANKING order="8" place="-1" resultid="5666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1393" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4542" />
                    <RANKING order="2" place="2" resultid="4897" />
                    <RANKING order="3" place="3" resultid="3665" />
                    <RANKING order="4" place="4" resultid="2569" />
                    <RANKING order="5" place="5" resultid="2873" />
                    <RANKING order="6" place="-1" resultid="3674" />
                    <RANKING order="7" place="-1" resultid="6078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1394" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4038" />
                    <RANKING order="2" place="2" resultid="3407" />
                    <RANKING order="3" place="3" resultid="4699" />
                    <RANKING order="4" place="4" resultid="4017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1395" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5349" />
                    <RANKING order="2" place="2" resultid="3556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1396" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4737" />
                    <RANKING order="2" place="2" resultid="3569" />
                    <RANKING order="3" place="3" resultid="3550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3485" />
                    <RANKING order="2" place="2" resultid="3919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1399" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1400" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1401" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7581" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7582" daytime="16:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7583" daytime="16:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7584" daytime="16:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7585" daytime="16:27" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7586" daytime="16:29" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7587" daytime="16:32" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7588" daytime="16:34" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7589" daytime="16:36" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7590" daytime="16:38" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7591" daytime="16:40" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1402" daytime="16:42" gender="M" number="21" order="23" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1403" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6341" />
                    <RANKING order="2" place="2" resultid="7230" />
                    <RANKING order="3" place="3" resultid="7201" />
                    <RANKING order="4" place="4" resultid="4242" />
                    <RANKING order="5" place="5" resultid="2640" />
                    <RANKING order="6" place="-1" resultid="6487" />
                    <RANKING order="7" place="-1" resultid="7154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1404" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4383" />
                    <RANKING order="2" place="2" resultid="5690" />
                    <RANKING order="3" place="3" resultid="5181" />
                    <RANKING order="4" place="4" resultid="2791" />
                    <RANKING order="5" place="5" resultid="4615" />
                    <RANKING order="6" place="6" resultid="5169" />
                    <RANKING order="7" place="7" resultid="5154" />
                    <RANKING order="8" place="8" resultid="2749" />
                    <RANKING order="9" place="9" resultid="2753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1405" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7959" />
                    <RANKING order="2" place="2" resultid="2798" />
                    <RANKING order="3" place="3" resultid="5694" />
                    <RANKING order="4" place="4" resultid="4328" />
                    <RANKING order="5" place="5" resultid="5065" />
                    <RANKING order="6" place="6" resultid="2908" />
                    <RANKING order="7" place="7" resultid="3963" />
                    <RANKING order="8" place="8" resultid="5030" />
                    <RANKING order="9" place="9" resultid="2743" />
                    <RANKING order="10" place="10" resultid="5911" />
                    <RANKING order="11" place="11" resultid="2898" />
                    <RANKING order="12" place="12" resultid="3243" />
                    <RANKING order="13" place="13" resultid="3248" />
                    <RANKING order="14" place="14" resultid="2891" />
                    <RANKING order="15" place="15" resultid="6329" />
                    <RANKING order="16" place="16" resultid="2758" />
                    <RANKING order="17" place="17" resultid="2939" />
                    <RANKING order="18" place="-1" resultid="2956" />
                    <RANKING order="19" place="-1" resultid="6453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1406" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5982" />
                    <RANKING order="2" place="2" resultid="5518" />
                    <RANKING order="3" place="3" resultid="5301" />
                    <RANKING order="4" place="4" resultid="4941" />
                    <RANKING order="5" place="5" resultid="4843" />
                    <RANKING order="6" place="6" resultid="5150" />
                    <RANKING order="7" place="7" resultid="3968" />
                    <RANKING order="8" place="-1" resultid="6422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1407" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3033" />
                    <RANKING order="2" place="2" resultid="4608" />
                    <RANKING order="3" place="3" resultid="3744" />
                    <RANKING order="4" place="4" resultid="3756" />
                    <RANKING order="5" place="5" resultid="2880" />
                    <RANKING order="6" place="6" resultid="6122" />
                    <RANKING order="7" place="7" resultid="3186" />
                    <RANKING order="8" place="8" resultid="3226" />
                    <RANKING order="9" place="9" resultid="3817" />
                    <RANKING order="10" place="10" resultid="5611" />
                    <RANKING order="11" place="11" resultid="5769" />
                    <RANKING order="12" place="12" resultid="3903" />
                    <RANKING order="13" place="13" resultid="5713" />
                    <RANKING order="14" place="-1" resultid="2810" />
                    <RANKING order="15" place="-1" resultid="5617" />
                    <RANKING order="16" place="-1" resultid="7315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1408" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3826" />
                    <RANKING order="2" place="2" resultid="3493" />
                    <RANKING order="3" place="3" resultid="4933" />
                    <RANKING order="4" place="4" resultid="3973" />
                    <RANKING order="5" place="5" resultid="6260" />
                    <RANKING order="6" place="6" resultid="5499" />
                    <RANKING order="7" place="7" resultid="6254" />
                    <RANKING order="8" place="8" resultid="3580" />
                    <RANKING order="9" place="9" resultid="4995" />
                    <RANKING order="10" place="10" resultid="4517" />
                    <RANKING order="11" place="11" resultid="4677" />
                    <RANKING order="12" place="12" resultid="4556" />
                    <RANKING order="13" place="-1" resultid="2492" />
                    <RANKING order="14" place="-1" resultid="3220" />
                    <RANKING order="15" place="-1" resultid="4106" />
                    <RANKING order="16" place="-1" resultid="5101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1409" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5377" />
                    <RANKING order="2" place="2" resultid="3059" />
                    <RANKING order="3" place="3" resultid="2611" />
                    <RANKING order="4" place="4" resultid="6241" />
                    <RANKING order="5" place="5" resultid="4407" />
                    <RANKING order="6" place="-1" resultid="3682" />
                    <RANKING order="7" place="-1" resultid="4561" />
                    <RANKING order="8" place="-1" resultid="5340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5780" />
                    <RANKING order="2" place="2" resultid="5337" />
                    <RANKING order="3" place="3" resultid="2866" />
                    <RANKING order="4" place="4" resultid="3136" />
                    <RANKING order="5" place="5" resultid="6222" />
                    <RANKING order="6" place="6" resultid="7060" />
                    <RANKING order="7" place="7" resultid="5454" />
                    <RANKING order="8" place="8" resultid="4652" />
                    <RANKING order="9" place="9" resultid="2553" />
                    <RANKING order="10" place="10" resultid="5256" />
                    <RANKING order="11" place="-1" resultid="4452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5309" />
                    <RANKING order="2" place="2" resultid="3370" />
                    <RANKING order="3" place="3" resultid="3460" />
                    <RANKING order="4" place="4" resultid="4632" />
                    <RANKING order="5" place="5" resultid="2692" />
                    <RANKING order="6" place="6" resultid="5932" />
                    <RANKING order="7" place="7" resultid="3606" />
                    <RANKING order="8" place="8" resultid="3863" />
                    <RANKING order="9" place="-1" resultid="6111" />
                    <RANKING order="10" place="-1" resultid="3381" />
                    <RANKING order="11" place="-1" resultid="3398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1412" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5426" />
                    <RANKING order="2" place="2" resultid="5466" />
                    <RANKING order="3" place="3" resultid="5877" />
                    <RANKING order="4" place="4" resultid="4446" />
                    <RANKING order="5" place="5" resultid="3596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4732" />
                    <RANKING order="2" place="2" resultid="4026" />
                    <RANKING order="3" place="-1" resultid="3631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3415" />
                    <RANKING order="2" place="2" resultid="4980" />
                    <RANKING order="3" place="3" resultid="5797" />
                    <RANKING order="4" place="-1" resultid="5889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1415" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1417" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1418" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7592" daytime="16:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7593" daytime="16:43" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7594" daytime="16:47" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7595" daytime="16:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7596" daytime="16:53" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7597" daytime="16:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7598" daytime="16:57" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7599" daytime="16:59" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7600" daytime="17:01" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7601" daytime="17:03" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7602" daytime="17:05" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7603" daytime="17:07" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7604" daytime="17:09" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7605" daytime="17:11" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7606" daytime="17:13" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7607" daytime="17:14" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7608" daytime="17:16" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7609" daytime="17:18" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7610" daytime="17:20" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7611" daytime="17:21" number="20" order="20" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1419" daytime="17:23" gender="F" number="22" order="24" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1420" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7256" />
                    <RANKING order="2" place="2" resultid="3950" />
                    <RANKING order="3" place="3" resultid="7328" />
                    <RANKING order="4" place="4" resultid="6448" />
                    <RANKING order="5" place="-1" resultid="7321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1421" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2364" />
                    <RANKING order="2" place="2" resultid="5816" />
                    <RANKING order="3" place="3" resultid="4259" />
                    <RANKING order="4" place="4" resultid="5974" />
                    <RANKING order="5" place="5" resultid="3931" />
                    <RANKING order="6" place="6" resultid="3253" />
                    <RANKING order="7" place="7" resultid="2719" />
                    <RANKING order="8" place="8" resultid="2707" />
                    <RANKING order="9" place="9" resultid="4988" />
                    <RANKING order="10" place="10" resultid="2802" />
                    <RANKING order="11" place="11" resultid="5053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1422" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4950" />
                    <RANKING order="2" place="2" resultid="3152" />
                    <RANKING order="3" place="3" resultid="5925" />
                    <RANKING order="4" place="4" resultid="4288" />
                    <RANKING order="5" place="5" resultid="6388" />
                    <RANKING order="6" place="6" resultid="6128" />
                    <RANKING order="7" place="7" resultid="5531" />
                    <RANKING order="8" place="8" resultid="6041" />
                    <RANKING order="9" place="9" resultid="4435" />
                    <RANKING order="10" place="-1" resultid="2825" />
                    <RANKING order="11" place="-1" resultid="5699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1423" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3719" />
                    <RANKING order="2" place="2" resultid="5919" />
                    <RANKING order="3" place="3" resultid="4521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1424" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5748" />
                    <RANKING order="2" place="2" resultid="5512" />
                    <RANKING order="3" place="3" resultid="4414" />
                    <RANKING order="4" place="4" resultid="5129" />
                    <RANKING order="5" place="5" resultid="4429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4399" />
                    <RANKING order="2" place="2" resultid="4536" />
                    <RANKING order="3" place="3" resultid="4853" />
                    <RANKING order="4" place="-1" resultid="4233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5437" />
                    <RANKING order="2" place="2" resultid="2518" />
                    <RANKING order="3" place="3" resultid="4475" />
                    <RANKING order="4" place="-1" resultid="5344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6190" />
                    <RANKING order="2" place="2" resultid="4898" />
                    <RANKING order="3" place="3" resultid="2860" />
                    <RANKING order="4" place="4" resultid="4466" />
                    <RANKING order="5" place="5" resultid="3666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3408" />
                    <RANKING order="2" place="2" resultid="4904" />
                    <RANKING order="3" place="3" resultid="5459" />
                    <RANKING order="4" place="4" resultid="4441" />
                    <RANKING order="5" place="5" resultid="3542" />
                    <RANKING order="6" place="6" resultid="3981" />
                    <RANKING order="7" place="-1" resultid="3389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4493" />
                    <RANKING order="2" place="2" resultid="3557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1431" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1432" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1433" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1434" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1435" agemax="-1" agemin="95" name="O: 95 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5677" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7612" daytime="17:23" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7613" daytime="17:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7614" daytime="17:27" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7615" daytime="17:29" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7616" daytime="17:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7617" daytime="17:31" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7618" daytime="17:32" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7619" daytime="17:33" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7620" daytime="17:34" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7621" daytime="17:36" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1436" daytime="17:37" gender="M" number="23" order="25" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1437" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7185" />
                    <RANKING order="2" place="2" resultid="2507" />
                    <RANKING order="3" place="3" resultid="5660" />
                    <RANKING order="4" place="4" resultid="6357" />
                    <RANKING order="5" place="5" resultid="7231" />
                    <RANKING order="6" place="6" resultid="7065" />
                    <RANKING order="7" place="7" resultid="6167" />
                    <RANKING order="8" place="-1" resultid="6489" />
                    <RANKING order="9" place="-1" resultid="7202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1438" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7224" />
                    <RANKING order="2" place="2" resultid="6429" />
                    <RANKING order="3" place="3" resultid="5672" />
                    <RANKING order="4" place="4" resultid="6160" />
                    <RANKING order="5" place="5" resultid="5108" />
                    <RANKING order="6" place="6" resultid="4384" />
                    <RANKING order="7" place="7" resultid="4616" />
                    <RANKING order="8" place="8" resultid="6444" />
                    <RANKING order="9" place="9" resultid="5089" />
                    <RANKING order="10" place="10" resultid="5187" />
                    <RANKING order="11" place="11" resultid="2765" />
                    <RANKING order="12" place="12" resultid="4458" />
                    <RANKING order="13" place="13" resultid="5650" />
                    <RANKING order="14" place="14" resultid="5155" />
                    <RANKING order="15" place="15" resultid="5120" />
                    <RANKING order="16" place="16" resultid="3182" />
                    <RANKING order="17" place="-1" resultid="3231" />
                    <RANKING order="18" place="-1" resultid="4226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1439" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2964" />
                    <RANKING order="2" place="2" resultid="6454" />
                    <RANKING order="3" place="3" resultid="4124" />
                    <RANKING order="4" place="4" resultid="6466" />
                    <RANKING order="5" place="5" resultid="2558" />
                    <RANKING order="6" place="6" resultid="5199" />
                    <RANKING order="7" place="7" resultid="2909" />
                    <RANKING order="8" place="8" resultid="6335" />
                    <RANKING order="9" place="9" resultid="3964" />
                    <RANKING order="10" place="10" resultid="6461" />
                    <RANKING order="11" place="11" resultid="6320" />
                    <RANKING order="12" place="12" resultid="2903" />
                    <RANKING order="13" place="13" resultid="5863" />
                    <RANKING order="14" place="14" resultid="5948" />
                    <RANKING order="15" place="15" resultid="2744" />
                    <RANKING order="16" place="16" resultid="5902" />
                    <RANKING order="17" place="17" resultid="5192" />
                    <RANKING order="18" place="-1" resultid="2588" />
                    <RANKING order="19" place="-1" resultid="2971" />
                    <RANKING order="20" place="-1" resultid="4141" />
                    <RANKING order="21" place="-1" resultid="6063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1440" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3436" />
                    <RANKING order="2" place="2" resultid="6295" />
                    <RANKING order="3" place="3" resultid="6153" />
                    <RANKING order="4" place="4" resultid="6314" />
                    <RANKING order="5" place="5" resultid="4789" />
                    <RANKING order="6" place="6" resultid="4270" />
                    <RANKING order="7" place="7" resultid="5478" />
                    <RANKING order="8" place="8" resultid="6302" />
                    <RANKING order="9" place="9" resultid="2914" />
                    <RANKING order="10" place="10" resultid="5082" />
                    <RANKING order="11" place="11" resultid="5317" />
                    <RANKING order="12" place="12" resultid="4942" />
                    <RANKING order="13" place="13" resultid="2984" />
                    <RANKING order="14" place="14" resultid="3750" />
                    <RANKING order="15" place="15" resultid="2924" />
                    <RANKING order="16" place="16" resultid="5870" />
                    <RANKING order="17" place="17" resultid="6032" />
                    <RANKING order="18" place="18" resultid="2399" />
                    <RANKING order="19" place="19" resultid="5023" />
                    <RANKING order="20" place="20" resultid="4551" />
                    <RANKING order="21" place="21" resultid="3969" />
                    <RANKING order="22" place="-1" resultid="2932" />
                    <RANKING order="23" place="-1" resultid="5519" />
                    <RANKING order="24" place="-1" resultid="7130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1441" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5371" />
                    <RANKING order="2" place="2" resultid="4798" />
                    <RANKING order="3" place="3" resultid="4297" />
                    <RANKING order="4" place="4" resultid="5575" />
                    <RANKING order="5" place="5" resultid="4391" />
                    <RANKING order="6" place="6" resultid="5248" />
                    <RANKING order="7" place="7" resultid="3763" />
                    <RANKING order="8" place="8" resultid="4757" />
                    <RANKING order="9" place="9" resultid="4323" />
                    <RANKING order="10" place="10" resultid="5041" />
                    <RANKING order="11" place="11" resultid="4313" />
                    <RANKING order="12" place="12" resultid="3757" />
                    <RANKING order="13" place="13" resultid="4825" />
                    <RANKING order="14" place="14" resultid="3771" />
                    <RANKING order="15" place="15" resultid="3688" />
                    <RANKING order="16" place="16" resultid="4340" />
                    <RANKING order="17" place="17" resultid="5002" />
                    <RANKING order="18" place="-1" resultid="3745" />
                    <RANKING order="19" place="-1" resultid="3831" />
                    <RANKING order="20" place="-1" resultid="5594" />
                    <RANKING order="21" place="-1" resultid="5612" />
                    <RANKING order="22" place="-1" resultid="6307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5136" />
                    <RANKING order="2" place="2" resultid="3494" />
                    <RANKING order="3" place="3" resultid="2649" />
                    <RANKING order="4" place="4" resultid="4097" />
                    <RANKING order="5" place="5" resultid="4861" />
                    <RANKING order="6" place="6" resultid="2376" />
                    <RANKING order="7" place="7" resultid="3937" />
                    <RANKING order="8" place="8" resultid="4807" />
                    <RANKING order="9" place="9" resultid="4048" />
                    <RANKING order="10" place="10" resultid="6255" />
                    <RANKING order="11" place="11" resultid="3888" />
                    <RANKING order="12" place="12" resultid="3639" />
                    <RANKING order="13" place="13" resultid="3192" />
                    <RANKING order="14" place="-1" resultid="5333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4623" />
                    <RANKING order="2" place="2" resultid="2536" />
                    <RANKING order="3" place="3" resultid="5378" />
                    <RANKING order="4" place="4" resultid="6234" />
                    <RANKING order="5" place="5" resultid="4508" />
                    <RANKING order="6" place="6" resultid="2439" />
                    <RANKING order="7" place="7" resultid="6249" />
                    <RANKING order="8" place="8" resultid="2498" />
                    <RANKING order="9" place="9" resultid="5524" />
                    <RANKING order="10" place="10" resultid="4010" />
                    <RANKING order="11" place="-1" resultid="5445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6106" />
                    <RANKING order="2" place="2" resultid="4306" />
                    <RANKING order="3" place="3" resultid="4666" />
                    <RANKING order="4" place="4" resultid="5774" />
                    <RANKING order="5" place="5" resultid="2447" />
                    <RANKING order="6" place="6" resultid="2847" />
                    <RANKING order="7" place="7" resultid="4650" />
                    <RANKING order="8" place="8" resultid="6072" />
                    <RANKING order="9" place="9" resultid="5047" />
                    <RANKING order="10" place="10" resultid="3167" />
                    <RANKING order="11" place="-1" resultid="4693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2469" />
                    <RANKING order="2" place="2" resultid="5755" />
                    <RANKING order="3" place="3" resultid="5940" />
                    <RANKING order="4" place="4" resultid="3648" />
                    <RANKING order="5" place="5" resultid="2693" />
                    <RANKING order="6" place="6" resultid="5964" />
                    <RANKING order="7" place="7" resultid="7240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4742" />
                    <RANKING order="2" place="2" resultid="2408" />
                    <RANKING order="3" place="3" resultid="5495" />
                    <RANKING order="4" place="4" resultid="4763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6135" />
                    <RANKING order="2" place="2" resultid="4918" />
                    <RANKING order="3" place="3" resultid="4570" />
                    <RANKING order="4" place="-1" resultid="3615" />
                    <RANKING order="5" place="-1" resultid="5894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2385" />
                    <RANKING order="2" place="2" resultid="4642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3871" />
                    <RANKING order="2" place="-1" resultid="5329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1451" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1452" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7622" daytime="17:37" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7623" daytime="17:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7624" daytime="17:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7625" daytime="17:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7626" daytime="17:43" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7627" daytime="17:44" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7628" daytime="17:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7629" daytime="17:47" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7630" daytime="17:48" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7631" daytime="17:49" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7632" daytime="17:50" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7633" daytime="17:51" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7634" daytime="17:52" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7635" daytime="17:53" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7636" daytime="17:54" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7637" daytime="17:55" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7638" daytime="17:56" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7639" daytime="17:57" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7640" daytime="17:58" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7641" daytime="17:59" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="7642" daytime="18:00" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="7643" daytime="18:01" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="7644" daytime="18:02" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="7645" daytime="18:03" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="7646" daytime="18:04" number="25" order="25" status="OFFICIAL" />
                <HEAT heatid="7647" daytime="18:05" number="26" order="26" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1453" daytime="18:06" gender="F" number="24" order="26" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1454" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7218" />
                    <RANKING order="2" place="2" resultid="2701" />
                    <RANKING order="3" place="3" resultid="3882" />
                    <RANKING order="4" place="4" resultid="3951" />
                    <RANKING order="5" place="5" resultid="3521" />
                    <RANKING order="6" place="6" resultid="5176" />
                    <RANKING order="7" place="-1" resultid="7322" />
                    <RANKING order="8" place="-1" resultid="7329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1455" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2365" />
                    <RANKING order="2" place="2" resultid="7137" />
                    <RANKING order="3" place="3" resultid="4501" />
                    <RANKING order="4" place="4" resultid="4131" />
                    <RANKING order="5" place="5" resultid="2526" />
                    <RANKING order="6" place="6" resultid="2784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1456" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5355" />
                    <RANKING order="2" place="2" resultid="6172" />
                    <RANKING order="3" place="3" resultid="5014" />
                    <RANKING order="4" place="4" resultid="3162" />
                    <RANKING order="5" place="5" resultid="4289" />
                    <RANKING order="6" place="6" resultid="6144" />
                    <RANKING order="7" place="-1" resultid="2826" />
                    <RANKING order="8" place="-1" resultid="5837" />
                    <RANKING order="9" place="-1" resultid="6363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1457" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3712" />
                    <RANKING order="2" place="2" resultid="3735" />
                    <RANKING order="3" place="3" resultid="5019" />
                    <RANKING order="4" place="4" resultid="3912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1458" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5506" />
                    <RANKING order="2" place="2" resultid="3836" />
                    <RANKING order="3" place="3" resultid="4415" />
                    <RANKING order="4" place="4" resultid="6208" />
                    <RANKING order="5" place="5" resultid="3529" />
                    <RANKING order="6" place="6" resultid="3727" />
                    <RANKING order="7" place="7" resultid="4430" />
                    <RANKING order="8" place="8" resultid="5710" />
                    <RANKING order="9" place="9" resultid="7248" />
                    <RANKING order="10" place="-1" resultid="6369" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5685" />
                    <RANKING order="2" place="2" resultid="3473" />
                    <RANKING order="3" place="3" resultid="2832" />
                    <RANKING order="4" place="4" resultid="6048" />
                    <RANKING order="5" place="5" resultid="3896" />
                    <RANKING order="6" place="-1" resultid="4234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1460" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5438" />
                    <RANKING order="2" place="2" resultid="6203" />
                    <RANKING order="3" place="3" resultid="6094" />
                    <RANKING order="4" place="4" resultid="5387" />
                    <RANKING order="5" place="-1" resultid="6087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1461" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4684" />
                    <RANKING order="2" place="2" resultid="5325" />
                    <RANKING order="3" place="3" resultid="3506" />
                    <RANKING order="4" place="-1" resultid="4543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1462" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3390" />
                    <RANKING order="2" place="2" resultid="3575" />
                    <RANKING order="3" place="-1" resultid="3563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1463" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6024" />
                    <RANKING order="2" place="2" resultid="6100" />
                    <RANKING order="3" place="3" resultid="4704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1464" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4729" />
                    <RANKING order="2" place="2" resultid="5785" />
                    <RANKING order="3" place="3" resultid="2475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1466" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1468" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1469" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7648" daytime="18:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7649" daytime="18:09" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7650" daytime="18:13" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7651" daytime="18:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7652" daytime="18:17" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7653" daytime="18:19" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7654" daytime="18:21" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7655" daytime="18:23" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7656" daytime="18:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7657" daytime="18:27" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7658" daytime="18:29" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1470" daytime="18:31" gender="M" number="25" order="27" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1471" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7186" />
                    <RANKING order="2" place="2" resultid="7210" />
                    <RANKING order="3" place="3" resultid="2641" />
                    <RANKING order="4" place="-1" resultid="6480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1472" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5704" />
                    <RANKING order="2" place="2" resultid="6430" />
                    <RANKING order="3" place="3" resultid="7145" />
                    <RANKING order="4" place="4" resultid="6161" />
                    <RANKING order="5" place="5" resultid="2739" />
                    <RANKING order="6" place="6" resultid="5718" />
                    <RANKING order="7" place="-1" resultid="5090" />
                    <RANKING order="8" place="-1" resultid="6177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1473" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3028" />
                    <RANKING order="2" place="2" resultid="2564" />
                    <RANKING order="3" place="3" resultid="2589" />
                    <RANKING order="4" place="4" resultid="2957" />
                    <RANKING order="5" place="5" resultid="6348" />
                    <RANKING order="6" place="6" resultid="5912" />
                    <RANKING order="7" place="7" resultid="2979" />
                    <RANKING order="8" place="8" resultid="2947" />
                    <RANKING order="9" place="-1" resultid="2940" />
                    <RANKING order="10" place="-1" resultid="3999" />
                    <RANKING order="11" place="-1" resultid="5949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1474" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3437" />
                    <RANKING order="2" place="2" resultid="4790" />
                    <RANKING order="3" place="3" resultid="3144" />
                    <RANKING order="4" place="4" resultid="5956" />
                    <RANKING order="5" place="5" resultid="4271" />
                    <RANKING order="6" place="6" resultid="3991" />
                    <RANKING order="7" place="7" resultid="5871" />
                    <RANKING order="8" place="8" resultid="3778" />
                    <RANKING order="9" place="9" resultid="4514" />
                    <RANKING order="10" place="-1" resultid="5829" />
                    <RANKING order="11" place="-1" resultid="6154" />
                    <RANKING order="12" place="-1" resultid="6315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1475" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5618" />
                    <RANKING order="2" place="2" resultid="3179" />
                    <RANKING order="3" place="3" resultid="3832" />
                    <RANKING order="4" place="4" resultid="4826" />
                    <RANKING order="5" place="-1" resultid="3175" />
                    <RANKING order="6" place="-1" resultid="4069" />
                    <RANKING order="7" place="-1" resultid="5823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1476" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5682" />
                    <RANKING order="2" place="2" resultid="4968" />
                    <RANKING order="3" place="3" resultid="2521" />
                    <RANKING order="4" place="4" resultid="3848" />
                    <RANKING order="5" place="5" resultid="2582" />
                    <RANKING order="6" place="6" resultid="4098" />
                    <RANKING order="7" place="7" resultid="3581" />
                    <RANKING order="8" place="8" resultid="4862" />
                    <RANKING order="9" place="9" resultid="5656" />
                    <RANKING order="10" place="10" resultid="2634" />
                    <RANKING order="11" place="-1" resultid="3051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1477" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6435" />
                    <RANKING order="2" place="2" resultid="6020" />
                    <RANKING order="3" place="3" resultid="4624" />
                    <RANKING order="4" place="4" resultid="3060" />
                    <RANKING order="5" place="5" resultid="2440" />
                    <RANKING order="6" place="6" resultid="3822" />
                    <RANKING order="7" place="7" resultid="3683" />
                    <RANKING order="8" place="-1" resultid="2537" />
                    <RANKING order="9" place="-1" resultid="2612" />
                    <RANKING order="10" place="-1" resultid="4239" />
                    <RANKING order="11" place="-1" resultid="4509" />
                    <RANKING order="12" place="-1" resultid="4834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1478" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4667" />
                    <RANKING order="2" place="2" resultid="5537" />
                    <RANKING order="3" place="3" resultid="4926" />
                    <RANKING order="4" place="4" resultid="2685" />
                    <RANKING order="5" place="5" resultid="4750" />
                    <RANKING order="6" place="6" resultid="3168" />
                    <RANKING order="7" place="-1" resultid="4453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1479" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4957" />
                    <RANKING order="2" place="2" resultid="3649" />
                    <RANKING order="3" place="3" resultid="2430" />
                    <RANKING order="4" place="4" resultid="3864" />
                    <RANKING order="5" place="-1" resultid="5310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1480" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4816" />
                    <RANKING order="2" place="2" resultid="4709" />
                    <RANKING order="3" place="3" resultid="4211" />
                    <RANKING order="4" place="4" resultid="5878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4919" />
                    <RANKING order="2" place="2" resultid="5008" />
                    <RANKING order="3" place="3" resultid="5895" />
                    <RANKING order="4" place="4" resultid="4027" />
                    <RANKING order="5" place="5" resultid="3588" />
                    <RANKING order="6" place="-1" resultid="3632" />
                    <RANKING order="7" place="-1" resultid="4530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4643" />
                    <RANKING order="2" place="2" resultid="5798" />
                    <RANKING order="3" place="3" resultid="4981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1484" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1485" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1486" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7659" daytime="18:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7660" daytime="18:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7661" daytime="18:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7662" daytime="18:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7663" daytime="18:43" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7664" daytime="18:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7665" daytime="18:47" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7666" daytime="18:49" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7667" daytime="18:51" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7668" daytime="18:52" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7669" daytime="18:54" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7670" daytime="18:56" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7671" daytime="18:58" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7672" daytime="18:59" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7673" daytime="19:01" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7674" daytime="19:02" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1487" daytime="19:04" gender="F" number="26" order="28" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1488" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2666" />
                    <RANKING order="2" place="2" resultid="2702" />
                    <RANKING order="3" place="3" resultid="7219" />
                    <RANKING order="4" place="4" resultid="5077" />
                    <RANKING order="5" place="-1" resultid="6449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1489" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7138" />
                    <RANKING order="2" place="2" resultid="2529" />
                    <RANKING order="3" place="3" resultid="5071" />
                    <RANKING order="4" place="4" resultid="4220" />
                    <RANKING order="5" place="5" resultid="5588" />
                    <RANKING order="6" place="6" resultid="5162" />
                    <RANKING order="7" place="7" resultid="6385" />
                    <RANKING order="8" place="8" resultid="2785" />
                    <RANKING order="9" place="9" resultid="4989" />
                    <RANKING order="10" place="10" resultid="5054" />
                    <RANKING order="11" place="11" resultid="4083" />
                    <RANKING order="12" place="12" resultid="7943" />
                    <RANKING order="13" place="-1" resultid="2713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1490" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4951" />
                    <RANKING order="2" place="2" resultid="3153" />
                    <RANKING order="3" place="3" resultid="5356" />
                    <RANKING order="4" place="4" resultid="4335" />
                    <RANKING order="5" place="5" resultid="4436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1491" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2816" />
                    <RANKING order="2" place="2" resultid="3720" />
                    <RANKING order="3" place="3" resultid="6056" />
                    <RANKING order="4" place="4" resultid="3736" />
                    <RANKING order="5" place="5" resultid="7073" />
                    <RANKING order="6" place="6" resultid="5020" />
                    <RANKING order="7" place="7" resultid="3660" />
                    <RANKING order="8" place="8" resultid="4522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1492" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2461" />
                    <RANKING order="2" place="2" resultid="3728" />
                    <RANKING order="3" place="3" resultid="7249" />
                    <RANKING order="4" place="4" resultid="2674" />
                    <RANKING order="5" place="-1" resultid="5392" />
                    <RANKING order="6" place="-1" resultid="5607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3474" />
                    <RANKING order="2" place="2" resultid="4279" />
                    <RANKING order="3" place="3" resultid="3843" />
                    <RANKING order="4" place="4" resultid="2833" />
                    <RANKING order="5" place="5" resultid="4537" />
                    <RANKING order="6" place="-1" resultid="3810" />
                    <RANKING order="7" place="-1" resultid="5686" />
                    <RANKING order="8" place="-1" resultid="3501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6198" />
                    <RANKING order="2" place="2" resultid="5488" />
                    <RANKING order="3" place="3" resultid="4476" />
                    <RANKING order="4" place="4" resultid="5096" />
                    <RANKING order="5" place="5" resultid="5601" />
                    <RANKING order="6" place="-1" resultid="5667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1495" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6191" />
                    <RANKING order="2" place="2" resultid="4467" />
                    <RANKING order="3" place="3" resultid="2840" />
                    <RANKING order="4" place="4" resultid="2874" />
                    <RANKING order="5" place="-1" resultid="3675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1496" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4905" />
                    <RANKING order="2" place="2" resultid="5460" />
                    <RANKING order="3" place="3" resultid="3543" />
                    <RANKING order="4" place="4" resultid="4746" />
                    <RANKING order="5" place="5" resultid="3982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1497" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5061" />
                    <RANKING order="2" place="2" resultid="4494" />
                    <RANKING order="3" place="3" resultid="3621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1498" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1499" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1500" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1502" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1503" agemax="-1" agemin="95" name="O: 95 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5678" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7675" daytime="19:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7676" daytime="19:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7677" daytime="19:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7678" daytime="19:19" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7679" daytime="19:23" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7680" daytime="19:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7681" daytime="19:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7682" daytime="19:33" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7683" daytime="19:36" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7684" daytime="19:40" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7685" daytime="19:42" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1504" daytime="19:46" gender="M" number="27" order="29" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1505" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7194" />
                    <RANKING order="2" place="2" resultid="2508" />
                    <RANKING order="3" place="3" resultid="2603" />
                    <RANKING order="4" place="4" resultid="4868" />
                    <RANKING order="5" place="5" resultid="4005" />
                    <RANKING order="6" place="6" resultid="4723" />
                    <RANKING order="7" place="7" resultid="4137" />
                    <RANKING order="8" place="-1" resultid="2457" />
                    <RANKING order="9" place="-1" resultid="6342" />
                    <RANKING order="10" place="-1" resultid="7155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1506" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5673" />
                    <RANKING order="2" place="2" resultid="6178" />
                    <RANKING order="3" place="3" resultid="2792" />
                    <RANKING order="4" place="4" resultid="4459" />
                    <RANKING order="5" place="5" resultid="5121" />
                    <RANKING order="6" place="6" resultid="3232" />
                    <RANKING order="7" place="7" resultid="3183" />
                    <RANKING order="8" place="-1" resultid="4227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1507" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2965" />
                    <RANKING order="2" place="2" resultid="2726" />
                    <RANKING order="3" place="3" resultid="2546" />
                    <RANKING order="4" place="4" resultid="6467" />
                    <RANKING order="5" place="5" resultid="3958" />
                    <RANKING order="6" place="6" resultid="3879" />
                    <RANKING order="7" place="7" resultid="5193" />
                    <RANKING order="8" place="8" resultid="4319" />
                    <RANKING order="9" place="9" resultid="4974" />
                    <RANKING order="10" place="-1" resultid="2565" />
                    <RANKING order="11" place="-1" resultid="4142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1508" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5983" />
                    <RANKING order="2" place="2" resultid="3210" />
                    <RANKING order="3" place="3" resultid="5083" />
                    <RANKING order="4" place="4" resultid="3992" />
                    <RANKING order="5" place="5" resultid="4423" />
                    <RANKING order="6" place="6" resultid="2925" />
                    <RANKING order="7" place="7" resultid="2733" />
                    <RANKING order="8" place="8" resultid="4673" />
                    <RANKING order="9" place="9" resultid="4552" />
                    <RANKING order="10" place="10" resultid="6324" />
                    <RANKING order="11" place="-1" resultid="2915" />
                    <RANKING order="12" place="-1" resultid="2933" />
                    <RANKING order="13" place="-1" resultid="4094" />
                    <RANKING order="14" place="-1" resultid="5479" />
                    <RANKING order="15" place="-1" resultid="6296" />
                    <RANKING order="16" place="-1" resultid="6423" />
                    <RANKING order="17" place="-1" resultid="7131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1509" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4799" />
                    <RANKING order="2" place="2" resultid="3238" />
                    <RANKING order="3" place="3" resultid="4298" />
                    <RANKING order="4" place="4" resultid="3158" />
                    <RANKING order="5" place="5" resultid="3764" />
                    <RANKING order="6" place="6" resultid="5249" />
                    <RANKING order="7" place="7" resultid="3454" />
                    <RANKING order="8" place="8" resultid="5042" />
                    <RANKING order="9" place="9" resultid="4392" />
                    <RANKING order="10" place="10" resultid="2452" />
                    <RANKING order="11" place="11" resultid="4314" />
                    <RANKING order="12" place="12" resultid="6123" />
                    <RANKING order="13" place="13" resultid="3772" />
                    <RANKING order="14" place="14" resultid="2652" />
                    <RANKING order="15" place="15" resultid="3924" />
                    <RANKING order="16" place="16" resultid="4341" />
                    <RANKING order="17" place="17" resultid="5003" />
                    <RANKING order="18" place="18" resultid="3689" />
                    <RANKING order="19" place="-1" resultid="2811" />
                    <RANKING order="20" place="-1" resultid="4070" />
                    <RANKING order="21" place="-1" resultid="4961" />
                    <RANKING order="22" place="-1" resultid="5361" />
                    <RANKING order="23" place="-1" resultid="5714" />
                    <RANKING order="24" place="-1" resultid="6308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4077" />
                    <RANKING order="2" place="2" resultid="3043" />
                    <RANKING order="3" place="3" resultid="5137" />
                    <RANKING order="4" place="4" resultid="6266" />
                    <RANKING order="5" place="5" resultid="6261" />
                    <RANKING order="6" place="6" resultid="3938" />
                    <RANKING order="7" place="7" resultid="5764" />
                    <RANKING order="8" place="8" resultid="4934" />
                    <RANKING order="9" place="9" resultid="3849" />
                    <RANKING order="10" place="10" resultid="2658" />
                    <RANKING order="11" place="11" resultid="4808" />
                    <RANKING order="12" place="12" resultid="4346" />
                    <RANKING order="13" place="13" resultid="3640" />
                    <RANKING order="14" place="14" resultid="4518" />
                    <RANKING order="15" place="15" resultid="3193" />
                    <RANKING order="16" place="-1" resultid="2416" />
                    <RANKING order="17" place="-1" resultid="2493" />
                    <RANKING order="18" place="-1" resultid="3516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1511" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2595" />
                    <RANKING order="2" place="2" resultid="3511" />
                    <RANKING order="3" place="3" resultid="2575" />
                    <RANKING order="4" place="4" resultid="4562" />
                    <RANKING order="5" place="-1" resultid="5115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1512" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4307" />
                    <RANKING order="2" place="2" resultid="6107" />
                    <RANKING order="3" place="3" resultid="2448" />
                    <RANKING order="4" place="4" resultid="4694" />
                    <RANKING order="5" place="5" resultid="6073" />
                    <RANKING order="6" place="6" resultid="6228" />
                    <RANKING order="7" place="7" resultid="5048" />
                    <RANKING order="8" place="8" resultid="5257" />
                    <RANKING order="9" place="-1" resultid="2848" />
                    <RANKING order="10" place="-1" resultid="3944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1513" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2395" />
                    <RANKING order="2" place="2" resultid="6116" />
                    <RANKING order="3" place="3" resultid="5941" />
                    <RANKING order="4" place="4" resultid="3399" />
                    <RANKING order="5" place="5" resultid="5756" />
                    <RANKING order="6" place="6" resultid="7241" />
                    <RANKING order="7" place="-1" resultid="2431" />
                    <RANKING order="8" place="-1" resultid="6276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1514" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4484" />
                    <RANKING order="2" place="2" resultid="2856" />
                    <RANKING order="3" place="3" resultid="5883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5009" />
                    <RANKING order="2" place="2" resultid="6136" />
                    <RANKING order="3" place="3" resultid="4531" />
                    <RANKING order="4" place="4" resultid="4250" />
                    <RANKING order="5" place="-1" resultid="3626" />
                    <RANKING order="6" place="-1" resultid="4571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3872" />
                    <RANKING order="2" place="2" resultid="7180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1518" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1519" agemax="94" agemin="90" name="N: 90 - 94 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1520" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7686" daytime="19:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7687" daytime="19:51" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7688" daytime="19:57" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7689" daytime="20:01" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7690" daytime="20:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7691" daytime="20:09" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7692" daytime="20:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7693" daytime="20:16" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7694" daytime="20:19" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7695" daytime="20:22" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7696" daytime="20:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7697" daytime="20:28" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7698" daytime="20:31" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7699" daytime="20:34" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7700" daytime="20:37" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7701" daytime="20:40" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7702" daytime="20:43" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7703" daytime="20:46" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7704" daytime="20:48" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7705" daytime="20:51" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="7706" daytime="20:54" number="21" order="21" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1521" daytime="20:56" gender="F" number="28" order="31" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2338" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2339" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5202" />
                    <RANKING order="2" place="2" resultid="4351" />
                    <RANKING order="3" place="3" resultid="3780" />
                    <RANKING order="4" place="4" resultid="6394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2340" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4578" />
                    <RANKING order="2" place="2" resultid="5546" />
                    <RANKING order="3" place="3" resultid="5621" />
                    <RANKING order="4" place="-1" resultid="5401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2341" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6284" />
                    <RANKING order="2" place="2" resultid="4579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2342" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2343" agemax="319" agemin="280" name="F: 280 - 319 lat " calculate="TOTAL" />
                <AGEGROUP agegroupid="2344" agemax="359" agemin="320" name="G: 320 - 359 lat " calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7707" daytime="20:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7708" daytime="21:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1528" daytime="21:03" gender="M" number="29" order="32" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2345" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5204" />
                    <RANKING order="2" place="2" resultid="2776" />
                    <RANKING order="3" place="3" resultid="7997" />
                    <RANKING order="4" place="-1" resultid="5724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2346" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3446" />
                    <RANKING order="2" place="2" resultid="2986" />
                    <RANKING order="3" place="3" resultid="6396" />
                    <RANKING order="4" place="4" resultid="2614" />
                    <RANKING order="5" place="5" resultid="5207" />
                    <RANKING order="6" place="6" resultid="4354" />
                    <RANKING order="7" place="7" resultid="2987" />
                    <RANKING order="8" place="8" resultid="3255" />
                    <RANKING order="9" place="9" resultid="2778" />
                    <RANKING order="10" place="10" resultid="5208" />
                    <RANKING order="11" place="11" resultid="2988" />
                    <RANKING order="12" place="12" resultid="2989" />
                    <RANKING order="13" place="-1" resultid="3195" />
                    <RANKING order="14" place="-1" resultid="5992" />
                    <RANKING order="15" place="-1" resultid="6462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2347" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4874" />
                    <RANKING order="2" place="2" resultid="5396" />
                    <RANKING order="3" place="3" resultid="5206" />
                    <RANKING order="4" place="4" resultid="4654" />
                    <RANKING order="5" place="5" resultid="3785" />
                    <RANKING order="6" place="6" resultid="5626" />
                    <RANKING order="7" place="7" resultid="3852" />
                    <RANKING order="8" place="8" resultid="2423" />
                    <RANKING order="9" place="9" resultid="4348" />
                    <RANKING order="10" place="10" resultid="3700" />
                    <RANKING order="11" place="-1" resultid="5723" />
                    <RANKING order="12" place="-1" resultid="5990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2348" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6282" />
                    <RANKING order="2" place="2" resultid="5548" />
                    <RANKING order="3" place="3" resultid="4875" />
                    <RANKING order="4" place="4" resultid="2617" />
                    <RANKING order="5" place="-1" resultid="5400" />
                    <RANKING order="6" place="-1" resultid="5841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2349" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4769" />
                    <RANKING order="2" place="2" resultid="4583" />
                    <RANKING order="3" place="3" resultid="5550" />
                    <RANKING order="4" place="-1" resultid="3420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2350" agemax="319" agemin="280" name="F: 280 - 319 lat " calculate="TOTAL" />
                <AGEGROUP agegroupid="2351" agemax="359" agemin="320" name="G: 320 - 359 lat " calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7709" daytime="21:03" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7710" daytime="21:07" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7711" daytime="21:11" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7712" daytime="21:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7713" daytime="21:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7714" daytime="21:19" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7715" daytime="21:21" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7716" daytime="21:24" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1542" daytime="21:26" gender="F" number="30" order="34" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1543" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3522" />
                    <RANKING order="2" place="2" resultid="5856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1544" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5817" />
                    <RANKING order="2" place="2" resultid="4260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1545" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4116" />
                    <RANKING order="2" place="2" resultid="6145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1546" agemax="39" agemin="35" name="C: 35 - 39 lat" />
                <AGEGROUP agegroupid="1547" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1548" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1549" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4911" />
                    <RANKING order="2" place="2" resultid="4088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1550" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1551" agemax="64" agemin="60" name="H: 60 - 64 lat" />
                <AGEGROUP agegroupid="1552" agemax="69" agemin="65" name="I: 65 - 69 lat" />
                <AGEGROUP agegroupid="1553" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1554" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1555" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1556" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1557" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1558" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7717" daytime="21:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7718" daytime="21:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1559" daytime="21:42" gender="M" number="31" order="35" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1560" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2604" />
                    <RANKING order="2" place="2" resultid="4869" />
                    <RANKING order="3" place="3" resultid="7211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1561" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7146" />
                    <RANKING order="2" place="2" resultid="3480" />
                    <RANKING order="3" place="3" resultid="6184" />
                    <RANKING order="4" place="-1" resultid="2766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1562" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4628" />
                    <RANKING order="2" place="2" resultid="2547" />
                    <RANKING order="3" place="3" resultid="8003" />
                    <RANKING order="4" place="4" resultid="4329" />
                    <RANKING order="5" place="-1" resultid="2948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1563" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3211" />
                    <RANKING order="2" place="2" resultid="5145" />
                    <RANKING order="3" place="3" resultid="4844" />
                    <RANKING order="4" place="4" resultid="5318" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1564" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3034" />
                    <RANKING order="2" place="2" resultid="8002" />
                    <RANKING order="3" place="-1" resultid="3904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1565" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3044" />
                    <RANKING order="2" place="2" resultid="2523" />
                    <RANKING order="3" place="3" resultid="7984" />
                    <RANKING order="4" place="4" resultid="4107" />
                    <RANKING order="5" place="5" resultid="4049" />
                    <RANKING order="6" place="6" resultid="4996" />
                    <RANKING order="7" place="-1" resultid="3889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1566" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6235" />
                    <RANKING order="2" place="2" resultid="4835" />
                    <RANKING order="3" place="3" resultid="2499" />
                    <RANKING order="4" place="4" resultid="7987" />
                    <RANKING order="5" place="5" resultid="2576" />
                    <RANKING order="6" place="6" resultid="5446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1567" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5538" />
                    <RANKING order="2" place="2" resultid="2867" />
                    <RANKING order="3" place="3" resultid="3137" />
                    <RANKING order="4" place="4" resultid="4927" />
                    <RANKING order="5" place="5" resultid="2679" />
                    <RANKING order="6" place="-1" resultid="2686" />
                    <RANKING order="7" place="-1" resultid="5781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1568" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4633" />
                    <RANKING order="2" place="2" resultid="5933" />
                    <RANKING order="3" place="3" resultid="5965" />
                    <RANKING order="4" place="4" resultid="3607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1569" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4817" />
                    <RANKING order="2" place="2" resultid="2409" />
                    <RANKING order="3" place="3" resultid="4485" />
                    <RANKING order="4" place="4" resultid="4212" />
                    <RANKING order="5" place="5" resultid="3597" />
                    <RANKING order="6" place="-1" resultid="5884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3616" />
                    <RANKING order="2" place="2" resultid="4251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1571" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1572" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1573" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1574" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1575" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7974" daytime="21:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7975" daytime="21:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7976" daytime="22:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7977" daytime="22:11" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7978" daytime="22:19" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7979" daytime="22:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7980" daytime="22:33" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7981" daytime="22:39" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7982" daytime="22:46" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7983" daytime="22:52" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2014-11-16" daytime="09:00" name="IV Blok (Niedziela)" number="4" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1577" daytime="09:00" gender="F" number="32" order="36" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1578" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3952" />
                    <RANKING order="2" place="2" resultid="3523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1579" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5975" />
                    <RANKING order="2" place="2" resultid="4261" />
                    <RANKING order="3" place="3" resultid="5163" />
                    <RANKING order="4" place="4" resultid="4990" />
                    <RANKING order="5" place="-1" resultid="5055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1580" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4952" />
                    <RANKING order="2" place="2" resultid="3154" />
                    <RANKING order="3" place="3" resultid="5926" />
                    <RANKING order="4" place="4" resultid="4117" />
                    <RANKING order="5" place="5" resultid="4290" />
                    <RANKING order="6" place="6" resultid="4283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1581" agemax="39" agemin="35" name="C: 35 - 39 lat" />
                <AGEGROUP agegroupid="1582" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5513" />
                    <RANKING order="2" place="2" resultid="2462" />
                    <RANKING order="3" place="3" resultid="4431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4538" />
                    <RANKING order="2" place="2" resultid="4854" />
                    <RANKING order="3" place="-1" resultid="4235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1584" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4912" />
                    <RANKING order="2" place="2" resultid="5439" />
                    <RANKING order="3" place="3" resultid="2519" />
                    <RANKING order="4" place="4" resultid="4477" />
                    <RANKING order="5" place="5" resultid="4089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6192" />
                    <RANKING order="2" place="2" resultid="4468" />
                    <RANKING order="3" place="3" resultid="3667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1586" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3409" />
                    <RANKING order="2" place="2" resultid="3544" />
                    <RANKING order="3" place="3" resultid="3391" />
                    <RANKING order="4" place="-1" resultid="5461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1587" agemax="69" agemin="65" name="I: 65 - 69 lat" />
                <AGEGROUP agegroupid="1588" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1589" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1590" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1591" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1592" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1593" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7730" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7731" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7732" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7733" daytime="09:07" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7734" daytime="09:09" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7735" daytime="09:11" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1594" daytime="09:13" gender="M" number="33" order="37" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1595" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2509" />
                    <RANKING order="2" place="2" resultid="2605" />
                    <RANKING order="3" place="3" resultid="6343" />
                    <RANKING order="4" place="4" resultid="6358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1596" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5791" />
                    <RANKING order="2" place="2" resultid="2767" />
                    <RANKING order="3" place="3" resultid="4460" />
                    <RANKING order="4" place="4" resultid="5170" />
                    <RANKING order="5" place="-1" resultid="3481" />
                    <RANKING order="6" place="-1" resultid="4228" />
                    <RANKING order="7" place="-1" resultid="5156" />
                    <RANKING order="8" place="-1" resultid="5719" />
                    <RANKING order="9" place="-1" resultid="6162" />
                    <RANKING order="10" place="-1" resultid="5110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1597" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2966" />
                    <RANKING order="2" place="2" resultid="4125" />
                    <RANKING order="3" place="3" resultid="2559" />
                    <RANKING order="4" place="4" resultid="5032" />
                    <RANKING order="5" place="5" resultid="2590" />
                    <RANKING order="6" place="6" resultid="2548" />
                    <RANKING order="7" place="7" resultid="5950" />
                    <RANKING order="8" place="8" resultid="5864" />
                    <RANKING order="9" place="-1" resultid="2949" />
                    <RANKING order="10" place="-1" resultid="4143" />
                    <RANKING order="11" place="-1" resultid="5904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3438" />
                    <RANKING order="2" place="2" resultid="3212" />
                    <RANKING order="3" place="3" resultid="2916" />
                    <RANKING order="4" place="3" resultid="5831" />
                    <RANKING order="5" place="5" resultid="5146" />
                    <RANKING order="6" place="6" resultid="5084" />
                    <RANKING order="7" place="7" resultid="5319" />
                    <RANKING order="8" place="8" resultid="2926" />
                    <RANKING order="9" place="9" resultid="6033" />
                    <RANKING order="10" place="-1" resultid="3751" />
                    <RANKING order="11" place="-1" resultid="4272" />
                    <RANKING order="12" place="-1" resultid="5480" />
                    <RANKING order="13" place="-1" resultid="5958" />
                    <RANKING order="14" place="-1" resultid="6155" />
                    <RANKING order="15" place="-1" resultid="6297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4800" />
                    <RANKING order="2" place="2" resultid="4299" />
                    <RANKING order="3" place="3" resultid="5250" />
                    <RANKING order="4" place="4" resultid="5577" />
                    <RANKING order="5" place="5" resultid="3159" />
                    <RANKING order="6" place="6" resultid="3833" />
                    <RANKING order="7" place="7" resultid="3765" />
                    <RANKING order="8" place="8" resultid="4758" />
                    <RANKING order="9" place="9" resultid="4827" />
                    <RANKING order="10" place="-1" resultid="3905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3495" />
                    <RANKING order="2" place="2" resultid="4078" />
                    <RANKING order="3" place="3" resultid="2378" />
                    <RANKING order="4" place="4" resultid="4935" />
                    <RANKING order="5" place="5" resultid="6262" />
                    <RANKING order="6" place="6" resultid="4863" />
                    <RANKING order="7" place="7" resultid="4050" />
                    <RANKING order="8" place="8" resultid="4347" />
                    <RANKING order="9" place="9" resultid="3641" />
                    <RANKING order="10" place="10" resultid="4809" />
                    <RANKING order="11" place="11" resultid="4997" />
                    <RANKING order="12" place="-1" resultid="3194" />
                    <RANKING order="13" place="-1" resultid="3890" />
                    <RANKING order="14" place="-1" resultid="5138" />
                    <RANKING order="15" place="-1" resultid="5334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6236" />
                    <RANKING order="2" place="2" resultid="2538" />
                    <RANKING order="3" place="3" resultid="4836" />
                    <RANKING order="4" place="4" resultid="2577" />
                    <RANKING order="5" place="-1" resultid="2596" />
                    <RANKING order="6" place="-1" resultid="4012" />
                    <RANKING order="7" place="-1" resultid="5447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4308" />
                    <RANKING order="2" place="2" resultid="6108" />
                    <RANKING order="3" place="3" resultid="5775" />
                    <RANKING order="4" place="4" resultid="3138" />
                    <RANKING order="5" place="5" resultid="3169" />
                    <RANKING order="6" place="-1" resultid="2849" />
                    <RANKING order="7" place="-1" resultid="5539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5757" />
                    <RANKING order="2" place="2" resultid="3650" />
                    <RANKING order="3" place="3" resultid="5942" />
                    <RANKING order="4" place="4" resultid="2694" />
                    <RANKING order="5" place="5" resultid="5966" />
                    <RANKING order="6" place="-1" resultid="2470" />
                    <RANKING order="7" place="-1" resultid="3383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2410" />
                    <RANKING order="2" place="2" resultid="4486" />
                    <RANKING order="3" place="3" resultid="4213" />
                    <RANKING order="4" place="-1" resultid="5496" />
                    <RANKING order="5" place="-1" resultid="5885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6137" />
                    <RANKING order="2" place="2" resultid="3617" />
                    <RANKING order="3" place="-1" resultid="4252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1606" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3416" />
                    <RANKING order="2" place="-1" resultid="2387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1607" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1608" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1609" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1610" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7736" daytime="09:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7737" daytime="09:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7738" daytime="09:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7739" daytime="09:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7740" daytime="09:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7741" daytime="09:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7742" daytime="09:28" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7743" daytime="09:30" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7744" daytime="09:32" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7745" daytime="09:34" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7746" daytime="09:36" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7747" daytime="09:37" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7748" daytime="09:39" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7749" daytime="09:41" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7750" daytime="09:42" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7751" daytime="09:44" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7752" daytime="09:46" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1611" daytime="09:47" gender="F" number="34" order="38" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1612" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7220" />
                    <RANKING order="2" place="2" resultid="3524" />
                    <RANKING order="3" place="3" resultid="5857" />
                    <RANKING order="4" place="4" resultid="7330" />
                    <RANKING order="5" place="-1" resultid="3883" />
                    <RANKING order="6" place="-1" resultid="7323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1613" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2366" />
                    <RANKING order="2" place="2" resultid="4502" />
                    <RANKING order="3" place="3" resultid="4132" />
                    <RANKING order="4" place="4" resultid="7139" />
                    <RANKING order="5" place="5" resultid="2527" />
                    <RANKING order="6" place="6" resultid="2786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1614" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5357" />
                    <RANKING order="2" place="2" resultid="6173" />
                    <RANKING order="3" place="3" resultid="4291" />
                    <RANKING order="4" place="-1" resultid="5838" />
                    <RANKING order="5" place="-1" resultid="6146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1615" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3713" />
                    <RANKING order="2" place="2" resultid="3737" />
                    <RANKING order="3" place="-1" resultid="6058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1616" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5507" />
                    <RANKING order="2" place="2" resultid="3837" />
                    <RANKING order="3" place="3" resultid="3530" />
                    <RANKING order="4" place="4" resultid="3729" />
                    <RANKING order="5" place="5" resultid="6209" />
                    <RANKING order="6" place="6" resultid="4432" />
                    <RANKING order="7" place="-1" resultid="7250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1617" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3475" />
                    <RANKING order="2" place="2" resultid="5687" />
                    <RANKING order="3" place="3" resultid="2834" />
                    <RANKING order="4" place="4" resultid="3897" />
                    <RANKING order="5" place="-1" resultid="4236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6095" />
                    <RANKING order="2" place="2" resultid="5440" />
                    <RANKING order="3" place="3" resultid="6088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4686" />
                    <RANKING order="2" place="2" resultid="3507" />
                    <RANKING order="3" place="3" resultid="3676" />
                    <RANKING order="4" place="4" resultid="2875" />
                    <RANKING order="5" place="-1" resultid="6080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1620" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3392" />
                    <RANKING order="2" place="2" resultid="3576" />
                    <RANKING order="3" place="3" resultid="3983" />
                    <RANKING order="4" place="-1" resultid="3564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1621" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6025" />
                    <RANKING order="2" place="2" resultid="6101" />
                    <RANKING order="3" place="-1" resultid="4705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1622" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2476" />
                    <RANKING order="2" place="-1" resultid="5786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1623" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1624" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1625" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1626" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1627" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7753" daytime="09:47" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7754" daytime="09:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7755" daytime="10:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7756" daytime="10:07" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7757" daytime="10:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7758" daytime="10:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7759" daytime="10:19" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7760" daytime="10:23" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7761" daytime="10:26" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1628" daytime="10:29" gender="M" number="35" order="39" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1629" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7212" />
                    <RANKING order="2" place="2" resultid="4870" />
                    <RANKING order="3" place="-1" resultid="2642" />
                    <RANKING order="4" place="-1" resultid="6482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1630" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5705" />
                    <RANKING order="2" place="2" resultid="7147" />
                    <RANKING order="3" place="3" resultid="4419" />
                    <RANKING order="4" place="-1" resultid="5091" />
                    <RANKING order="5" place="-1" resultid="6163" />
                    <RANKING order="6" place="-1" resultid="6179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1631" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2591" />
                    <RANKING order="2" place="2" resultid="2566" />
                    <RANKING order="3" place="3" resultid="2959" />
                    <RANKING order="4" place="4" resultid="2821" />
                    <RANKING order="5" place="-1" resultid="2893" />
                    <RANKING order="6" place="-1" resultid="5913" />
                    <RANKING order="7" place="-1" resultid="6349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1632" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4791" />
                    <RANKING order="2" place="2" resultid="3145" />
                    <RANKING order="3" place="3" resultid="3993" />
                    <RANKING order="4" place="4" resultid="5832" />
                    <RANKING order="5" place="5" resultid="4845" />
                    <RANKING order="6" place="-1" resultid="3439" />
                    <RANKING order="7" place="-1" resultid="5872" />
                    <RANKING order="8" place="-1" resultid="5959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4801" />
                    <RANKING order="2" place="2" resultid="4610" />
                    <RANKING order="3" place="3" resultid="4828" />
                    <RANKING order="4" place="-1" resultid="3455" />
                    <RANKING order="5" place="-1" resultid="4071" />
                    <RANKING order="6" place="-1" resultid="5619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5683" />
                    <RANKING order="2" place="2" resultid="4969" />
                    <RANKING order="3" place="3" resultid="2522" />
                    <RANKING order="4" place="4" resultid="3850" />
                    <RANKING order="5" place="5" resultid="2583" />
                    <RANKING order="6" place="6" resultid="3582" />
                    <RANKING order="7" place="7" resultid="3802" />
                    <RANKING order="8" place="8" resultid="4864" />
                    <RANKING order="9" place="-1" resultid="2635" />
                    <RANKING order="10" place="-1" resultid="3052" />
                    <RANKING order="11" place="-1" resultid="4100" />
                    <RANKING order="12" place="-1" resultid="5657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2539" />
                    <RANKING order="2" place="2" resultid="3061" />
                    <RANKING order="3" place="3" resultid="4837" />
                    <RANKING order="4" place="4" resultid="3823" />
                    <RANKING order="5" place="5" resultid="2441" />
                    <RANKING order="6" place="6" resultid="6243" />
                    <RANKING order="7" place="-1" resultid="3512" />
                    <RANKING order="8" place="-1" resultid="5448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6109" />
                    <RANKING order="2" place="2" resultid="4668" />
                    <RANKING order="3" place="3" resultid="2868" />
                    <RANKING order="4" place="4" resultid="4928" />
                    <RANKING order="5" place="5" resultid="2687" />
                    <RANKING order="6" place="-1" resultid="5540" />
                    <RANKING order="7" place="-1" resultid="4751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4958" />
                    <RANKING order="2" place="2" resultid="3651" />
                    <RANKING order="3" place="3" resultid="2432" />
                    <RANKING order="4" place="-1" resultid="3865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1638" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4818" />
                    <RANKING order="2" place="2" resultid="4710" />
                    <RANKING order="3" place="3" resultid="4214" />
                    <RANKING order="4" place="4" resultid="3598" />
                    <RANKING order="5" place="-1" resultid="5886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1639" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4920" />
                    <RANKING order="2" place="2" resultid="5010" />
                    <RANKING order="3" place="3" resultid="4572" />
                    <RANKING order="4" place="4" resultid="3589" />
                    <RANKING order="5" place="-1" resultid="4028" />
                    <RANKING order="6" place="-1" resultid="5896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1640" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4644" />
                    <RANKING order="2" place="2" resultid="4982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1641" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1642" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1643" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1644" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7762" daytime="10:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7763" daytime="10:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7764" daytime="10:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7765" daytime="10:47" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7766" daytime="10:51" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7767" daytime="10:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7768" daytime="10:58" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7769" daytime="11:02" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7770" daytime="11:05" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7771" daytime="11:08" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7772" daytime="11:12" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7773" daytime="11:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7774" daytime="11:18" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1645" daytime="11:21" gender="F" number="36" order="40" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1646" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2667" />
                    <RANKING order="2" place="2" resultid="5177" />
                    <RANKING order="3" place="3" resultid="6474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1647" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7140" />
                    <RANKING order="2" place="2" resultid="3932" />
                    <RANKING order="3" place="3" resultid="5976" />
                    <RANKING order="4" place="4" resultid="2708" />
                    <RANKING order="5" place="5" resultid="6472" />
                    <RANKING order="6" place="6" resultid="4991" />
                    <RANKING order="7" place="-1" resultid="4262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1648" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5927" />
                    <RANKING order="2" place="2" resultid="4148" />
                    <RANKING order="3" place="3" resultid="4118" />
                    <RANKING order="4" place="4" resultid="6129" />
                    <RANKING order="5" place="5" resultid="6042" />
                    <RANKING order="6" place="6" resultid="6374" />
                    <RANKING order="7" place="-1" resultid="5015" />
                    <RANKING order="8" place="-1" resultid="5037" />
                    <RANKING order="9" place="-1" resultid="5700" />
                    <RANKING order="10" place="-1" resultid="5839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1649" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3714" />
                    <RANKING order="2" place="2" resultid="5920" />
                    <RANKING order="3" place="3" resultid="7074" />
                    <RANKING order="4" place="4" resultid="3913" />
                    <RANKING order="5" place="5" resultid="3661" />
                    <RANKING order="6" place="6" resultid="4523" />
                    <RANKING order="7" place="7" resultid="4042" />
                    <RANKING order="8" place="-1" resultid="5422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5749" />
                    <RANKING order="2" place="2" resultid="5130" />
                    <RANKING order="3" place="3" resultid="5608" />
                    <RANKING order="4" place="4" resultid="5584" />
                    <RANKING order="5" place="-1" resultid="5393" />
                    <RANKING order="6" place="-1" resultid="6271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4400" />
                    <RANKING order="2" place="2" resultid="3844" />
                    <RANKING order="3" place="3" resultid="4855" />
                    <RANKING order="4" place="4" resultid="3502" />
                    <RANKING order="5" place="5" resultid="3814" />
                    <RANKING order="6" place="6" resultid="6381" />
                    <RANKING order="7" place="7" resultid="3898" />
                    <RANKING order="8" place="-1" resultid="6049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5489" />
                    <RANKING order="2" place="2" resultid="5097" />
                    <RANKING order="3" place="3" resultid="2515" />
                    <RANKING order="4" place="4" resultid="5668" />
                    <RANKING order="5" place="5" resultid="6204" />
                    <RANKING order="6" place="6" resultid="5388" />
                    <RANKING order="7" place="-1" resultid="5602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1653" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4899" />
                    <RANKING order="2" place="2" resultid="4544" />
                    <RANKING order="3" place="3" resultid="2861" />
                    <RANKING order="4" place="4" resultid="3677" />
                    <RANKING order="5" place="5" resultid="3668" />
                    <RANKING order="6" place="6" resultid="2570" />
                    <RANKING order="7" place="7" resultid="6081" />
                    <RANKING order="8" place="-1" resultid="2841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1654" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4039" />
                    <RANKING order="2" place="2" resultid="3410" />
                    <RANKING order="3" place="3" resultid="4906" />
                    <RANKING order="4" place="4" resultid="4442" />
                    <RANKING order="5" place="5" resultid="4700" />
                    <RANKING order="6" place="6" resultid="4018" />
                    <RANKING order="7" place="7" resultid="3577" />
                    <RANKING order="8" place="-1" resultid="5374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1655" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4706" />
                    <RANKING order="2" place="2" resultid="5350" />
                    <RANKING order="3" place="3" resultid="4495" />
                    <RANKING order="4" place="4" resultid="3558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1656" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4738" />
                    <RANKING order="2" place="2" resultid="3570" />
                    <RANKING order="3" place="3" resultid="2477" />
                    <RANKING order="4" place="4" resultid="3551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1657" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3486" />
                    <RANKING order="2" place="2" resultid="3921" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1658" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1659" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1660" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1661" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7775" daytime="11:21" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7776" daytime="11:23" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7777" daytime="11:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7778" daytime="11:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7779" daytime="11:28" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7780" daytime="11:29" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7781" daytime="11:31" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7782" daytime="11:32" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7783" daytime="11:33" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7784" daytime="11:34" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7785" daytime="11:36" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7786" daytime="11:37" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7787" daytime="11:38" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1662" daytime="11:39" gender="M" number="37" order="41" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1663" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6344" />
                    <RANKING order="2" place="2" resultid="7232" />
                    <RANKING order="3" place="3" resultid="4243" />
                    <RANKING order="4" place="4" resultid="7066" />
                    <RANKING order="5" place="5" resultid="6168" />
                    <RANKING order="6" place="-1" resultid="2643" />
                    <RANKING order="7" place="-1" resultid="6490" />
                    <RANKING order="8" place="-1" resultid="7203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1664" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4385" />
                    <RANKING order="2" place="2" resultid="5691" />
                    <RANKING order="3" place="3" resultid="5182" />
                    <RANKING order="4" place="4" resultid="5171" />
                    <RANKING order="5" place="5" resultid="4617" />
                    <RANKING order="6" place="6" resultid="2793" />
                    <RANKING order="7" place="7" resultid="5157" />
                    <RANKING order="8" place="8" resultid="5092" />
                    <RANKING order="9" place="9" resultid="5188" />
                    <RANKING order="10" place="10" resultid="5122" />
                    <RANKING order="11" place="11" resultid="2754" />
                    <RANKING order="12" place="-1" resultid="2750" />
                    <RANKING order="13" place="-1" resultid="5111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1665" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2799" />
                    <RANKING order="2" place="2" resultid="6455" />
                    <RANKING order="3" place="3" resultid="4001" />
                    <RANKING order="4" place="4" resultid="5695" />
                    <RANKING order="5" place="5" resultid="4330" />
                    <RANKING order="6" place="6" resultid="2910" />
                    <RANKING order="7" place="7" resultid="2904" />
                    <RANKING order="8" place="8" resultid="2728" />
                    <RANKING order="9" place="9" resultid="3244" />
                    <RANKING order="10" place="10" resultid="2899" />
                    <RANKING order="11" place="11" resultid="2894" />
                    <RANKING order="12" place="12" resultid="3249" />
                    <RANKING order="13" place="13" resultid="6330" />
                    <RANKING order="14" place="14" resultid="2759" />
                    <RANKING order="15" place="15" resultid="2941" />
                    <RANKING order="16" place="16" resultid="5194" />
                    <RANKING order="17" place="17" resultid="5066" />
                    <RANKING order="18" place="-1" resultid="2745" />
                    <RANKING order="19" place="-1" resultid="2960" />
                    <RANKING order="20" place="-1" resultid="5914" />
                    <RANKING order="21" place="-1" resultid="6336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1666" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5984" />
                    <RANKING order="2" place="2" resultid="5520" />
                    <RANKING order="3" place="3" resultid="5481" />
                    <RANKING order="4" place="4" resultid="5302" />
                    <RANKING order="5" place="5" resultid="6156" />
                    <RANKING order="6" place="6" resultid="4943" />
                    <RANKING order="7" place="7" resultid="4846" />
                    <RANKING order="8" place="8" resultid="4792" />
                    <RANKING order="9" place="9" resultid="5085" />
                    <RANKING order="10" place="10" resultid="6303" />
                    <RANKING order="11" place="11" resultid="2985" />
                    <RANKING order="12" place="12" resultid="6316" />
                    <RANKING order="13" place="13" resultid="2885" />
                    <RANKING order="14" place="14" resultid="3752" />
                    <RANKING order="15" place="15" resultid="2920" />
                    <RANKING order="16" place="16" resultid="6034" />
                    <RANKING order="17" place="-1" resultid="2400" />
                    <RANKING order="18" place="-1" resultid="2927" />
                    <RANKING order="19" place="-1" resultid="4273" />
                    <RANKING order="20" place="-1" resultid="5024" />
                    <RANKING order="21" place="-1" resultid="7132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1667" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5372" />
                    <RANKING order="2" place="2" resultid="3035" />
                    <RANKING order="3" place="3" resultid="3239" />
                    <RANKING order="4" place="4" resultid="3746" />
                    <RANKING order="5" place="5" resultid="3766" />
                    <RANKING order="6" place="6" resultid="5578" />
                    <RANKING order="7" place="7" resultid="4611" />
                    <RANKING order="8" place="8" resultid="3818" />
                    <RANKING order="9" place="9" resultid="3758" />
                    <RANKING order="10" place="10" resultid="3227" />
                    <RANKING order="11" place="11" resultid="5595" />
                    <RANKING order="12" place="12" resultid="5613" />
                    <RANKING order="13" place="13" resultid="3187" />
                    <RANKING order="14" place="14" resultid="3906" />
                    <RANKING order="15" place="15" resultid="5770" />
                    <RANKING order="16" place="16" resultid="4342" />
                    <RANKING order="17" place="17" resultid="3696" />
                    <RANKING order="18" place="-1" resultid="3690" />
                    <RANKING order="19" place="-1" resultid="6309" />
                    <RANKING order="20" place="-1" resultid="6352" />
                    <RANKING order="21" place="-1" resultid="7316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1668" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3827" />
                    <RANKING order="2" place="2" resultid="3496" />
                    <RANKING order="3" place="3" resultid="3975" />
                    <RANKING order="4" place="4" resultid="6263" />
                    <RANKING order="5" place="5" resultid="4936" />
                    <RANKING order="6" place="6" resultid="5500" />
                    <RANKING order="7" place="7" resultid="3891" />
                    <RANKING order="8" place="8" resultid="4998" />
                    <RANKING order="9" place="9" resultid="4678" />
                    <RANKING order="10" place="-1" resultid="8077" />
                    <RANKING order="11" place="-1" resultid="5102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5379" />
                    <RANKING order="2" place="2" resultid="6436" />
                    <RANKING order="3" place="3" resultid="3062" />
                    <RANKING order="4" place="4" resultid="4511" />
                    <RANKING order="5" place="5" resultid="2613" />
                    <RANKING order="6" place="6" resultid="6244" />
                    <RANKING order="7" place="7" resultid="2442" />
                    <RANKING order="8" place="8" resultid="6250" />
                    <RANKING order="9" place="9" resultid="3684" />
                    <RANKING order="10" place="10" resultid="4408" />
                    <RANKING order="11" place="11" resultid="5525" />
                    <RANKING order="12" place="-1" resultid="4563" />
                    <RANKING order="13" place="-1" resultid="5116" />
                    <RANKING order="14" place="-1" resultid="5305" />
                    <RANKING order="15" place="-1" resultid="5341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1670" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5782" />
                    <RANKING order="2" place="2" resultid="5338" />
                    <RANKING order="3" place="3" resultid="3139" />
                    <RANKING order="4" place="4" resultid="6223" />
                    <RANKING order="5" place="5" resultid="5455" />
                    <RANKING order="6" place="6" resultid="2554" />
                    <RANKING order="7" place="7" resultid="5258" />
                    <RANKING order="8" place="8" resultid="3170" />
                    <RANKING order="9" place="-1" resultid="4454" />
                    <RANKING order="10" place="-1" resultid="4695" />
                    <RANKING order="11" place="-1" resultid="7061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1671" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5311" />
                    <RANKING order="2" place="2" resultid="3461" />
                    <RANKING order="3" place="3" resultid="3371" />
                    <RANKING order="4" place="4" resultid="2695" />
                    <RANKING order="5" place="5" resultid="5934" />
                    <RANKING order="6" place="6" resultid="3608" />
                    <RANKING order="7" place="7" resultid="5967" />
                    <RANKING order="8" place="8" resultid="8005" />
                    <RANKING order="9" place="-1" resultid="3384" />
                    <RANKING order="10" place="-1" resultid="3400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1672" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5427" />
                    <RANKING order="2" place="2" resultid="5467" />
                    <RANKING order="3" place="3" resultid="2411" />
                    <RANKING order="4" place="4" resultid="3599" />
                    <RANKING order="5" place="-1" resultid="4447" />
                    <RANKING order="6" place="-1" resultid="5879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1673" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4733" />
                    <RANKING order="2" place="2" resultid="4921" />
                    <RANKING order="3" place="3" resultid="3618" />
                    <RANKING order="4" place="4" resultid="3633" />
                    <RANKING order="5" place="5" resultid="3590" />
                    <RANKING order="6" place="-1" resultid="4029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1674" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3417" />
                    <RANKING order="2" place="2" resultid="4983" />
                    <RANKING order="3" place="3" resultid="5799" />
                    <RANKING order="4" place="-1" resultid="4645" />
                    <RANKING order="5" place="-1" resultid="5890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1675" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3376" />
                    <RANKING order="2" place="2" resultid="3873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1676" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1677" agemax="94" agemin="90" name="N: 90 - 94 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1678" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7788" daytime="11:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7789" daytime="11:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7790" daytime="11:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7791" daytime="11:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7792" daytime="11:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7793" daytime="11:47" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7794" daytime="11:48" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7795" daytime="11:49" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7796" daytime="11:51" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7797" daytime="11:52" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7798" daytime="11:53" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7799" daytime="11:54" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7800" daytime="11:55" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7801" daytime="11:56" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7802" daytime="11:58" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7803" daytime="11:59" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7804" daytime="12:00" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7805" daytime="12:01" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7806" daytime="12:02" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7807" daytime="12:03" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="7808" daytime="12:04" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="7809" daytime="12:05" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="7810" daytime="12:06" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="7811" daytime="12:07" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="7812" daytime="12:08" number="25" order="25" status="OFFICIAL" />
                <HEAT heatid="7813" daytime="12:10" number="26" order="26" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1679" daytime="12:11" gender="X" number="38" order="42" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2352" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5210" />
                    <RANKING order="2" place="2" resultid="2770" />
                    <RANKING order="3" place="-1" resultid="2772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2353" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5209" />
                    <RANKING order="2" place="2" resultid="5988" />
                    <RANKING order="3" place="3" resultid="5260" />
                    <RANKING order="4" place="4" resultid="4355" />
                    <RANKING order="5" place="5" resultid="6392" />
                    <RANKING order="6" place="6" resultid="6390" />
                    <RANKING order="7" place="7" resultid="6399" />
                    <RANKING order="8" place="-1" resultid="5843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2354" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5542" />
                    <RANKING order="2" place="2" resultid="5725" />
                    <RANKING order="3" place="3" resultid="3853" />
                    <RANKING order="4" place="4" resultid="4945" />
                    <RANKING order="5" place="5" resultid="3783" />
                    <RANKING order="6" place="6" resultid="5623" />
                    <RANKING order="7" place="7" resultid="4357" />
                    <RANKING order="8" place="-1" resultid="5394" />
                    <RANKING order="9" place="-1" resultid="5726" />
                    <RANKING order="10" place="-1" resultid="6286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2355" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5544" />
                    <RANKING order="2" place="2" resultid="4575" />
                    <RANKING order="3" place="3" resultid="5551" />
                    <RANKING order="4" place="4" resultid="3697" />
                    <RANKING order="5" place="-1" resultid="6285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2356" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4765" />
                    <RANKING order="2" place="2" resultid="5398" />
                    <RANKING order="3" place="3" resultid="4577" />
                    <RANKING order="4" place="-1" resultid="3418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2357" agemax="319" agemin="280" name="F: 280 - 319 lat " calculate="TOTAL" />
                <AGEGROUP agegroupid="2358" agemax="359" agemin="320" name="G: 320 - 359 lat " calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7814" daytime="12:11" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7815" daytime="12:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7816" daytime="12:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7817" daytime="12:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7818" daytime="12:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7819" daytime="12:27" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1693" daytime="12:30" gender="F" number="39" order="43" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1694" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2668" />
                    <RANKING order="2" place="-1" resultid="2703" />
                    <RANKING order="3" place="-1" resultid="5078" />
                    <RANKING order="4" place="-1" resultid="5858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1695" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5818" />
                    <RANKING order="2" place="2" resultid="2530" />
                    <RANKING order="3" place="3" resultid="5072" />
                    <RANKING order="4" place="4" resultid="4503" />
                    <RANKING order="5" place="5" resultid="5589" />
                    <RANKING order="6" place="6" resultid="5164" />
                    <RANKING order="7" place="7" resultid="8061" />
                    <RANKING order="8" place="8" resultid="4084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1696" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5358" />
                    <RANKING order="2" place="2" resultid="4149" />
                    <RANKING order="3" place="3" resultid="4336" />
                    <RANKING order="4" place="4" resultid="6147" />
                    <RANKING order="5" place="5" resultid="4284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1697" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2817" />
                    <RANKING order="2" place="2" resultid="3721" />
                    <RANKING order="3" place="3" resultid="4266" />
                    <RANKING order="4" place="4" resultid="3738" />
                    <RANKING order="5" place="5" resultid="7075" />
                    <RANKING order="6" place="6" resultid="3914" />
                    <RANKING order="7" place="7" resultid="4524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1698" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4717" />
                    <RANKING order="2" place="2" resultid="3838" />
                    <RANKING order="3" place="3" resultid="3730" />
                    <RANKING order="4" place="4" resultid="7251" />
                    <RANKING order="5" place="5" resultid="2675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1699" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3476" />
                    <RANKING order="2" place="2" resultid="4281" />
                    <RANKING order="3" place="3" resultid="2835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1700" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4478" />
                    <RANKING order="2" place="2" resultid="5603" />
                    <RANKING order="3" place="3" resultid="4090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1701" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4687" />
                    <RANKING order="2" place="2" resultid="4469" />
                    <RANKING order="3" place="3" resultid="2876" />
                    <RANKING order="4" place="-1" resultid="2842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1702" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3545" />
                    <RANKING order="2" place="2" resultid="5462" />
                    <RANKING order="3" place="3" resultid="3984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1703" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5062" />
                    <RANKING order="2" place="2" resultid="4496" />
                    <RANKING order="3" place="3" resultid="3622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1704" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1705" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1706" agemax="84" agemin="80" name="L: 80 - 84 lat " />
                <AGEGROUP agegroupid="1707" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1708" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1709" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8018" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8019" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8020" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8021" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8022" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8023" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8024" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8025" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1710" daytime="13:43" gender="M" number="40" order="44" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1711" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2606" />
                    <RANKING order="2" place="2" resultid="2510" />
                    <RANKING order="3" place="3" resultid="7233" />
                    <RANKING order="4" place="4" resultid="4871" />
                    <RANKING order="5" place="5" resultid="4724" />
                    <RANKING order="6" place="6" resultid="4138" />
                    <RANKING order="7" place="-1" resultid="7157" />
                    <RANKING order="8" place="-1" resultid="7195" />
                    <RANKING order="9" place="-1" resultid="7204" />
                    <RANKING order="10" place="-1" resultid="7213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1712" agemax="29" agemin="25" name="A: 25 - 29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5792" />
                    <RANKING order="2" place="2" resultid="3482" />
                    <RANKING order="3" place="3" resultid="4386" />
                    <RANKING order="4" place="4" resultid="2794" />
                    <RANKING order="5" place="5" resultid="5123" />
                    <RANKING order="6" place="6" resultid="3184" />
                    <RANKING order="7" place="7" resultid="3233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1713" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4126" />
                    <RANKING order="2" place="2" resultid="2549" />
                    <RANKING order="3" place="3" resultid="2560" />
                    <RANKING order="4" place="4" resultid="5033" />
                    <RANKING order="5" place="5" resultid="5195" />
                    <RANKING order="6" place="6" resultid="4320" />
                    <RANKING order="7" place="7" resultid="2950" />
                    <RANKING order="8" place="-1" resultid="2729" />
                    <RANKING order="9" place="-1" resultid="4144" />
                    <RANKING order="10" place="-1" resultid="4975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1714" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3213" />
                    <RANKING order="2" place="2" resultid="4424" />
                    <RANKING order="3" place="3" resultid="5320" />
                    <RANKING order="4" place="4" resultid="2934" />
                    <RANKING order="5" place="5" resultid="5873" />
                    <RANKING order="6" place="6" resultid="3532" />
                    <RANKING order="7" place="-1" resultid="2734" />
                    <RANKING order="8" place="-1" resultid="5147" />
                    <RANKING order="9" place="-1" resultid="5985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1715" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4300" />
                    <RANKING order="2" place="2" resultid="3036" />
                    <RANKING order="3" place="3" resultid="2453" />
                    <RANKING order="4" place="4" resultid="3773" />
                    <RANKING order="5" place="-1" resultid="3456" />
                    <RANKING order="6" place="-1" resultid="3925" />
                    <RANKING order="7" place="-1" resultid="4315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1716" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3517" />
                    <RANKING order="2" place="2" resultid="4079" />
                    <RANKING order="3" place="3" resultid="3045" />
                    <RANKING order="4" place="4" resultid="6267" />
                    <RANKING order="5" place="5" resultid="5765" />
                    <RANKING order="6" place="6" resultid="2524" />
                    <RANKING order="7" place="7" resultid="4108" />
                    <RANKING order="8" place="8" resultid="4051" />
                    <RANKING order="9" place="9" resultid="4548" />
                    <RANKING order="10" place="10" resultid="3642" />
                    <RANKING order="11" place="-1" resultid="2417" />
                    <RANKING order="12" place="-1" resultid="4810" />
                    <RANKING order="13" place="-1" resultid="5139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1717" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2597" />
                    <RANKING order="2" place="2" resultid="6437" />
                    <RANKING order="3" place="3" resultid="3513" />
                    <RANKING order="4" place="4" resultid="2500" />
                    <RANKING order="5" place="5" resultid="4409" />
                    <RANKING order="6" place="6" resultid="2578" />
                    <RANKING order="7" place="7" resultid="4154" />
                    <RANKING order="8" place="8" resultid="4564" />
                    <RANKING order="9" place="9" resultid="4013" />
                    <RANKING order="10" place="-1" resultid="6237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1718" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4309" />
                    <RANKING order="2" place="2" resultid="2869" />
                    <RANKING order="3" place="3" resultid="4696" />
                    <RANKING order="4" place="4" resultid="8072" />
                    <RANKING order="5" place="5" resultid="6074" />
                    <RANKING order="6" place="6" resultid="2680" />
                    <RANKING order="7" place="7" resultid="5049" />
                    <RANKING order="8" place="8" resultid="5259" />
                    <RANKING order="9" place="-1" resultid="2850" />
                    <RANKING order="10" place="-1" resultid="6229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1719" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8060" />
                    <RANKING order="2" place="2" resultid="2396" />
                    <RANKING order="3" place="3" resultid="3401" />
                    <RANKING order="4" place="4" resultid="5943" />
                    <RANKING order="5" place="5" resultid="2433" />
                    <RANKING order="6" place="6" resultid="3609" />
                    <RANKING order="7" place="-1" resultid="7242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1720" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4819" />
                    <RANKING order="2" place="2" resultid="4487" />
                    <RANKING order="3" place="3" resultid="2857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1721" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5011" />
                    <RANKING order="2" place="2" resultid="6138" />
                    <RANKING order="3" place="3" resultid="4532" />
                    <RANKING order="4" place="4" resultid="4253" />
                    <RANKING order="5" place="5" resultid="4573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1722" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1723" agemax="84" agemin="80" name="L: 80 - 84 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3874" />
                    <RANKING order="2" place="-1" resultid="7181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1724" agemax="89" agemin="85" name="M: 85 - 89 lat " />
                <AGEGROUP agegroupid="1725" agemax="94" agemin="90" name="N: 90 - 94 lat " />
                <AGEGROUP agegroupid="1726" agemax="-1" agemin="95" name="O: 95 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8043" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8044" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8045" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8046" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8047" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8048" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8049" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8050" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8051" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8052" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="8053" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="8054" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="8055" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="8056" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="8057" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="8058" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" name="MUKS Lider Chełm" nation="POL">
          <CONTACT city="Chełm" email="agnieszkakargol@onet.eu" name="Kargol" phone="798408133" state="LUBEL" street="Połaniecka 10" zip="22-100" />
          <ATHLETES>
            <ATHLETE birthdate="1989-08-19" firstname="Agnieszka" gender="F" lastname="Kargol" nation="POL" license="100403100009" athleteid="2360">
              <RESULTS>
                <RESULT eventid="1058" points="523" reactiontime="+77" swimtime="00:00:28.85" resultid="2361" heatid="7344" lane="3" entrytime="00:00:27.47" entrycourse="SCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1183" points="575" reactiontime="+72" swimtime="00:00:30.90" resultid="2362" heatid="7441" lane="3" entrytime="00:00:30.01" entrycourse="SCM" />
                <RESULT eventid="1285" points="562" swimtime="00:01:09.95" resultid="2363" heatid="7537" lane="5" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="609" reactiontime="+78" swimtime="00:00:28.76" resultid="2364" heatid="7621" lane="3" entrytime="00:00:27.70" entrycourse="SCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1453" points="547" reactiontime="+76" swimtime="00:01:07.51" resultid="2365" heatid="7658" lane="3" entrytime="00:01:05.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1611" points="529" reactiontime="+70" swimtime="00:02:28.37" resultid="2366" heatid="7761" lane="4" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:51.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Tri Negu" nation="POL">
          <CONTACT city="Dawidy Bankowe" email="biuro@q-kwadrat.pl" name="Palysa" state="MAZ" street="Szlachecka 33" zip="05090" />
          <ATHLETES>
            <ATHLETE birthdate="1974-11-22" firstname="Pałysa" gender="M" lastname="Marek" nation="POL" athleteid="2368" />
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5130" name="TG Lage 1862" nation="GER" region="17">
          <CONTACT city="Lage" email="tg-schwimmen@gmx.de" name="Lange Ute" state="NO" street="Ringstr. 3" zip="32791" />
          <ATHLETES>
            <ATHLETE birthdate="1968-04-07" firstname="Konstantin" gender="M" lastname="Sklyar" nation="GER" license="321129" athleteid="2371">
              <RESULTS>
                <RESULT eventid="1109" points="332" reactiontime="+94" swimtime="00:02:38.85" resultid="2372" heatid="7400" lane="3" entrytime="00:02:43.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:16.60" />
                    <SPLIT distance="150" swimtime="00:02:02.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="325" reactiontime="+98" swimtime="00:02:55.50" resultid="2373" heatid="7479" lane="3" entrytime="00:03:00.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                    <SPLIT distance="100" swimtime="00:01:25.03" />
                    <SPLIT distance="150" swimtime="00:02:10.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="342" reactiontime="+86" swimtime="00:01:04.25" resultid="2374" heatid="7516" lane="4" entrytime="00:01:03.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="3 start w bloku." eventid="1336" status="DSQ" swimtime="00:02:50.26" resultid="2375" heatid="7569" lane="5" entrytime="00:02:48.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:20.25" />
                    <SPLIT distance="150" swimtime="00:02:07.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="317" reactiontime="+83" swimtime="00:00:31.96" resultid="2376" heatid="7635" lane="3" entrytime="00:00:31.85" entrycourse="SCM" />
                <RESULT eventid="1594" points="312" reactiontime="+87" swimtime="00:01:11.41" resultid="2378" heatid="7746" lane="6" entrytime="00:01:10.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="305" reactiontime="+96" swimtime="00:05:49.56" resultid="7984" heatid="7974" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="150" swimtime="00:02:05.78" />
                    <SPLIT distance="200" swimtime="00:02:52.72" />
                    <SPLIT distance="250" swimtime="00:03:42.72" />
                    <SPLIT distance="300" swimtime="00:04:33.24" />
                    <SPLIT distance="350" swimtime="00:05:12.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="UKS SP8 Chrzanów" nation="POL" region="06">
          <CONTACT email="abalp@poczta.onet.pl" name="Zabrzański Alfred" phone="692076808" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="2390">
              <RESULTS>
                <RESULT eventid="1075" points="292" reactiontime="+89" swimtime="00:00:30.57" resultid="2391" heatid="7361" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2392" heatid="7911" lane="6" entrytime="00:24:45.00" />
                <RESULT eventid="1200" points="193" reactiontime="+76" swimtime="00:00:39.06" resultid="2393" heatid="7447" lane="1" entrytime="00:00:40.80" />
                <RESULT eventid="1268" points="277" reactiontime="+90" swimtime="00:01:08.89" resultid="2394" heatid="7511" lane="1" entrytime="00:01:09.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="249" swimtime="00:02:37.91" resultid="2395" heatid="7694" lane="5" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:15.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="215" reactiontime="+98" swimtime="00:05:54.65" resultid="2396" heatid="8048" lane="2" entrytime="00:06:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:01:19.94" />
                    <SPLIT distance="150" swimtime="00:02:03.68" />
                    <SPLIT distance="200" swimtime="00:02:49.87" />
                    <SPLIT distance="250" swimtime="00:03:36.85" />
                    <SPLIT distance="300" swimtime="00:04:23.07" />
                    <SPLIT distance="350" swimtime="00:05:10.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Niezrzeszeni" nation="POL">
          <CONTACT email="piotr_urbanczyk@onet.pl" name="PIOTR URBAŃCZYK" phone="608172201" />
          <ATHLETES>
            <ATHLETE birthdate="1937-09-19" firstname="Zygmunt" gender="M" lastname="Lewandowski" nation="POL" athleteid="2381">
              <RESULTS>
                <RESULT eventid="1075" points="127" reactiontime="+99" swimtime="00:00:40.38" resultid="2382" heatid="7349" lane="6" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="1165" points="101" reactiontime="+115" swimtime="00:30:22.20" resultid="2383" heatid="7908" lane="6" entrytime="00:35:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.03" />
                    <SPLIT distance="100" swimtime="00:01:46.64" />
                    <SPLIT distance="150" swimtime="00:02:44.13" />
                    <SPLIT distance="200" swimtime="00:03:42.55" />
                    <SPLIT distance="250" swimtime="00:04:40.35" />
                    <SPLIT distance="300" swimtime="00:05:38.87" />
                    <SPLIT distance="350" swimtime="00:06:37.08" />
                    <SPLIT distance="400" swimtime="00:07:37.46" />
                    <SPLIT distance="450" swimtime="00:08:38.95" />
                    <SPLIT distance="500" swimtime="00:09:40.57" />
                    <SPLIT distance="550" swimtime="00:10:43.53" />
                    <SPLIT distance="600" swimtime="00:11:45.77" />
                    <SPLIT distance="650" swimtime="00:12:48.37" />
                    <SPLIT distance="700" swimtime="00:13:51.33" />
                    <SPLIT distance="750" swimtime="00:14:55.82" />
                    <SPLIT distance="800" swimtime="00:15:56.97" />
                    <SPLIT distance="850" swimtime="00:16:58.43" />
                    <SPLIT distance="900" swimtime="00:17:59.81" />
                    <SPLIT distance="950" swimtime="00:19:01.63" />
                    <SPLIT distance="1000" swimtime="00:20:04.49" />
                    <SPLIT distance="1050" swimtime="00:21:08.71" />
                    <SPLIT distance="1100" swimtime="00:22:10.47" />
                    <SPLIT distance="1150" swimtime="00:23:11.67" />
                    <SPLIT distance="1200" swimtime="00:24:13.58" />
                    <SPLIT distance="1250" swimtime="00:25:16.88" />
                    <SPLIT distance="1300" swimtime="00:26:20.14" />
                    <SPLIT distance="1350" swimtime="00:27:21.53" />
                    <SPLIT distance="1400" swimtime="00:28:21.22" />
                    <SPLIT distance="1450" swimtime="00:29:22.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="90" swimtime="00:01:52.94" resultid="2384" heatid="7539" lane="5" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="79" reactiontime="+108" swimtime="00:00:50.72" resultid="2385" heatid="7623" lane="3" entrytime="00:01:05.00" entrycourse="SCM" />
                <RESULT eventid="1504" points="103" swimtime="00:03:31.57" resultid="2386" heatid="7688" lane="5" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.34" />
                    <SPLIT distance="100" swimtime="00:01:42.22" />
                    <SPLIT distance="150" swimtime="00:02:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="2387" heatid="7738" lane="1" entrytime="00:02:05.00" entrycourse="SCM" />
                <RESULT eventid="1710" points="98" swimtime="00:07:41.18" resultid="2388" heatid="8045" lane="5" entrytime="00:08:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.66" />
                    <SPLIT distance="100" swimtime="00:01:49.40" />
                    <SPLIT distance="150" swimtime="00:02:48.22" />
                    <SPLIT distance="200" swimtime="00:03:47.51" />
                    <SPLIT distance="250" swimtime="00:04:47.80" />
                    <SPLIT distance="300" swimtime="00:05:44.96" />
                    <SPLIT distance="350" swimtime="00:06:43.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Michał" gender="M" lastname="Syryca" nation="POL" athleteid="2397">
              <RESULTS>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="2398" heatid="7456" lane="1" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="1436" points="251" swimtime="00:00:34.52" resultid="2399" heatid="7639" lane="5" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="2400" heatid="7801" lane="4" entrytime="00:00:38.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Włodzimierz " gender="M" lastname="Zieleziński" nation="POL" athleteid="2425">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="2426" heatid="7355" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1165" points="152" reactiontime="+121" swimtime="00:26:31.15" resultid="2427" heatid="7909" lane="1" entrytime="00:27:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="100" swimtime="00:01:28.96" />
                    <SPLIT distance="150" swimtime="00:02:20.08" />
                    <SPLIT distance="200" swimtime="00:03:12.38" />
                    <SPLIT distance="250" swimtime="00:04:04.81" />
                    <SPLIT distance="300" swimtime="00:04:57.75" />
                    <SPLIT distance="350" swimtime="00:05:50.53" />
                    <SPLIT distance="400" swimtime="00:06:44.00" />
                    <SPLIT distance="450" swimtime="00:07:37.51" />
                    <SPLIT distance="500" swimtime="00:08:30.41" />
                    <SPLIT distance="550" swimtime="00:09:24.28" />
                    <SPLIT distance="600" swimtime="00:10:18.39" />
                    <SPLIT distance="650" swimtime="00:11:12.27" />
                    <SPLIT distance="700" swimtime="00:12:05.85" />
                    <SPLIT distance="750" swimtime="00:13:00.13" />
                    <SPLIT distance="800" swimtime="00:13:53.98" />
                    <SPLIT distance="850" swimtime="00:14:47.48" />
                    <SPLIT distance="900" swimtime="00:15:41.64" />
                    <SPLIT distance="950" swimtime="00:16:37.12" />
                    <SPLIT distance="1000" swimtime="00:17:33.27" />
                    <SPLIT distance="1050" swimtime="00:18:27.83" />
                    <SPLIT distance="1100" swimtime="00:19:23.13" />
                    <SPLIT distance="1150" swimtime="00:20:17.91" />
                    <SPLIT distance="1200" swimtime="00:21:11.75" />
                    <SPLIT distance="1250" swimtime="00:22:05.87" />
                    <SPLIT distance="1300" swimtime="00:23:00.38" />
                    <SPLIT distance="1350" swimtime="00:23:54.53" />
                    <SPLIT distance="1400" swimtime="00:24:48.94" />
                    <SPLIT distance="1450" swimtime="00:25:41.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="159" reactiontime="+88" swimtime="00:00:41.72" resultid="2428" heatid="7446" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="2429" heatid="7505" lane="1" entrytime="00:01:18.00" />
                <RESULT eventid="1470" points="145" reactiontime="+90" swimtime="00:01:33.06" resultid="2430" heatid="7663" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="2431" heatid="7690" lane="3" entrytime="00:03:00.00" />
                <RESULT eventid="1628" points="131" reactiontime="+95" swimtime="00:03:28.76" resultid="2432" heatid="7765" lane="1" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                    <SPLIT distance="100" swimtime="00:01:40.86" />
                    <SPLIT distance="150" swimtime="00:02:35.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="176" reactiontime="+112" swimtime="00:06:19.65" resultid="2433" heatid="8047" lane="3" entrytime="00:06:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:01:24.97" />
                    <SPLIT distance="150" swimtime="00:02:13.72" />
                    <SPLIT distance="200" swimtime="00:03:03.50" />
                    <SPLIT distance="250" swimtime="00:03:54.18" />
                    <SPLIT distance="300" swimtime="00:04:43.97" />
                    <SPLIT distance="350" swimtime="00:05:34.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Szozda " gender="M" lastname="Zbigniew" nation="POL" athleteid="2434">
              <RESULTS>
                <RESULT eventid="1075" points="266" swimtime="00:00:31.55" resultid="2435" heatid="7359" lane="5" entrytime="00:00:31.70" />
                <RESULT eventid="1109" points="238" swimtime="00:02:57.43" resultid="2436" heatid="7397" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:21.68" />
                    <SPLIT distance="150" swimtime="00:02:14.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="237" reactiontime="+83" swimtime="00:00:36.49" resultid="2437" heatid="7449" lane="4" entrytime="00:00:36.80" />
                <RESULT eventid="1302" points="278" reactiontime="+104" swimtime="00:01:17.69" resultid="2438" heatid="7547" lane="6" entrytime="00:01:19.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="275" swimtime="00:00:33.52" resultid="2439" heatid="7632" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1470" points="222" reactiontime="+75" swimtime="00:01:20.73" resultid="2440" heatid="7664" lane="3" entrytime="00:01:23.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="189" reactiontime="+78" swimtime="00:03:04.81" resultid="2441" heatid="7766" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="100" swimtime="00:01:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="269" reactiontime="+101" swimtime="00:00:39.08" resultid="2442" heatid="7796" lane="3" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-18" firstname="Kazimierz" gender="M" lastname="Sinicki" nation="POL" athleteid="2444">
              <RESULTS>
                <RESULT eventid="1075" points="342" reactiontime="+85" swimtime="00:00:29.02" resultid="2445" heatid="7365" lane="3" entrytime="00:00:29.50" />
                <RESULT eventid="1268" points="313" reactiontime="+86" swimtime="00:01:06.16" resultid="2446" heatid="7511" lane="3" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="270" reactiontime="+85" swimtime="00:00:33.71" resultid="2447" heatid="7629" lane="3" entrytime="00:00:35.50" />
                <RESULT eventid="1504" points="269" reactiontime="+94" swimtime="00:02:33.93" resultid="2448" heatid="7695" lane="1" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:55.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="DAMIAN " gender="M" lastname="KĄDZIELEWSKI" nation="POL" athleteid="2454">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="2455" heatid="7350" lane="4" entrytime="00:00:38.24" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="2456" heatid="7501" lane="4" entrytime="00:01:40.10" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="2457" heatid="7688" lane="6" entrytime="00:04:02.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="JUDYTA " gender="F" lastname="SOŁTYK" nation="POL" athleteid="2459">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1319" points="372" reactiontime="+89" swimtime="00:02:47.90" resultid="2460" heatid="7563" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:19.84" />
                    <SPLIT distance="150" swimtime="00:02:04.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="463" reactiontime="+86" swimtime="00:02:23.61" resultid="2461" heatid="7683" lane="4" entrytime="00:02:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:09.67" />
                    <SPLIT distance="150" swimtime="00:01:46.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="409" reactiontime="+84" swimtime="00:01:14.13" resultid="2462" heatid="7735" lane="6" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="Alina " gender="F" lastname="Wieczorkiewicz" nation="POL" athleteid="2471">
              <RESULTS>
                <RESULT eventid="1058" points="18" reactiontime="+126" swimtime="00:01:27.27" resultid="2472" heatid="7332" lane="2" entrytime="00:01:20.00" />
                <RESULT eventid="1183" points="30" reactiontime="+105" swimtime="00:01:22.21" resultid="2473" heatid="7432" lane="5" entrytime="00:01:25.00" />
                <RESULT eventid="1285" points="25" reactiontime="+116" swimtime="00:03:16.80" resultid="2474" heatid="7526" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="27" reactiontime="+83" swimtime="00:03:02.90" resultid="2475" heatid="7649" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="25" reactiontime="+95" swimtime="00:06:46.53" resultid="2476" heatid="7754" lane="5" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:38.47" />
                    <SPLIT distance="100" swimtime="00:03:24.08" />
                    <SPLIT distance="150" swimtime="00:05:09.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="30" reactiontime="+126" swimtime="00:01:32.53" resultid="2477" heatid="7776" lane="6" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Patryk " gender="M" lastname="Poniatowski" nation="POL" athleteid="2478">
              <RESULTS>
                <RESULT eventid="1075" points="608" reactiontime="+76" swimtime="00:00:23.95" resultid="2479" heatid="7381" lane="1" entrytime="00:00:24.01" />
                <RESULT eventid="1268" points="606" reactiontime="+73" swimtime="00:00:53.09" resultid="2480" heatid="7525" lane="6" entrytime="00:00:54.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="549" reactiontime="+65" swimtime="00:00:27.61" resultid="2481" heatid="7460" lane="6" entrytime="00:00:27.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="2531">
              <RESULTS>
                <RESULT eventid="1075" points="395" reactiontime="+80" swimtime="00:00:27.65" resultid="2532" heatid="7369" lane="6" entrytime="00:00:28.25" />
                <RESULT eventid="1109" points="364" swimtime="00:02:34.08" resultid="2533" heatid="7403" lane="5" entrytime="00:02:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:11.20" />
                    <SPLIT distance="150" swimtime="00:01:57.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="399" reactiontime="+81" swimtime="00:01:01.04" resultid="2534" heatid="7518" lane="3" entrytime="00:01:01.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="378" reactiontime="+88" swimtime="00:01:10.19" resultid="2535" heatid="7552" lane="2" entrytime="00:01:10.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="384" swimtime="00:00:29.98" resultid="2536" heatid="7638" lane="5" entrytime="00:00:30.55" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="2537" heatid="7668" lane="6" entrytime="00:01:14.50" />
                <RESULT eventid="1594" points="357" reactiontime="+88" swimtime="00:01:08.31" resultid="2538" heatid="7749" lane="1" entrytime="00:01:08.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="281" reactiontime="+70" swimtime="00:02:41.94" resultid="2539" heatid="7769" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                    <SPLIT distance="100" swimtime="00:01:19.44" />
                    <SPLIT distance="150" swimtime="00:02:00.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="ANNA" gender="F" lastname="KOTUSIŃSKA " nation="POL" athleteid="2800">
              <RESULTS>
                <RESULT eventid="1251" points="222" swimtime="00:01:24.18" resultid="2801" heatid="7492" lane="5" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="195" reactiontime="+91" swimtime="00:00:42.00" resultid="2802" heatid="7616" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Igor" gender="M" lastname="Okarmus " nation="POL" athleteid="2803">
              <RESULTS>
                <RESULT eventid="1165" points="303" reactiontime="+116" swimtime="00:21:04.56" resultid="2804" heatid="7913" lane="1" entrytime="00:22:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:12.79" />
                    <SPLIT distance="150" swimtime="00:01:53.37" />
                    <SPLIT distance="200" swimtime="00:02:34.65" />
                    <SPLIT distance="250" swimtime="00:03:16.40" />
                    <SPLIT distance="300" swimtime="00:03:59.31" />
                    <SPLIT distance="350" swimtime="00:04:41.78" />
                    <SPLIT distance="400" swimtime="00:05:23.57" />
                    <SPLIT distance="450" swimtime="00:06:05.95" />
                    <SPLIT distance="500" swimtime="00:06:47.87" />
                    <SPLIT distance="550" swimtime="00:07:29.97" />
                    <SPLIT distance="600" swimtime="00:08:12.17" />
                    <SPLIT distance="650" swimtime="00:08:54.63" />
                    <SPLIT distance="700" swimtime="00:09:37.22" />
                    <SPLIT distance="750" swimtime="00:10:20.02" />
                    <SPLIT distance="800" swimtime="00:11:02.81" />
                    <SPLIT distance="850" swimtime="00:11:45.30" />
                    <SPLIT distance="900" swimtime="00:12:28.51" />
                    <SPLIT distance="950" swimtime="00:13:11.40" />
                    <SPLIT distance="1000" swimtime="00:13:54.29" />
                    <SPLIT distance="1050" swimtime="00:14:37.61" />
                    <SPLIT distance="1100" swimtime="00:15:21.16" />
                    <SPLIT distance="1150" swimtime="00:16:04.60" />
                    <SPLIT distance="1200" swimtime="00:16:47.37" />
                    <SPLIT distance="1250" swimtime="00:17:30.03" />
                    <SPLIT distance="1300" swimtime="00:18:13.91" />
                    <SPLIT distance="1350" swimtime="00:18:57.59" />
                    <SPLIT distance="1400" swimtime="00:19:40.59" />
                    <SPLIT distance="1450" swimtime="00:20:23.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-01" firstname="Jolanta" gender="F" lastname="Zawadzka" nation="POL" athleteid="2859">
              <RESULTS>
                <RESULT eventid="1419" points="184" reactiontime="+88" swimtime="00:00:42.85" resultid="2860" heatid="7615" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1645" points="245" swimtime="00:00:45.97" resultid="2861" heatid="7783" lane="2" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-16" firstname="Piotr" gender="M" lastname="Urbańczyk" nation="POL" athleteid="3026">
              <RESULTS>
                <RESULT eventid="1200" points="491" reactiontime="+63" swimtime="00:00:28.65" resultid="3027" heatid="7459" lane="2" entrytime="00:00:28.40" />
                <RESULT eventid="1470" points="498" reactiontime="+64" swimtime="00:01:01.72" resultid="3028" heatid="7674" lane="5" entrytime="00:01:00.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jolanta" gender="F" lastname="Lipińska " nation="POL" athleteid="3977">
              <RESULTS>
                <RESULT eventid="1092" points="33" reactiontime="+122" swimtime="00:06:26.32" resultid="3978" heatid="7382" lane="4" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.14" />
                    <SPLIT distance="100" swimtime="00:03:18.72" />
                    <SPLIT distance="150" swimtime="00:05:02.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="56" swimtime="00:05:51.61" resultid="3979" heatid="7462" lane="5" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.95" />
                    <SPLIT distance="100" swimtime="00:02:50.84" />
                    <SPLIT distance="150" swimtime="00:04:23.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="34" swimtime="00:02:57.23" resultid="3980" heatid="7526" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="12" reactiontime="+134" swimtime="00:01:44.91" resultid="3981" heatid="7612" lane="3" entrytime="00:01:45.00" />
                <RESULT eventid="1487" points="30" swimtime="00:05:56.27" resultid="3982" heatid="7675" lane="5" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.24" />
                    <SPLIT distance="100" swimtime="00:02:56.15" />
                    <SPLIT distance="150" swimtime="00:04:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="37" reactiontime="+86" swimtime="00:05:58.46" resultid="3983" heatid="7754" lane="1" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.23" />
                    <SPLIT distance="100" swimtime="00:02:53.07" />
                    <SPLIT distance="150" swimtime="00:04:26.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="38" reactiontime="+132" swimtime="00:11:36.80" resultid="3984" heatid="8019" lane="6" entrytime="00:11:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.23" />
                    <SPLIT distance="100" swimtime="00:02:51.92" />
                    <SPLIT distance="150" swimtime="00:04:19.41" />
                    <SPLIT distance="200" swimtime="00:05:48.24" />
                    <SPLIT distance="250" swimtime="00:07:16.64" />
                    <SPLIT distance="300" swimtime="00:08:43.48" />
                    <SPLIT distance="350" swimtime="00:10:11.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="KRZYSZTOF " gender="M" lastname="DRÓZD" nation="POL" athleteid="4002">
              <RESULTS>
                <RESULT eventid="1075" points="388" swimtime="00:00:27.83" resultid="4003" heatid="7374" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="4004" heatid="7546" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1504" points="288" reactiontime="+64" swimtime="00:02:30.32" resultid="4005" heatid="7695" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:08.67" />
                    <SPLIT distance="150" swimtime="00:01:49.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Norbert" gender="M" lastname="Tchorzewski " nation="POL" athleteid="4043">
              <RESULTS>
                <RESULT eventid="1075" points="303" reactiontime="+83" swimtime="00:00:30.20" resultid="4044" heatid="7361" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1165" points="230" reactiontime="+114" swimtime="00:23:05.50" resultid="4045" heatid="7912" lane="1" entrytime="00:23:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="150" swimtime="00:02:05.41" />
                    <SPLIT distance="200" swimtime="00:02:51.06" />
                    <SPLIT distance="250" swimtime="00:03:38.27" />
                    <SPLIT distance="300" swimtime="00:04:23.65" />
                    <SPLIT distance="350" swimtime="00:05:10.81" />
                    <SPLIT distance="400" swimtime="00:05:57.86" />
                    <SPLIT distance="450" swimtime="00:06:44.92" />
                    <SPLIT distance="500" swimtime="00:07:31.43" />
                    <SPLIT distance="550" swimtime="00:08:18.87" />
                    <SPLIT distance="600" swimtime="00:09:05.21" />
                    <SPLIT distance="650" swimtime="00:09:52.53" />
                    <SPLIT distance="700" swimtime="00:10:40.04" />
                    <SPLIT distance="750" swimtime="00:11:27.26" />
                    <SPLIT distance="800" swimtime="00:12:14.35" />
                    <SPLIT distance="850" swimtime="00:13:01.56" />
                    <SPLIT distance="900" swimtime="00:13:47.77" />
                    <SPLIT distance="950" swimtime="00:14:34.20" />
                    <SPLIT distance="1000" swimtime="00:15:21.90" />
                    <SPLIT distance="1050" swimtime="00:16:08.55" />
                    <SPLIT distance="1100" swimtime="00:16:55.00" />
                    <SPLIT distance="1150" swimtime="00:17:40.86" />
                    <SPLIT distance="1200" swimtime="00:18:27.84" />
                    <SPLIT distance="1250" swimtime="00:19:14.55" />
                    <SPLIT distance="1300" swimtime="00:20:01.27" />
                    <SPLIT distance="1350" swimtime="00:20:47.95" />
                    <SPLIT distance="1400" swimtime="00:21:34.46" />
                    <SPLIT distance="1450" swimtime="00:22:21.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="305" reactiontime="+82" swimtime="00:01:06.74" resultid="4046" heatid="7510" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="257" reactiontime="+81" swimtime="00:01:19.79" resultid="4047" heatid="7543" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="277" reactiontime="+82" swimtime="00:00:33.43" resultid="4048" heatid="7635" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1559" points="182" swimtime="00:06:55.41" resultid="4049" heatid="7977" lane="5" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="100" swimtime="00:01:26.93" />
                    <SPLIT distance="150" swimtime="00:02:20.73" />
                    <SPLIT distance="200" swimtime="00:03:20.81" />
                    <SPLIT distance="250" swimtime="00:04:23.37" />
                    <SPLIT distance="300" swimtime="00:05:25.50" />
                    <SPLIT distance="350" swimtime="00:06:10.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="239" reactiontime="+103" swimtime="00:01:18.02" resultid="4050" heatid="7743" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="228" reactiontime="+120" swimtime="00:05:47.82" resultid="4051" heatid="8049" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:16.17" />
                    <SPLIT distance="150" swimtime="00:01:59.68" />
                    <SPLIT distance="200" swimtime="00:02:43.99" />
                    <SPLIT distance="250" swimtime="00:03:29.60" />
                    <SPLIT distance="300" swimtime="00:04:15.66" />
                    <SPLIT distance="350" swimtime="00:05:02.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Piotr" gender="M" lastname="Dąmbski " nation="POL" athleteid="4221">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4222" heatid="7391" lane="1" />
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4223" heatid="7353" lane="4" entrytime="00:00:34.51" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="4224" heatid="7506" lane="6" entrytime="00:01:16.96" />
                <RESULT eventid="1336" status="DNS" swimtime="00:00:00.00" resultid="4225" heatid="7564" lane="2" />
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="4226" heatid="7626" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="4227" heatid="7687" lane="5" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="4228" heatid="7738" lane="3" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Małgorzata " gender="F" lastname="Bogdan" nation="POL" athleteid="4230">
              <RESULTS>
                <RESULT eventid="1285" status="DNS" swimtime="00:00:00.00" resultid="4231" heatid="7530" lane="2" entrytime="00:01:30.00" />
                <RESULT eventid="1319" status="DNS" swimtime="00:00:00.00" resultid="4232" heatid="7562" lane="5" entrytime="00:03:45.00" />
                <RESULT eventid="1419" status="DNS" swimtime="00:00:00.00" resultid="4233" heatid="7617" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="4234" heatid="7652" lane="2" entrytime="00:01:30.00" />
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="4235" heatid="7732" lane="2" entrytime="00:01:40.00" />
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="4236" heatid="7756" lane="4" entrytime="00:03:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Artur" gender="M" lastname="Rutkowski " nation="POL" athleteid="4237">
              <RESULTS>
                <RESULT eventid="1200" points="47" reactiontime="+79" swimtime="00:01:02.47" resultid="4238" heatid="7448" lane="6" entrytime="00:00:38.50" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="4239" heatid="7666" lane="4" entrytime="00:01:18.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Jakub" gender="M" lastname="Rutkowski " nation="POL" athleteid="4240">
              <RESULTS>
                <RESULT eventid="1234" points="488" reactiontime="+92" swimtime="00:02:33.27" resultid="4241" heatid="7485" lane="1" entrytime="00:02:29.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:12.20" />
                    <SPLIT distance="150" swimtime="00:01:51.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="512" reactiontime="+81" swimtime="00:01:09.48" resultid="4242" heatid="7611" lane="6" entrytime="00:01:08.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="498" swimtime="00:00:31.85" resultid="4243" heatid="7812" lane="5" entrytime="00:00:31.14" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Zbigniew" gender="M" lastname="Dymecki" nation="POL" athleteid="4245">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4246" heatid="7392" lane="6" entrytime="00:04:30.00" />
                <RESULT eventid="1302" points="79" reactiontime="+115" swimtime="00:01:58.26" resultid="4248" heatid="7539" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="34" swimtime="00:05:35.60" resultid="4249" heatid="7565" lane="5" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.87" />
                    <SPLIT distance="100" swimtime="00:02:30.26" />
                    <SPLIT distance="150" swimtime="00:04:04.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="75" reactiontime="+121" swimtime="00:03:54.77" resultid="4250" heatid="7688" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                    <SPLIT distance="100" swimtime="00:01:48.06" />
                    <SPLIT distance="150" swimtime="00:02:45.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="58" swimtime="00:10:08.17" resultid="4251" heatid="7975" lane="5" entrytime="00:09:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.71" />
                    <SPLIT distance="100" swimtime="00:02:41.43" />
                    <SPLIT distance="150" swimtime="00:04:06.34" />
                    <SPLIT distance="200" swimtime="00:05:28.40" />
                    <SPLIT distance="250" swimtime="00:06:43.28" />
                    <SPLIT distance="300" swimtime="00:07:59.65" />
                    <SPLIT distance="350" swimtime="00:09:02.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="4252" heatid="7737" lane="4" entrytime="00:02:10.00" />
                <RESULT eventid="1710" points="62" reactiontime="+115" swimtime="00:08:57.35" resultid="4253" heatid="8044" lane="3" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.73" />
                    <SPLIT distance="100" swimtime="00:01:58.19" />
                    <SPLIT distance="150" swimtime="00:03:06.51" />
                    <SPLIT distance="200" swimtime="00:04:15.94" />
                    <SPLIT distance="250" swimtime="00:05:24.88" />
                    <SPLIT distance="300" swimtime="00:06:35.27" />
                    <SPLIT distance="350" swimtime="00:07:47.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="61" reactiontime="+110" swimtime="00:35:57.84" resultid="7936" heatid="7907" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.06" />
                    <SPLIT distance="100" swimtime="00:02:02.75" />
                    <SPLIT distance="150" swimtime="00:03:09.42" />
                    <SPLIT distance="200" swimtime="00:04:18.49" />
                    <SPLIT distance="250" swimtime="00:05:27.90" />
                    <SPLIT distance="300" swimtime="00:06:39.49" />
                    <SPLIT distance="350" swimtime="00:07:49.11" />
                    <SPLIT distance="400" swimtime="00:09:00.20" />
                    <SPLIT distance="450" swimtime="00:10:12.30" />
                    <SPLIT distance="500" swimtime="00:11:21.26" />
                    <SPLIT distance="550" swimtime="00:12:35.26" />
                    <SPLIT distance="600" swimtime="00:13:47.79" />
                    <SPLIT distance="650" swimtime="00:14:59.76" />
                    <SPLIT distance="700" swimtime="00:16:12.86" />
                    <SPLIT distance="750" swimtime="00:17:25.16" />
                    <SPLIT distance="800" swimtime="00:18:38.00" />
                    <SPLIT distance="850" swimtime="00:19:52.22" />
                    <SPLIT distance="900" swimtime="00:21:03.51" />
                    <SPLIT distance="950" swimtime="00:22:17.73" />
                    <SPLIT distance="1000" swimtime="00:23:33.26" />
                    <SPLIT distance="1050" swimtime="00:24:47.76" />
                    <SPLIT distance="1100" swimtime="00:26:03.82" />
                    <SPLIT distance="1150" swimtime="00:27:17.98" />
                    <SPLIT distance="1200" swimtime="00:28:30.15" />
                    <SPLIT distance="1250" swimtime="00:29:44.54" />
                    <SPLIT distance="1300" swimtime="00:31:00.42" />
                    <SPLIT distance="1350" swimtime="00:32:15.19" />
                    <SPLIT distance="1400" swimtime="00:33:28.60" />
                    <SPLIT distance="1450" swimtime="00:34:43.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname=" KATARZYNA" gender="F" lastname="BUBIENKO" nation="POL" athleteid="6124">
              <RESULTS>
                <RESULT eventid="1251" points="217" reactiontime="+113" swimtime="00:01:24.76" resultid="6125" heatid="7492" lane="6" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="99" reactiontime="+129" swimtime="00:04:20.64" resultid="6126" heatid="7561" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.58" />
                    <SPLIT distance="100" swimtime="00:03:15.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="239" reactiontime="+113" swimtime="00:01:40.90" resultid="6127" heatid="7585" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="206" swimtime="00:00:41.26" resultid="6128" heatid="7615" lane="5" entrytime="00:00:41.45" />
                <RESULT eventid="1645" points="246" reactiontime="+106" swimtime="00:00:45.96" resultid="6129" heatid="7782" lane="3" entrytime="00:00:44.81" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-10" firstname="Edward " gender="M" lastname="Dziekoński " nation="POL" athleteid="6130">
              <RESULTS>
                <RESULT eventid="1075" points="134" reactiontime="+105" swimtime="00:00:39.66" resultid="6131" heatid="7351" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1165" points="128" reactiontime="+115" swimtime="00:28:05.66" resultid="6132" heatid="7908" lane="3" entrytime="00:28:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.02" />
                    <SPLIT distance="100" swimtime="00:01:49.82" />
                    <SPLIT distance="150" swimtime="00:02:47.07" />
                    <SPLIT distance="200" swimtime="00:03:44.75" />
                    <SPLIT distance="250" swimtime="00:04:41.60" />
                    <SPLIT distance="300" swimtime="00:05:38.52" />
                    <SPLIT distance="350" swimtime="00:06:34.18" />
                    <SPLIT distance="400" swimtime="00:07:31.38" />
                    <SPLIT distance="450" swimtime="00:08:27.20" />
                    <SPLIT distance="500" swimtime="00:09:23.64" />
                    <SPLIT distance="550" swimtime="00:10:20.62" />
                    <SPLIT distance="600" swimtime="00:11:17.04" />
                    <SPLIT distance="650" swimtime="00:12:13.13" />
                    <SPLIT distance="700" swimtime="00:13:09.04" />
                    <SPLIT distance="750" swimtime="00:14:04.86" />
                    <SPLIT distance="800" swimtime="00:15:00.56" />
                    <SPLIT distance="850" swimtime="00:15:56.01" />
                    <SPLIT distance="900" swimtime="00:16:51.82" />
                    <SPLIT distance="950" swimtime="00:17:47.31" />
                    <SPLIT distance="1000" swimtime="00:18:42.51" />
                    <SPLIT distance="1050" swimtime="00:19:39.59" />
                    <SPLIT distance="1100" swimtime="00:20:36.71" />
                    <SPLIT distance="1150" swimtime="00:21:34.44" />
                    <SPLIT distance="1200" swimtime="00:22:30.25" />
                    <SPLIT distance="1250" swimtime="00:23:28.27" />
                    <SPLIT distance="1300" swimtime="00:24:25.28" />
                    <SPLIT distance="1350" swimtime="00:25:21.13" />
                    <SPLIT distance="1400" swimtime="00:26:17.99" />
                    <SPLIT distance="1450" swimtime="00:27:13.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="130" reactiontime="+107" swimtime="00:01:28.55" resultid="6133" heatid="7503" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="99" swimtime="00:01:49.37" resultid="6134" heatid="7540" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="143" reactiontime="+116" swimtime="00:00:41.63" resultid="6135" heatid="7627" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1504" points="109" swimtime="00:03:27.97" resultid="6136" heatid="7689" lane="5" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.12" />
                    <SPLIT distance="100" swimtime="00:01:37.60" />
                    <SPLIT distance="150" swimtime="00:02:33.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="68" reactiontime="+120" swimtime="00:01:58.32" resultid="6137" heatid="7739" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="118" reactiontime="+114" swimtime="00:07:13.66" resultid="6138" heatid="8045" lane="3" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.34" />
                    <SPLIT distance="100" swimtime="00:01:43.41" />
                    <SPLIT distance="150" swimtime="00:02:40.61" />
                    <SPLIT distance="200" swimtime="00:03:36.26" />
                    <SPLIT distance="250" swimtime="00:04:32.10" />
                    <SPLIT distance="300" swimtime="00:05:27.05" />
                    <SPLIT distance="350" swimtime="00:06:21.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="Sabrina" gender="F" lastname="Staniewska " nation="POL" athleteid="6139">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="6140" heatid="7385" lane="2" entrytime="00:03:15.00" />
                <RESULT eventid="1285" points="276" reactiontime="+105" swimtime="00:01:28.68" resultid="6142" heatid="7530" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="166" swimtime="00:03:39.51" resultid="6143" heatid="7563" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                    <SPLIT distance="100" swimtime="00:01:41.40" />
                    <SPLIT distance="150" swimtime="00:02:05.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="239" reactiontime="+91" swimtime="00:01:28.97" resultid="6144" heatid="7654" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="261" reactiontime="+109" swimtime="00:06:48.31" resultid="6145" heatid="7717" lane="4" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.34" />
                    <SPLIT distance="100" swimtime="00:01:37.86" />
                    <SPLIT distance="150" swimtime="00:02:29.59" />
                    <SPLIT distance="200" swimtime="00:03:20.65" />
                    <SPLIT distance="250" swimtime="00:04:20.28" />
                    <SPLIT distance="300" swimtime="00:05:21.96" />
                    <SPLIT distance="350" swimtime="00:06:05.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="6146" heatid="7759" lane="2" entrytime="00:03:00.00" />
                <RESULT eventid="1693" points="318" reactiontime="+100" swimtime="00:05:43.84" resultid="6147" heatid="8022" lane="4" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:18.20" />
                    <SPLIT distance="150" swimtime="00:02:01.93" />
                    <SPLIT distance="200" swimtime="00:02:46.26" />
                    <SPLIT distance="250" swimtime="00:03:30.67" />
                    <SPLIT distance="300" swimtime="00:04:15.62" />
                    <SPLIT distance="350" swimtime="00:05:00.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="MARIUSZ" gender="M" lastname="GOLON  " nation="POL" athleteid="6148">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="6149" heatid="7368" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1109" points="339" reactiontime="+94" swimtime="00:02:37.87" resultid="6150" heatid="7399" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:02:00.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="352" reactiontime="+77" swimtime="00:00:32.02" resultid="6151" heatid="7452" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1302" points="417" reactiontime="+86" swimtime="00:01:07.90" resultid="6152" heatid="7551" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="431" reactiontime="+83" swimtime="00:00:28.85" resultid="6153" heatid="7639" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="6154" heatid="7667" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="6155" heatid="7743" lane="2" entrytime="00:01:20.00" />
                <RESULT eventid="1662" points="396" reactiontime="+87" swimtime="00:00:34.36" resultid="6156" heatid="7804" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Marcin " gender="M" lastname="Górka" nation="POL" athleteid="6157">
              <RESULTS>
                <RESULT eventid="1200" points="495" swimtime="00:00:28.58" resultid="6158" heatid="7457" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1302" points="447" reactiontime="+79" swimtime="00:01:06.38" resultid="6159" heatid="7557" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="523" reactiontime="+76" swimtime="00:00:27.05" resultid="6160" heatid="7645" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1470" points="453" reactiontime="+58" swimtime="00:01:03.69" resultid="6161" heatid="7673" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="6162" heatid="7750" lane="3" entrytime="00:01:04.00" />
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="6163" heatid="7773" lane="5" entrytime="00:02:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Michał" gender="M" lastname="Gawroński " nation="POL" athleteid="6164">
              <RESULTS>
                <RESULT eventid="1200" points="435" reactiontime="+71" swimtime="00:00:29.84" resultid="6165" heatid="7455" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1302" points="420" reactiontime="+81" swimtime="00:01:07.74" resultid="6166" heatid="7558" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="404" reactiontime="+79" swimtime="00:00:29.48" resultid="6167" heatid="7635" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1662" points="403" reactiontime="+80" swimtime="00:00:34.16" resultid="6168" heatid="7803" lane="4" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Hanna " gender="F" lastname="Kozak " nation="POL" athleteid="6170">
              <RESULTS>
                <RESULT eventid="1453" points="342" reactiontime="+63" swimtime="00:01:18.94" resultid="6172" heatid="7655" lane="4" entrytime="00:01:20.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="325" reactiontime="+65" swimtime="00:02:54.41" resultid="6173" heatid="7760" lane="4" entrytime="00:02:48.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:01:22.55" />
                    <SPLIT distance="150" swimtime="00:02:09.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" status="DNS" swimtime="00:00:00.00" resultid="6174" heatid="7534" lane="1" entrytime="00:01:21.50" />
                <RESULT eventid="1183" points="348" reactiontime="+58" swimtime="00:00:36.52" resultid="7175" heatid="7439" lane="2" entrytime="00:00:36.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Mateusz " gender="M" lastname="Dymiter" nation="POL" athleteid="6183">
              <RESULTS>
                <RESULT eventid="1559" points="305" swimtime="00:05:49.62" resultid="6184" heatid="7979" lane="5" entrytime="00:06:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="150" swimtime="00:02:05.78" />
                    <SPLIT distance="200" swimtime="00:02:52.12" />
                    <SPLIT distance="250" swimtime="00:03:42.07" />
                    <SPLIT distance="300" swimtime="00:04:30.19" />
                    <SPLIT distance="350" swimtime="00:05:09.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="KATARZYNA " gender="F" lastname="MICHAŁOWSKA" nation="POL" athleteid="6446">
              <RESULTS>
                <RESULT eventid="1251" points="286" reactiontime="+107" swimtime="00:01:17.35" resultid="6447" heatid="7494" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="247" reactiontime="+105" swimtime="00:00:38.84" resultid="6448" heatid="7617" lane="6" entrytime="00:00:39.50" />
                <RESULT eventid="1487" status="DNS" swimtime="00:00:00.00" resultid="6449" heatid="7681" lane="6" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Mateusz" gender="M" lastname="Czwartosz " nation="POL" athleteid="7062">
              <RESULTS>
                <RESULT eventid="1200" points="401" reactiontime="+66" swimtime="00:00:30.65" resultid="7063" heatid="7455" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1302" points="419" reactiontime="+83" swimtime="00:01:07.83" resultid="7064" heatid="7557" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="434" swimtime="00:00:28.78" resultid="7065" heatid="7635" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1662" points="435" reactiontime="+79" swimtime="00:00:33.32" resultid="7066" heatid="7803" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Karolina" gender="F" lastname="Kreczmer " nation="POL" athleteid="7317">
              <RESULTS>
                <RESULT eventid="1183" status="DNS" swimtime="00:00:00.00" resultid="7318" heatid="7438" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="7319" heatid="7494" lane="1" entrytime="00:01:15.00" />
                <RESULT eventid="1285" status="DNS" swimtime="00:00:00.00" resultid="7320" heatid="7533" lane="2" entrytime="00:01:25.00" />
                <RESULT eventid="1419" status="DNS" swimtime="00:00:00.00" resultid="7321" heatid="7617" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="7322" heatid="7654" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="7323" heatid="7758" lane="5" entrytime="00:03:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Zofia" gender="F" lastname="Brunka" nation="POL" athleteid="7324">
              <RESULTS>
                <RESULT eventid="1183" points="282" reactiontime="+66" swimtime="00:00:39.18" resultid="7325" heatid="7437" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="7326" heatid="7494" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1285" points="289" swimtime="00:01:27.24" resultid="7327" heatid="7533" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="286" reactiontime="+75" swimtime="00:00:36.99" resultid="7328" heatid="7617" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="7329" heatid="7655" lane="6" entrytime="00:01:24.00" />
                <RESULT eventid="1611" points="255" reactiontime="+66" swimtime="00:03:09.10" resultid="7330" heatid="7758" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:30.28" />
                    <SPLIT distance="150" swimtime="00:02:19.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="MOSiR KSZO Ostrowiec" nation="POL">
          <CONTACT name="Różalski" street="Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" athleteid="2403">
              <RESULTS>
                <RESULT eventid="1075" points="262" reactiontime="+78" swimtime="00:00:31.71" resultid="2404" heatid="7357" lane="3" entrytime="00:00:32.50" />
                <RESULT eventid="1109" points="162" reactiontime="+100" swimtime="00:03:21.93" resultid="2405" heatid="7395" lane="4" entrytime="00:03:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:38.23" />
                    <SPLIT distance="150" swimtime="00:02:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="223" reactiontime="+91" swimtime="00:01:23.59" resultid="2406" heatid="7544" lane="4" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="105" reactiontime="+107" swimtime="00:03:50.98" resultid="2407" heatid="7566" lane="2" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.35" />
                    <SPLIT distance="100" swimtime="00:01:50.02" />
                    <SPLIT distance="150" swimtime="00:02:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="227" reactiontime="+93" swimtime="00:00:35.71" resultid="2408" heatid="7631" lane="4" entrytime="00:00:34.80" />
                <RESULT eventid="1559" points="144" reactiontime="+102" swimtime="00:07:28.49" resultid="2409" heatid="7976" lane="4" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.80" />
                    <SPLIT distance="100" swimtime="00:01:47.74" />
                    <SPLIT distance="150" swimtime="00:02:47.29" />
                    <SPLIT distance="200" swimtime="00:03:46.11" />
                    <SPLIT distance="250" swimtime="00:04:49.85" />
                    <SPLIT distance="300" swimtime="00:05:53.06" />
                    <SPLIT distance="350" swimtime="00:06:42.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="121" reactiontime="+102" swimtime="00:01:37.75" resultid="2410" heatid="7740" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="217" swimtime="00:00:42.00" resultid="2411" heatid="7795" lane="5" entrytime="00:00:42.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="MOSiR Częstochowa" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1969-01-01" firstname="Ireneusz " gender="M" lastname="Stachurski" nation="POL" athleteid="2413">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="2414" heatid="7350" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="2416" heatid="7690" lane="2" entrytime="00:03:00.00" />
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="2417" heatid="8047" lane="5" entrytime="00:06:30.00" />
                <RESULT eventid="1470" points="121" reactiontime="+86" swimtime="00:01:38.78" resultid="2634" heatid="7662" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="2635" heatid="7765" lane="6" entrytime="00:03:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00811" name="Pałac Katowice Masters" nation="POL" region="11">
          <CONTACT email="tsplywak@wp.pl" name="Bucholz" phone="606 135 860" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-26" firstname="Tomasz" gender="M" lastname="Bucholz" nation="POL" athleteid="2419" />
            <ATHLETE birthdate="1973-11-03" firstname="Sławomir" gender="M" lastname="Szafarczyk" nation="POL" athleteid="2420" />
            <ATHLETE birthdate="1973-08-28" firstname="Jacek" gender="M" lastname="Kobylczak" nation="POL" athleteid="2422" />
            <ATHLETE birthdate="1972-01-01" firstname="Matysiewicz" gender="M" lastname="Mateusz" nation="POL" athleteid="7947" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="298" reactiontime="+62" swimtime="00:02:17.38" resultid="7162" heatid="7932" lane="5" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="150" swimtime="00:01:47.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2420" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="2422" number="2" />
                    <RELAYPOSITION athleteid="7947" number="3" />
                    <RELAYPOSITION athleteid="2419" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1528" points="302" reactiontime="+83" swimtime="00:02:00.35" resultid="2423" heatid="7711" lane="3" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                    <SPLIT distance="100" swimtime="00:00:52.41" />
                    <SPLIT distance="150" swimtime="00:01:30.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2420" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="7947" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2419" number="3" />
                    <RELAYPOSITION athleteid="2422" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="HTF" name="Happy Tri Friends" nation="POL" region="KR">
          <CONTACT city="Kraków" email="m-lewandowski@o2.pl" name="Lewandowski Marcin" phone="501486298" state="MAŁOP" street="Twardowskiego 37" zip="30-312" />
          <ATHLETES>
            <ATHLETE birthdate="1973-04-13" firstname="Marcin" gender="M" lastname="Lewandowski" nation="POL" license="ML" athleteid="2450">
              <RESULTS>
                <RESULT eventid="1165" points="308" reactiontime="+96" swimtime="00:20:58.05" resultid="2451" heatid="7915" lane="2" entrytime="00:20:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:17.98" />
                    <SPLIT distance="150" swimtime="00:01:58.69" />
                    <SPLIT distance="200" swimtime="00:02:39.42" />
                    <SPLIT distance="250" swimtime="00:03:20.92" />
                    <SPLIT distance="300" swimtime="00:04:02.35" />
                    <SPLIT distance="350" swimtime="00:04:44.07" />
                    <SPLIT distance="400" swimtime="00:05:26.00" />
                    <SPLIT distance="450" swimtime="00:06:07.62" />
                    <SPLIT distance="500" swimtime="00:06:49.41" />
                    <SPLIT distance="550" swimtime="00:07:31.37" />
                    <SPLIT distance="600" swimtime="00:08:13.12" />
                    <SPLIT distance="650" swimtime="00:08:55.32" />
                    <SPLIT distance="700" swimtime="00:09:37.64" />
                    <SPLIT distance="750" swimtime="00:10:20.10" />
                    <SPLIT distance="800" swimtime="00:11:02.30" />
                    <SPLIT distance="850" swimtime="00:11:44.82" />
                    <SPLIT distance="900" swimtime="00:12:26.95" />
                    <SPLIT distance="950" swimtime="00:13:09.27" />
                    <SPLIT distance="1000" swimtime="00:13:51.44" />
                    <SPLIT distance="1050" swimtime="00:14:33.77" />
                    <SPLIT distance="1100" swimtime="00:15:16.33" />
                    <SPLIT distance="1150" swimtime="00:15:59.14" />
                    <SPLIT distance="1200" swimtime="00:16:41.97" />
                    <SPLIT distance="1250" swimtime="00:17:24.57" />
                    <SPLIT distance="1300" swimtime="00:18:07.77" />
                    <SPLIT distance="1350" swimtime="00:18:50.64" />
                    <SPLIT distance="1400" swimtime="00:19:33.25" />
                    <SPLIT distance="1450" swimtime="00:20:16.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="328" reactiontime="+83" swimtime="00:02:24.03" resultid="2452" heatid="7700" lane="2" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:46.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="325" reactiontime="+91" swimtime="00:05:09.30" resultid="2453" heatid="8053" lane="4" entrytime="00:05:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="150" swimtime="00:01:51.27" />
                    <SPLIT distance="200" swimtime="00:02:30.09" />
                    <SPLIT distance="250" swimtime="00:03:09.70" />
                    <SPLIT distance="300" swimtime="00:03:49.65" />
                    <SPLIT distance="350" swimtime="00:04:29.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01511" name="MTP Delfin Cieszyn" nation="POL" region="11">
          <ATHLETES>
            <ATHLETE birthdate="1986-05-25" firstname="Łukasz" gender="M" lastname="Widzik" nation="POL" athleteid="6175">
              <RESULTS>
                <RESULT eventid="1165" points="410" swimtime="00:19:04.19" resultid="6176" heatid="7907" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:07.33" />
                    <SPLIT distance="150" swimtime="00:01:44.51" />
                    <SPLIT distance="200" swimtime="00:02:21.73" />
                    <SPLIT distance="250" swimtime="00:02:59.60" />
                    <SPLIT distance="300" swimtime="00:03:37.50" />
                    <SPLIT distance="350" swimtime="00:04:15.01" />
                    <SPLIT distance="400" swimtime="00:04:52.85" />
                    <SPLIT distance="450" swimtime="00:05:30.89" />
                    <SPLIT distance="500" swimtime="00:06:09.43" />
                    <SPLIT distance="550" swimtime="00:06:47.75" />
                    <SPLIT distance="600" swimtime="00:07:26.37" />
                    <SPLIT distance="650" swimtime="00:08:04.94" />
                    <SPLIT distance="700" swimtime="00:08:43.73" />
                    <SPLIT distance="750" swimtime="00:09:22.61" />
                    <SPLIT distance="800" swimtime="00:10:01.93" />
                    <SPLIT distance="850" swimtime="00:10:40.97" />
                    <SPLIT distance="900" swimtime="00:11:20.51" />
                    <SPLIT distance="950" swimtime="00:11:59.56" />
                    <SPLIT distance="1000" swimtime="00:12:38.68" />
                    <SPLIT distance="1050" swimtime="00:13:17.75" />
                    <SPLIT distance="1100" swimtime="00:13:56.54" />
                    <SPLIT distance="1150" swimtime="00:14:36.05" />
                    <SPLIT distance="1200" swimtime="00:15:15.57" />
                    <SPLIT distance="1250" swimtime="00:15:54.22" />
                    <SPLIT distance="1300" swimtime="00:16:33.14" />
                    <SPLIT distance="1350" swimtime="00:17:12.16" />
                    <SPLIT distance="1400" swimtime="00:17:50.59" />
                    <SPLIT distance="1450" swimtime="00:18:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="6177" heatid="7673" lane="5" entrytime="00:01:03.78" />
                <RESULT eventid="1504" points="412" reactiontime="+73" swimtime="00:02:13.46" resultid="6178" heatid="7686" lane="6" entrytime="00:02:09.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                    <SPLIT distance="100" swimtime="00:01:03.09" />
                    <SPLIT distance="150" swimtime="00:01:38.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="6179" heatid="7773" lane="3" entrytime="00:02:19.76" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-16" firstname="Dominika" gender="F" lastname="Będlin" nation="POL" athleteid="6180">
              <RESULTS>
                <RESULT eventid="1058" points="192" reactiontime="+129" swimtime="00:00:40.30" resultid="6181" heatid="7331" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="6287" heatid="7496" lane="5" entrytime="00:01:08.00" />
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="6473" heatid="7591" lane="2" entrytime="00:01:20.70" />
                <RESULT eventid="1645" points="99" reactiontime="+116" swimtime="00:01:02.10" resultid="6474" heatid="7775" lane="6" entrytime="00:00:38.21" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="GöteborgSim" nation="SWE">
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Leonard" gender="M" lastname="Bielicz" nation="POL" athleteid="2465">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1075" points="414" reactiontime="+73" swimtime="00:00:27.23" resultid="2466" heatid="7375" lane="1" entrytime="00:00:26.80" />
                <RESULT comment="Rekord Polski Masters" eventid="1268" points="393" swimtime="00:01:01.35" resultid="2467" heatid="7519" lane="5" entrytime="00:01:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1302" points="357" reactiontime="+74" swimtime="00:01:11.53" resultid="2468" heatid="7550" lane="4" entrytime="00:01:13.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1436" points="399" reactiontime="+79" swimtime="00:00:29.59" resultid="2469" heatid="7641" lane="4" entrytime="00:00:29.06" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="2470" heatid="7751" lane="5" entrytime="00:01:07.37" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="VSK Slávia PF České Budějovice" nation="CZE">
          <ATHLETES>
            <ATHLETE birthdate="1956-08-31" firstname="Petr " gender="M" lastname="Ries" nation="CZE" athleteid="2483">
              <RESULTS>
                <RESULT eventid="1268" points="222" reactiontime="+87" swimtime="00:01:14.14" resultid="2484" heatid="7507" lane="3" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Iks Konstancin" nation="POL">
          <CONTACT name="Juchno" />
          <ATHLETES>
            <ATHLETE birthdate="1969-01-01" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" athleteid="2487">
              <RESULTS>
                <RESULT eventid="1075" points="410" reactiontime="+74" swimtime="00:00:27.31" resultid="2488" heatid="7372" lane="2" entrytime="00:00:27.50" />
                <RESULT eventid="1109" points="336" swimtime="00:02:38.26" resultid="2489" heatid="7400" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                    <SPLIT distance="150" swimtime="00:02:02.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="426" swimtime="00:00:59.70" resultid="2490" heatid="7520" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="342" reactiontime="+79" swimtime="00:01:12.58" resultid="2491" heatid="7549" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="2492" heatid="7606" lane="6" entrytime="00:01:21.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="2493" heatid="7701" lane="3" entrytime="00:02:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-03" firstname="Rafal" gender="M" lastname="Juchno" nation="POL" athleteid="6419">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="6420" heatid="7366" lane="6" entrytime="00:00:29.30" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="6421" heatid="7515" lane="6" entrytime="00:01:05.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="6422" heatid="7600" lane="2" entrytime="00:01:30.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="6423" heatid="7694" lane="6" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01711" name="UKS WODNIK Sieminanowice Śląskie" nation="POL" region="11" shortname="UKS WODNIK Sieminanowice Śląsk">
          <CONTACT city="Siemianowice Śląskie" email="vivisektor@interia.pl" name="Małyszek Leszek" phone="534039934" state="ŚLĄSK" street="Mikołaja 3" zip="41-106" />
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="2495">
              <RESULTS>
                <RESULT eventid="1109" points="229" reactiontime="+85" swimtime="00:02:59.75" resultid="2496" heatid="7397" lane="4" entrytime="00:02:55.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:25.20" />
                    <SPLIT distance="150" swimtime="00:02:17.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="276" swimtime="00:21:45.25" resultid="2497" heatid="7914" lane="5" entrytime="00:21:14.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                    <SPLIT distance="100" swimtime="00:01:19.75" />
                    <SPLIT distance="150" swimtime="00:02:02.94" />
                    <SPLIT distance="200" swimtime="00:02:46.18" />
                    <SPLIT distance="250" swimtime="00:03:29.32" />
                    <SPLIT distance="300" swimtime="00:04:13.46" />
                    <SPLIT distance="350" swimtime="00:04:57.42" />
                    <SPLIT distance="400" swimtime="00:05:42.15" />
                    <SPLIT distance="450" swimtime="00:06:26.62" />
                    <SPLIT distance="500" swimtime="00:07:10.45" />
                    <SPLIT distance="550" swimtime="00:07:54.56" />
                    <SPLIT distance="600" swimtime="00:08:38.65" />
                    <SPLIT distance="650" swimtime="00:09:22.72" />
                    <SPLIT distance="700" swimtime="00:10:06.98" />
                    <SPLIT distance="750" swimtime="00:10:51.01" />
                    <SPLIT distance="800" swimtime="00:11:34.79" />
                    <SPLIT distance="850" swimtime="00:12:18.90" />
                    <SPLIT distance="900" swimtime="00:13:02.65" />
                    <SPLIT distance="950" swimtime="00:13:46.55" />
                    <SPLIT distance="1000" swimtime="00:14:30.77" />
                    <SPLIT distance="1050" swimtime="00:15:14.55" />
                    <SPLIT distance="1100" swimtime="00:15:58.63" />
                    <SPLIT distance="1150" swimtime="00:16:42.23" />
                    <SPLIT distance="1200" swimtime="00:17:26.20" />
                    <SPLIT distance="1250" swimtime="00:18:09.86" />
                    <SPLIT distance="1300" swimtime="00:18:53.62" />
                    <SPLIT distance="1350" swimtime="00:19:38.25" />
                    <SPLIT distance="1400" swimtime="00:20:20.88" />
                    <SPLIT distance="1450" swimtime="00:21:04.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="218" reactiontime="+77" swimtime="00:00:36.21" resultid="2498" heatid="7630" lane="6" entrytime="00:00:35.20" />
                <RESULT eventid="1559" points="208" reactiontime="+86" swimtime="00:06:37.38" resultid="2499" heatid="7978" lane="4" entrytime="00:06:22.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                    <SPLIT distance="100" swimtime="00:01:38.36" />
                    <SPLIT distance="150" swimtime="00:02:30.99" />
                    <SPLIT distance="200" swimtime="00:03:21.29" />
                    <SPLIT distance="250" swimtime="00:04:17.28" />
                    <SPLIT distance="300" swimtime="00:05:13.01" />
                    <SPLIT distance="350" swimtime="00:05:55.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="256" reactiontime="+86" swimtime="00:05:34.85" resultid="2500" heatid="8051" lane="1" entrytime="00:05:35.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:01:19.92" />
                    <SPLIT distance="150" swimtime="00:02:02.31" />
                    <SPLIT distance="200" swimtime="00:02:44.53" />
                    <SPLIT distance="250" swimtime="00:03:26.98" />
                    <SPLIT distance="300" swimtime="00:04:09.66" />
                    <SPLIT distance="350" swimtime="00:04:52.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="CityZen Poznań" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Marcin " gender="M" lastname="Jabłoński" nation="POL" athleteid="2502">
              <RESULTS>
                <RESULT eventid="1075" points="582" reactiontime="+68" swimtime="00:00:24.31" resultid="2503" heatid="7381" lane="4" entrytime="00:00:23.42" />
                <RESULT eventid="1109" points="561" reactiontime="+71" swimtime="00:02:13.44" resultid="2504" heatid="7407" lane="4" entrytime="00:02:08.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="100" swimtime="00:01:02.19" />
                    <SPLIT distance="150" swimtime="00:01:41.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="532" reactiontime="+56" swimtime="00:00:27.89" resultid="2505" heatid="7460" lane="5" entrytime="00:00:27.02" />
                <RESULT eventid="1268" points="630" reactiontime="+70" swimtime="00:00:52.41" resultid="2506" heatid="7525" lane="3" entrytime="00:00:50.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="603" swimtime="00:00:25.79" resultid="2507" heatid="7647" lane="5" entrytime="00:00:25.21" />
                <RESULT eventid="1504" points="609" reactiontime="+73" swimtime="00:01:57.17" resultid="2508" heatid="7706" lane="4" entrytime="00:01:52.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                    <SPLIT distance="100" swimtime="00:00:57.13" />
                    <SPLIT distance="150" swimtime="00:01:28.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="635" reactiontime="+71" swimtime="00:00:56.39" resultid="2509" heatid="7752" lane="4" entrytime="00:00:55.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="556" reactiontime="+71" swimtime="00:04:18.70" resultid="2510" heatid="8058" lane="4" entrytime="00:04:05.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                    <SPLIT distance="100" swimtime="00:00:59.22" />
                    <SPLIT distance="150" swimtime="00:01:31.65" />
                    <SPLIT distance="200" swimtime="00:02:04.22" />
                    <SPLIT distance="250" swimtime="00:02:37.43" />
                    <SPLIT distance="300" swimtime="00:03:11.17" />
                    <SPLIT distance="350" swimtime="00:03:44.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KUPI" name="Športový plavecký klub Kúpele Piešťany " nation="SVK">
          <ATHLETES>
            <ATHLETE birthdate="1961-04-20" firstname="Anna " gender="F" lastname="Kičínová" nation="SVK" athleteid="2512">
              <RESULTS>
                <RESULT eventid="1645" points="280" reactiontime="+100" swimtime="00:00:44.00" resultid="2515" heatid="7783" lane="6" entrytime="00:00:44.40" />
                <RESULT eventid="1385" points="278" reactiontime="+99" swimtime="00:01:36.06" resultid="2516" heatid="7587" lane="4" entrytime="00:01:37.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="270" reactiontime="+91" swimtime="00:03:27.96" resultid="2517" heatid="7466" lane="4" entrytime="00:03:29.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                    <SPLIT distance="100" swimtime="00:01:36.77" />
                    <SPLIT distance="150" swimtime="00:02:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="227" reactiontime="+95" swimtime="00:00:39.96" resultid="2518" heatid="7615" lane="3" entrytime="00:00:40.30" />
                <RESULT eventid="1577" points="251" reactiontime="+99" swimtime="00:01:27.24" resultid="2519" heatid="7733" lane="6" entrytime="00:01:32.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="239" reactiontime="+101" swimtime="00:03:14.60" resultid="2520" heatid="7563" lane="6" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:01:30.97" />
                    <SPLIT distance="150" swimtime="00:02:22.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-10-27" firstname="Pavol " gender="M" lastname="Škodný" nation="SVK" athleteid="2513">
              <RESULTS>
                <RESULT eventid="1470" points="321" reactiontime="+71" swimtime="00:01:11.46" resultid="2521" heatid="7669" lane="3" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="311" reactiontime="+73" swimtime="00:02:36.60" resultid="2522" heatid="7771" lane="4" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:16.65" />
                    <SPLIT distance="150" swimtime="00:01:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="347" reactiontime="+94" swimtime="00:05:35.13" resultid="2523" heatid="7980" lane="2" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:16.50" />
                    <SPLIT distance="150" swimtime="00:01:59.41" />
                    <SPLIT distance="200" swimtime="00:02:41.62" />
                    <SPLIT distance="250" swimtime="00:03:31.19" />
                    <SPLIT distance="300" swimtime="00:04:20.50" />
                    <SPLIT distance="350" swimtime="00:04:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="326" swimtime="00:05:09.04" resultid="2524" heatid="8054" lane="5" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="150" swimtime="00:01:49.67" />
                    <SPLIT distance="200" swimtime="00:02:29.65" />
                    <SPLIT distance="250" swimtime="00:03:09.90" />
                    <SPLIT distance="300" swimtime="00:03:50.45" />
                    <SPLIT distance="350" swimtime="00:04:30.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-15" firstname="Lucia " gender="F" lastname="Vachanová" nation="SVK" athleteid="2514">
              <RESULTS>
                <RESULT eventid="1183" points="420" reactiontime="+70" swimtime="00:00:34.31" resultid="2525" heatid="7439" lane="6" entrytime="00:00:36.90" />
                <RESULT eventid="1453" points="411" reactiontime="+75" swimtime="00:01:14.28" resultid="2526" heatid="7656" lane="2" entrytime="00:01:19.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="395" reactiontime="+75" swimtime="00:02:43.48" resultid="2527" heatid="7760" lane="2" entrytime="00:02:49.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:19.86" />
                    <SPLIT distance="150" swimtime="00:02:02.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="436" reactiontime="+79" swimtime="00:01:07.27" resultid="2528" heatid="7496" lane="1" entrytime="00:01:08.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="496" reactiontime="+93" swimtime="00:02:20.39" resultid="2529" heatid="7683" lane="2" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:09.05" />
                    <SPLIT distance="150" swimtime="00:01:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="465" reactiontime="+91" swimtime="00:05:03.03" resultid="2530" heatid="8024" lane="1" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:11.39" />
                    <SPLIT distance="150" swimtime="00:01:49.64" />
                    <SPLIT distance="200" swimtime="00:02:28.41" />
                    <SPLIT distance="250" swimtime="00:03:07.15" />
                    <SPLIT distance="300" swimtime="00:03:45.88" />
                    <SPLIT distance="350" swimtime="00:04:25.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WARPOZ" name="KS Warta Poznań" nation="POL" region="WIE">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Thiem Jacek" phone="502499565" state="WIE" street="Os. Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1982-05-14" firstname="Przemysław" gender="M" lastname="Isalski" nation="POL" license="50011520013" athleteid="2541">
              <RESULTS>
                <RESULT eventid="1109" points="441" reactiontime="+81" swimtime="00:02:24.52" resultid="2542" heatid="7401" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="100" swimtime="00:01:07.70" />
                    <SPLIT distance="150" swimtime="00:01:49.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="460" reactiontime="+85" swimtime="00:18:20.95" resultid="2543" heatid="7917" lane="6" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:07.01" />
                    <SPLIT distance="150" swimtime="00:01:42.72" />
                    <SPLIT distance="200" swimtime="00:02:18.69" />
                    <SPLIT distance="250" swimtime="00:02:54.82" />
                    <SPLIT distance="300" swimtime="00:03:30.84" />
                    <SPLIT distance="350" swimtime="00:04:06.43" />
                    <SPLIT distance="400" swimtime="00:04:42.45" />
                    <SPLIT distance="450" swimtime="00:05:18.48" />
                    <SPLIT distance="500" swimtime="00:05:54.61" />
                    <SPLIT distance="550" swimtime="00:06:31.11" />
                    <SPLIT distance="600" swimtime="00:07:07.64" />
                    <SPLIT distance="650" swimtime="00:07:44.34" />
                    <SPLIT distance="700" swimtime="00:08:21.04" />
                    <SPLIT distance="750" swimtime="00:08:58.01" />
                    <SPLIT distance="800" swimtime="00:09:35.30" />
                    <SPLIT distance="850" swimtime="00:10:12.67" />
                    <SPLIT distance="900" swimtime="00:10:49.88" />
                    <SPLIT distance="950" swimtime="00:11:27.84" />
                    <SPLIT distance="1000" swimtime="00:12:06.12" />
                    <SPLIT distance="1050" swimtime="00:12:44.38" />
                    <SPLIT distance="1100" swimtime="00:13:22.06" />
                    <SPLIT distance="1150" swimtime="00:14:00.59" />
                    <SPLIT distance="1200" swimtime="00:14:38.20" />
                    <SPLIT distance="1250" swimtime="00:15:15.60" />
                    <SPLIT distance="1300" swimtime="00:15:52.89" />
                    <SPLIT distance="1350" swimtime="00:16:30.21" />
                    <SPLIT distance="1400" swimtime="00:17:07.51" />
                    <SPLIT distance="1450" swimtime="00:17:44.30" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K-14 - Dotkniecie ściany jedną ręka przy nawrocie" eventid="1234" reactiontime="+83" status="DSQ" swimtime="00:02:43.40" resultid="2544" heatid="7480" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:18.29" />
                    <SPLIT distance="150" swimtime="00:02:00.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="438" swimtime="00:01:06.80" resultid="2545" heatid="7551" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="476" swimtime="00:02:07.22" resultid="2546" heatid="7703" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="100" swimtime="00:01:01.83" />
                    <SPLIT distance="150" swimtime="00:01:34.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="427" reactiontime="+83" swimtime="00:05:12.56" resultid="2547" heatid="7982" lane="2" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:11.11" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                    <SPLIT distance="200" swimtime="00:02:34.17" />
                    <SPLIT distance="250" swimtime="00:03:18.85" />
                    <SPLIT distance="300" swimtime="00:04:04.00" />
                    <SPLIT distance="350" swimtime="00:04:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="293" reactiontime="+87" swimtime="00:01:12.91" resultid="2548" heatid="7746" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="481" reactiontime="+84" swimtime="00:04:31.49" resultid="2549" heatid="8056" lane="1" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:40.89" />
                    <SPLIT distance="200" swimtime="00:02:15.36" />
                    <SPLIT distance="250" swimtime="00:02:49.61" />
                    <SPLIT distance="300" swimtime="00:03:23.48" />
                    <SPLIT distance="350" swimtime="00:03:57.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-04-19" firstname="Marek" gender="M" lastname="Stanoch" nation="POL" athleteid="2550">
              <RESULTS>
                <RESULT eventid="1075" points="207" reactiontime="+99" swimtime="00:00:34.31" resultid="2551" heatid="7364" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1302" points="152" reactiontime="+96" swimtime="00:01:34.98" resultid="2552" heatid="7545" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="186" reactiontime="+98" swimtime="00:01:37.39" resultid="2553" heatid="7601" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="219" reactiontime="+87" swimtime="00:00:41.84" resultid="2554" heatid="7802" lane="6" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-05-19" firstname="Jakub" gender="M" lastname="Stanoch" nation="POL" license="50011520014" athleteid="2555">
              <RESULTS>
                <RESULT eventid="1165" points="399" reactiontime="+73" swimtime="00:19:14.30" resultid="2556" heatid="7914" lane="4" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:08.10" />
                    <SPLIT distance="150" swimtime="00:01:45.14" />
                    <SPLIT distance="200" swimtime="00:02:23.06" />
                    <SPLIT distance="250" swimtime="00:03:01.31" />
                    <SPLIT distance="300" swimtime="00:03:39.64" />
                    <SPLIT distance="350" swimtime="00:04:18.04" />
                    <SPLIT distance="400" swimtime="00:04:56.55" />
                    <SPLIT distance="450" swimtime="00:05:35.45" />
                    <SPLIT distance="500" swimtime="00:06:14.29" />
                    <SPLIT distance="550" swimtime="00:06:52.66" />
                    <SPLIT distance="600" swimtime="00:07:31.50" />
                    <SPLIT distance="650" swimtime="00:08:10.83" />
                    <SPLIT distance="700" swimtime="00:08:49.55" />
                    <SPLIT distance="750" swimtime="00:09:28.28" />
                    <SPLIT distance="800" swimtime="00:10:07.27" />
                    <SPLIT distance="850" swimtime="00:10:45.93" />
                    <SPLIT distance="900" swimtime="00:11:24.96" />
                    <SPLIT distance="950" swimtime="00:12:04.00" />
                    <SPLIT distance="1000" swimtime="00:12:42.91" />
                    <SPLIT distance="1050" swimtime="00:13:21.60" />
                    <SPLIT distance="1100" swimtime="00:14:00.85" />
                    <SPLIT distance="1150" swimtime="00:14:40.68" />
                    <SPLIT distance="1200" swimtime="00:15:19.85" />
                    <SPLIT distance="1250" swimtime="00:15:59.20" />
                    <SPLIT distance="1300" swimtime="00:16:38.40" />
                    <SPLIT distance="1350" swimtime="00:17:17.65" />
                    <SPLIT distance="1400" swimtime="00:17:56.82" />
                    <SPLIT distance="1450" swimtime="00:18:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="370" reactiontime="+67" swimtime="00:02:31.85" resultid="2557" heatid="7570" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:10.34" />
                    <SPLIT distance="150" swimtime="00:01:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="460" reactiontime="+68" swimtime="00:00:28.22" resultid="2558" heatid="7644" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1594" points="431" reactiontime="+70" swimtime="00:01:04.18" resultid="2559" heatid="7749" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="403" reactiontime="+68" swimtime="00:04:47.85" resultid="2560" heatid="8055" lane="1" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                    <SPLIT distance="150" swimtime="00:01:40.25" />
                    <SPLIT distance="200" swimtime="00:02:16.87" />
                    <SPLIT distance="250" swimtime="00:02:54.18" />
                    <SPLIT distance="300" swimtime="00:03:32.58" />
                    <SPLIT distance="350" swimtime="00:04:10.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="Tomaszewski" nation="POL" athleteid="2561">
              <RESULTS>
                <RESULT eventid="1075" points="449" swimtime="00:00:26.51" resultid="2562" heatid="7372" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="1200" points="449" reactiontime="+69" swimtime="00:00:29.51" resultid="2563" heatid="7457" lane="1" entrytime="00:00:30.30" />
                <RESULT eventid="1470" points="452" reactiontime="+70" swimtime="00:01:03.73" resultid="2564" heatid="7670" lane="3" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="2565" heatid="7697" lane="4" entrytime="00:02:26.00" />
                <RESULT eventid="1628" points="394" reactiontime="+72" swimtime="00:02:24.74" resultid="2566" heatid="7771" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Rusłana" gender="F" lastname="Dembecka" nation="POL" athleteid="2567">
              <RESULTS>
                <RESULT eventid="1217" points="137" reactiontime="+126" swimtime="00:04:20.52" resultid="2568" heatid="7463" lane="1" entrytime="00:04:46.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.02" />
                    <SPLIT distance="100" swimtime="00:02:13.26" />
                    <SPLIT distance="150" swimtime="00:03:18.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="135" reactiontime="+116" swimtime="00:02:02.06" resultid="2569" heatid="7584" lane="6" entrytime="00:02:01.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="155" reactiontime="+104" swimtime="00:00:53.50" resultid="2570" heatid="7778" lane="4" entrytime="00:00:53.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="50011520005" athleteid="2571">
              <RESULTS>
                <RESULT eventid="1075" points="243" reactiontime="+92" swimtime="00:00:32.49" resultid="2572" heatid="7357" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="1165" points="212" reactiontime="+118" swimtime="00:23:45.11" resultid="2573" heatid="7910" lane="2" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                    <SPLIT distance="100" swimtime="00:01:28.53" />
                    <SPLIT distance="150" swimtime="00:02:15.33" />
                    <SPLIT distance="200" swimtime="00:03:03.18" />
                    <SPLIT distance="250" swimtime="00:03:51.25" />
                    <SPLIT distance="300" swimtime="00:04:39.43" />
                    <SPLIT distance="350" swimtime="00:05:27.90" />
                    <SPLIT distance="400" swimtime="00:06:16.44" />
                    <SPLIT distance="450" swimtime="00:07:05.00" />
                    <SPLIT distance="500" swimtime="00:07:53.65" />
                    <SPLIT distance="550" swimtime="00:08:42.39" />
                    <SPLIT distance="600" swimtime="00:09:30.84" />
                    <SPLIT distance="650" swimtime="00:10:18.97" />
                    <SPLIT distance="700" swimtime="00:11:07.82" />
                    <SPLIT distance="750" swimtime="00:11:56.53" />
                    <SPLIT distance="800" swimtime="00:12:45.07" />
                    <SPLIT distance="850" swimtime="00:13:33.99" />
                    <SPLIT distance="900" swimtime="00:14:21.83" />
                    <SPLIT distance="950" swimtime="00:15:09.99" />
                    <SPLIT distance="1000" swimtime="00:15:58.40" />
                    <SPLIT distance="1050" swimtime="00:16:46.63" />
                    <SPLIT distance="1100" swimtime="00:17:34.05" />
                    <SPLIT distance="1150" swimtime="00:18:22.13" />
                    <SPLIT distance="1200" swimtime="00:19:10.06" />
                    <SPLIT distance="1250" swimtime="00:19:57.67" />
                    <SPLIT distance="1300" swimtime="00:20:44.98" />
                    <SPLIT distance="1350" swimtime="00:21:31.70" />
                    <SPLIT distance="1400" swimtime="00:22:17.82" />
                    <SPLIT distance="1450" swimtime="00:23:03.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="191" swimtime="00:03:09.19" resultid="2574" heatid="7568" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:31.07" />
                    <SPLIT distance="150" swimtime="00:02:19.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="216" reactiontime="+109" swimtime="00:02:45.48" resultid="2575" heatid="7693" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:22.92" />
                    <SPLIT distance="150" swimtime="00:02:05.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="168" reactiontime="+113" swimtime="00:07:06.53" resultid="2576" heatid="7977" lane="3" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:38.07" />
                    <SPLIT distance="150" swimtime="00:03:35.77" />
                    <SPLIT distance="200" swimtime="00:04:34.81" />
                    <SPLIT distance="250" swimtime="00:05:33.04" />
                    <SPLIT distance="300" swimtime="00:06:20.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="174" reactiontime="+108" swimtime="00:01:26.71" resultid="2577" heatid="7741" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="205" reactiontime="+111" swimtime="00:06:00.84" resultid="2578" heatid="8049" lane="3" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:26.58" />
                    <SPLIT distance="150" swimtime="00:02:12.96" />
                    <SPLIT distance="200" swimtime="00:02:59.95" />
                    <SPLIT distance="250" swimtime="00:03:46.11" />
                    <SPLIT distance="300" swimtime="00:04:33.26" />
                    <SPLIT distance="350" swimtime="00:05:18.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" license="50011520006" athleteid="2579">
              <RESULTS>
                <RESULT eventid="1165" points="322" reactiontime="+99" swimtime="00:20:40.19" resultid="2580" heatid="7915" lane="1" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:01:16.93" />
                    <SPLIT distance="150" swimtime="00:01:57.83" />
                    <SPLIT distance="200" swimtime="00:02:38.98" />
                    <SPLIT distance="250" swimtime="00:03:20.92" />
                    <SPLIT distance="300" swimtime="00:04:02.10" />
                    <SPLIT distance="350" swimtime="00:04:44.13" />
                    <SPLIT distance="400" swimtime="00:05:25.75" />
                    <SPLIT distance="450" swimtime="00:06:07.26" />
                    <SPLIT distance="500" swimtime="00:06:49.24" />
                    <SPLIT distance="550" swimtime="00:07:30.87" />
                    <SPLIT distance="600" swimtime="00:08:12.51" />
                    <SPLIT distance="650" swimtime="00:08:54.53" />
                    <SPLIT distance="700" swimtime="00:09:36.47" />
                    <SPLIT distance="750" swimtime="00:10:18.63" />
                    <SPLIT distance="800" swimtime="00:11:01.28" />
                    <SPLIT distance="850" swimtime="00:11:43.58" />
                    <SPLIT distance="900" swimtime="00:12:25.46" />
                    <SPLIT distance="950" swimtime="00:13:06.84" />
                    <SPLIT distance="1000" swimtime="00:13:48.53" />
                    <SPLIT distance="1050" swimtime="00:14:30.60" />
                    <SPLIT distance="1100" swimtime="00:15:11.76" />
                    <SPLIT distance="1150" swimtime="00:15:52.82" />
                    <SPLIT distance="1200" swimtime="00:16:33.85" />
                    <SPLIT distance="1250" swimtime="00:17:14.98" />
                    <SPLIT distance="1300" swimtime="00:17:56.48" />
                    <SPLIT distance="1350" swimtime="00:18:38.00" />
                    <SPLIT distance="1400" swimtime="00:19:20.27" />
                    <SPLIT distance="1450" swimtime="00:20:01.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="300" reactiontime="+90" swimtime="00:00:33.76" resultid="2581" heatid="7451" lane="4" entrytime="00:00:34.50" />
                <RESULT eventid="1470" points="305" reactiontime="+72" swimtime="00:01:12.65" resultid="2582" heatid="7669" lane="2" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="304" reactiontime="+73" swimtime="00:02:37.67" resultid="2583" heatid="7770" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:01:58.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-22" firstname="Piotr" gender="M" lastname="Kodur" nation="POL" athleteid="2584">
              <RESULTS>
                <RESULT eventid="1109" points="455" reactiontime="+76" swimtime="00:02:23.06" resultid="2585" heatid="7399" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="100" swimtime="00:01:05.83" />
                    <SPLIT distance="150" swimtime="00:01:48.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="432" reactiontime="+66" swimtime="00:00:29.90" resultid="2586" heatid="7449" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1302" points="487" reactiontime="+75" swimtime="00:01:04.48" resultid="2587" heatid="7549" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="2588" heatid="7637" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1470" points="438" reactiontime="+67" swimtime="00:01:04.41" resultid="2589" heatid="7670" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="336" reactiontime="+88" swimtime="00:01:09.70" resultid="2590" heatid="7747" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="414" reactiontime="+63" swimtime="00:02:22.27" resultid="2591" heatid="7769" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:07.99" />
                    <SPLIT distance="150" swimtime="00:01:44.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-02" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" license="50011520003" athleteid="2592">
              <RESULTS>
                <RESULT eventid="1075" points="383" swimtime="00:00:27.94" resultid="2593" heatid="7368" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="1268" points="411" reactiontime="+78" swimtime="00:01:00.43" resultid="2594" heatid="7519" lane="3" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="378" reactiontime="+88" swimtime="00:02:17.34" resultid="2595" heatid="7702" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:06.48" />
                    <SPLIT distance="150" swimtime="00:01:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="2596" heatid="7748" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="1710" points="384" swimtime="00:04:52.58" resultid="2597" heatid="8055" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:48.36" />
                    <SPLIT distance="200" swimtime="00:02:25.42" />
                    <SPLIT distance="250" swimtime="00:03:04.07" />
                    <SPLIT distance="300" swimtime="00:03:41.76" />
                    <SPLIT distance="350" swimtime="00:04:18.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-23" firstname="Przemysław" gender="M" lastname="Kuca" nation="POL" athleteid="2598">
              <RESULTS>
                <RESULT eventid="1075" points="555" swimtime="00:00:24.70" resultid="2599" heatid="7380" lane="5" entrytime="00:00:24.70" />
                <RESULT eventid="1109" points="584" swimtime="00:02:11.69" resultid="2600" heatid="7407" lane="5" entrytime="00:02:15.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                    <SPLIT distance="100" swimtime="00:01:03.09" />
                    <SPLIT distance="150" swimtime="00:01:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="584" reactiontime="+69" swimtime="00:00:53.76" resultid="2601" heatid="7525" lane="1" entrytime="00:00:52.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="619" reactiontime="+71" swimtime="00:02:08.00" resultid="2602" heatid="7571" lane="3" entrytime="00:02:07.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                    <SPLIT distance="100" swimtime="00:01:00.29" />
                    <SPLIT distance="150" swimtime="00:01:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="603" reactiontime="+70" swimtime="00:01:57.57" resultid="2603" heatid="7706" lane="1" entrytime="00:01:59.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                    <SPLIT distance="100" swimtime="00:00:57.31" />
                    <SPLIT distance="150" swimtime="00:01:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="583" reactiontime="+71" swimtime="00:04:41.75" resultid="2604" heatid="7983" lane="4" entrytime="00:04:53.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                    <SPLIT distance="100" swimtime="00:01:00.80" />
                    <SPLIT distance="150" swimtime="00:01:38.63" />
                    <SPLIT distance="200" swimtime="00:02:15.54" />
                    <SPLIT distance="250" swimtime="00:02:55.49" />
                    <SPLIT distance="300" swimtime="00:03:37.10" />
                    <SPLIT distance="350" swimtime="00:04:09.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="577" reactiontime="+70" swimtime="00:00:58.22" resultid="2605" heatid="7752" lane="2" entrytime="00:00:57.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="598" swimtime="00:04:12.41" resultid="2606" heatid="8058" lane="5" entrytime="00:04:23.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="100" swimtime="00:00:59.14" />
                    <SPLIT distance="150" swimtime="00:01:31.13" />
                    <SPLIT distance="200" swimtime="00:02:03.02" />
                    <SPLIT distance="250" swimtime="00:02:35.24" />
                    <SPLIT distance="300" swimtime="00:03:07.94" />
                    <SPLIT distance="350" swimtime="00:03:40.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" license="50011520004" athleteid="2607">
              <RESULTS>
                <RESULT eventid="1109" points="250" reactiontime="+98" swimtime="00:02:54.56" resultid="2608" heatid="7397" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                    <SPLIT distance="150" swimtime="00:02:13.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="279" swimtime="00:03:04.50" resultid="2609" heatid="7478" lane="5" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                    <SPLIT distance="100" swimtime="00:01:27.98" />
                    <SPLIT distance="150" swimtime="00:02:16.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="256" reactiontime="+97" swimtime="00:01:19.88" resultid="2610" heatid="7545" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="291" reactiontime="+87" swimtime="00:01:23.90" resultid="2611" heatid="7601" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="2612" heatid="7664" lane="5" entrytime="00:01:25.00" />
                <RESULT eventid="1662" points="278" reactiontime="+84" swimtime="00:00:38.65" resultid="2613" heatid="7799" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="485" reactiontime="+70" swimtime="00:01:56.81" resultid="2616" heatid="7934" lane="5" entrytime="00:01:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                    <SPLIT distance="100" swimtime="00:01:03.55" />
                    <SPLIT distance="150" swimtime="00:01:30.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2561" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="2584" number="2" />
                    <RELAYPOSITION athleteid="2555" number="3" />
                    <RELAYPOSITION athleteid="2541" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1377" points="287" reactiontime="+67" swimtime="00:02:19.01" resultid="2615" heatid="7931" lane="2" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:11.84" />
                    <SPLIT distance="150" swimtime="00:01:50.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2579" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="2607" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="2571" number="3" reactiontime="+101" />
                    <RELAYPOSITION athleteid="2592" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1528" points="459" swimtime="00:01:44.68" resultid="2614" heatid="7716" lane="5" entrytime="00:01:45.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.18" />
                    <SPLIT distance="100" swimtime="00:00:52.49" />
                    <SPLIT distance="150" swimtime="00:01:18.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2561" number="1" />
                    <RELAYPOSITION athleteid="2584" number="2" />
                    <RELAYPOSITION athleteid="2555" number="3" />
                    <RELAYPOSITION athleteid="2541" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1528" points="278" reactiontime="+94" swimtime="00:02:03.71" resultid="2617" heatid="7712" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="150" swimtime="00:01:35.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2579" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="2607" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2550" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2592" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AZSSUM" name="AZS Śląski Uniwersytet Medyczny" nation="POL" shortname="AZS Śląski Uniwersytet Medyczn">
          <CONTACT name="Pałka Karol" />
          <ATHLETES>
            <ATHLETE birthdate="1990-03-18" firstname="Karol" gender="M" lastname="Pałka" nation="POL" athleteid="2637">
              <RESULTS>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="2638" heatid="7450" lane="1" entrytime="00:00:35.50" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="2639" heatid="7480" lane="3" entrytime="00:02:58.00" />
                <RESULT eventid="1402" points="239" reactiontime="+78" swimtime="00:01:29.50" resultid="2640" heatid="7604" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="173" reactiontime="+72" swimtime="00:01:27.81" resultid="2641" heatid="7665" lane="1" entrytime="00:01:22.00" />
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="2642" heatid="7767" lane="5" entrytime="00:02:57.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="2643" heatid="7806" lane="5" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CM UJ MAST" name="Collegium Medicum UJ Masters Kraków" nation="POL" region="MAL" shortname="Collegium Medicum UJ Masters K">
          <CONTACT city="Kraków" email="MariuszBaranik@gmail.com" name="Mariusz Baranik" phone="698128222" state="MAŁOP" street="Białoprądnicka 32c/3" zip="31-221" />
          <ATHLETES>
            <ATHLETE birthdate="1969-06-29" firstname="Mariusz" gender="M" lastname="Baranik" nation="POL" athleteid="2645">
              <RESULTS>
                <RESULT eventid="1075" points="425" reactiontime="+79" swimtime="00:00:26.98" resultid="2646" heatid="7373" lane="6" entrytime="00:00:27.30" entrycourse="SCM" />
                <RESULT eventid="1268" points="405" reactiontime="+47" swimtime="00:01:00.74" resultid="2647" heatid="7518" lane="4" entrytime="00:01:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="2648" heatid="7553" lane="2" entrytime="00:01:10.00" entrycourse="SCM" />
                <RESULT eventid="1436" points="428" swimtime="00:00:28.91" resultid="2649" heatid="7641" lane="5" entrytime="00:00:29.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-11" firstname="Marcin" gender="M" lastname="Szczurek" nation="POL" athleteid="2650">
              <RESULTS>
                <RESULT eventid="1302" points="236" swimtime="00:01:22.10" resultid="2651" heatid="7549" lane="5" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="249" swimtime="00:02:37.86" resultid="2652" heatid="7695" lane="5" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:13.52" />
                    <SPLIT distance="150" swimtime="00:01:55.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-08-22" firstname="Mirosław" gender="M" lastname="Woźniak" nation="POL" athleteid="2654">
              <RESULTS>
                <RESULT eventid="1109" points="324" reactiontime="+83" swimtime="00:02:40.18" resultid="2655" heatid="7402" lane="3" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:15.85" />
                    <SPLIT distance="150" swimtime="00:02:03.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="350" reactiontime="+86" swimtime="00:01:03.74" resultid="2656" heatid="7518" lane="6" entrytime="00:01:02.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="342" reactiontime="+90" swimtime="00:01:12.56" resultid="2657" heatid="7551" lane="6" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="303" swimtime="00:02:27.82" resultid="2658" heatid="7697" lane="5" entrytime="00:02:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:50.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="UJ CM Kraków" nation="POL" region="MAL">
          <CONTACT city="Kraków" email="drab.magdalena@wp.pl" name="Drab" phone="604957110" state="MAL" street="Obozowa 76/10" zip="30-383" />
          <ATHLETES>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="2660">
              <RESULTS>
                <RESULT eventid="1058" points="554" reactiontime="+84" swimtime="00:00:28.30" resultid="2661" heatid="7344" lane="1" entrytime="00:00:28.31" />
                <RESULT eventid="1092" points="587" reactiontime="+84" swimtime="00:02:28.76" resultid="2662" heatid="7389" lane="3" entrytime="00:02:29.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="434" reactiontime="+87" swimtime="00:02:57.67" resultid="2663" heatid="7469" lane="4" entrytime="00:02:48.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:22.99" />
                    <SPLIT distance="150" swimtime="00:02:10.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="593" reactiontime="+87" swimtime="00:01:08.69" resultid="2664" heatid="7537" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="547" reactiontime="+82" swimtime="00:01:16.65" resultid="2665" heatid="7591" lane="3" entrytime="00:01:15.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="583" reactiontime="+85" swimtime="00:02:13.04" resultid="2666" heatid="7685" lane="3" entrytime="00:02:12.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:01:03.68" />
                    <SPLIT distance="150" swimtime="00:01:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="531" reactiontime="+84" swimtime="00:00:35.56" resultid="2667" heatid="7787" lane="3" entrytime="00:00:34.36" />
                <RESULT eventid="1693" points="530" reactiontime="+86" swimtime="00:04:50.27" resultid="2668" heatid="8025" lane="3" entrytime="00:04:48.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:45.45" />
                    <SPLIT distance="200" swimtime="00:02:22.83" />
                    <SPLIT distance="250" swimtime="00:03:00.03" />
                    <SPLIT distance="300" swimtime="00:03:37.15" />
                    <SPLIT distance="350" swimtime="00:04:14.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" name="KS niezrzeszeni.pl" nation="POL" region="WA">
          <CONTACT email="niezrzeszeni.pl@gmail.com" internet="niezrzeszeni.pl" name="wawer maylda katarzyna" />
          <ATHLETES>
            <ATHLETE birthdate="1973-08-26" firstname="Małgorzata" gender="F" lastname="Piechura" nation="POL" athleteid="2670">
              <RESULTS>
                <RESULT eventid="1092" points="116" reactiontime="+123" swimtime="00:04:15.01" resultid="2671" heatid="7384" lane="1" entrytime="00:04:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.31" />
                    <SPLIT distance="150" swimtime="00:03:16.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="129" reactiontime="+114" swimtime="00:01:40.93" resultid="2672" heatid="7488" lane="4" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="124" reactiontime="+113" swimtime="00:01:55.58" resultid="2673" heatid="7527" lane="3" entrytime="00:01:54.00" />
                <RESULT eventid="1487" points="116" reactiontime="+121" swimtime="00:03:47.72" resultid="2674" heatid="7676" lane="2" entrytime="00:03:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:52.94" />
                    <SPLIT distance="150" swimtime="00:02:54.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="130" reactiontime="+122" swimtime="00:07:42.79" resultid="2675" heatid="8019" lane="4" entrytime="00:07:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.42" />
                    <SPLIT distance="100" swimtime="00:01:47.16" />
                    <SPLIT distance="150" swimtime="00:02:46.54" />
                    <SPLIT distance="200" swimtime="00:03:48.63" />
                    <SPLIT distance="250" swimtime="00:04:47.87" />
                    <SPLIT distance="300" swimtime="00:05:48.36" />
                    <SPLIT distance="350" swimtime="00:06:50.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="2676">
              <RESULTS>
                <RESULT eventid="1165" points="158" reactiontime="+134" swimtime="00:26:10.47" resultid="2677" heatid="7909" lane="4" entrytime="00:26:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                    <SPLIT distance="100" swimtime="00:01:37.33" />
                    <SPLIT distance="150" swimtime="00:02:29.11" />
                    <SPLIT distance="200" swimtime="00:03:20.55" />
                    <SPLIT distance="250" swimtime="00:04:12.14" />
                    <SPLIT distance="300" swimtime="00:05:04.09" />
                    <SPLIT distance="350" swimtime="00:05:55.78" />
                    <SPLIT distance="400" swimtime="00:06:47.77" />
                    <SPLIT distance="450" swimtime="00:07:40.30" />
                    <SPLIT distance="500" swimtime="00:08:32.97" />
                    <SPLIT distance="550" swimtime="00:09:25.63" />
                    <SPLIT distance="600" swimtime="00:10:18.50" />
                    <SPLIT distance="650" swimtime="00:11:10.84" />
                    <SPLIT distance="700" swimtime="00:12:03.85" />
                    <SPLIT distance="750" swimtime="00:12:57.23" />
                    <SPLIT distance="800" swimtime="00:13:49.91" />
                    <SPLIT distance="850" swimtime="00:14:43.36" />
                    <SPLIT distance="900" swimtime="00:15:35.94" />
                    <SPLIT distance="950" swimtime="00:16:28.65" />
                    <SPLIT distance="1000" swimtime="00:17:21.94" />
                    <SPLIT distance="1050" swimtime="00:18:14.58" />
                    <SPLIT distance="1100" swimtime="00:19:07.74" />
                    <SPLIT distance="1150" swimtime="00:20:00.90" />
                    <SPLIT distance="1200" swimtime="00:20:54.52" />
                    <SPLIT distance="1250" swimtime="00:21:48.38" />
                    <SPLIT distance="1300" swimtime="00:22:42.07" />
                    <SPLIT distance="1350" swimtime="00:23:34.90" />
                    <SPLIT distance="1400" swimtime="00:24:28.96" />
                    <SPLIT distance="1450" swimtime="00:25:23.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="78" reactiontime="+136" swimtime="00:04:14.79" resultid="2678" heatid="7565" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.40" />
                    <SPLIT distance="100" swimtime="00:02:04.30" />
                    <SPLIT distance="150" swimtime="00:03:11.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="112" swimtime="00:08:07.82" resultid="2679" heatid="7974" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.23" />
                    <SPLIT distance="100" swimtime="00:01:57.07" />
                    <SPLIT distance="150" swimtime="00:03:09.47" />
                    <SPLIT distance="200" swimtime="00:04:21.19" />
                    <SPLIT distance="250" swimtime="00:05:25.38" />
                    <SPLIT distance="300" swimtime="00:06:27.20" />
                    <SPLIT distance="350" swimtime="00:07:19.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="154" reactiontime="+131" swimtime="00:06:36.16" resultid="2680" heatid="8046" lane="4" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.84" />
                    <SPLIT distance="100" swimtime="00:01:32.89" />
                    <SPLIT distance="150" swimtime="00:02:23.46" />
                    <SPLIT distance="200" swimtime="00:03:14.80" />
                    <SPLIT distance="250" swimtime="00:04:05.62" />
                    <SPLIT distance="300" swimtime="00:04:57.44" />
                    <SPLIT distance="350" swimtime="00:05:48.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="2681">
              <RESULTS>
                <RESULT eventid="1109" points="146" reactiontime="+114" swimtime="00:03:28.87" resultid="2682" heatid="7394" lane="2" entrytime="00:03:35.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.96" />
                    <SPLIT distance="100" swimtime="00:01:37.53" />
                    <SPLIT distance="150" swimtime="00:02:39.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="174" reactiontime="+130" swimtime="00:25:21.68" resultid="2683" heatid="7910" lane="1" entrytime="00:26:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:01:34.41" />
                    <SPLIT distance="150" swimtime="00:02:25.12" />
                    <SPLIT distance="200" swimtime="00:03:16.29" />
                    <SPLIT distance="250" swimtime="00:04:08.18" />
                    <SPLIT distance="300" swimtime="00:04:59.46" />
                    <SPLIT distance="350" swimtime="00:05:50.54" />
                    <SPLIT distance="400" swimtime="00:06:42.98" />
                    <SPLIT distance="450" swimtime="00:07:35.37" />
                    <SPLIT distance="500" swimtime="00:08:27.07" />
                    <SPLIT distance="550" swimtime="00:09:18.98" />
                    <SPLIT distance="600" swimtime="00:10:10.90" />
                    <SPLIT distance="650" swimtime="00:11:02.53" />
                    <SPLIT distance="700" swimtime="00:11:53.63" />
                    <SPLIT distance="750" swimtime="00:12:44.85" />
                    <SPLIT distance="800" swimtime="00:13:35.80" />
                    <SPLIT distance="850" swimtime="00:14:27.41" />
                    <SPLIT distance="900" swimtime="00:15:18.63" />
                    <SPLIT distance="950" swimtime="00:16:09.87" />
                    <SPLIT distance="1000" swimtime="00:17:53.00" />
                    <SPLIT distance="1050" swimtime="00:18:45.13" />
                    <SPLIT distance="1100" swimtime="00:19:35.49" />
                    <SPLIT distance="1150" swimtime="00:20:26.86" />
                    <SPLIT distance="1200" swimtime="00:21:17.43" />
                    <SPLIT distance="1250" swimtime="00:22:08.11" />
                    <SPLIT distance="1300" swimtime="00:22:58.80" />
                    <SPLIT distance="1350" swimtime="00:23:48.03" />
                    <SPLIT distance="1400" swimtime="00:24:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="177" reactiontime="+70" swimtime="00:00:40.20" resultid="2684" heatid="7446" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1470" points="164" reactiontime="+71" swimtime="00:01:29.26" resultid="2685" heatid="7663" lane="2" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="2686" heatid="7976" lane="3" entrytime="00:07:39.79" />
                <RESULT eventid="1628" points="171" reactiontime="+74" swimtime="00:03:11.11" resultid="2687" heatid="7765" lane="3" entrytime="00:03:16.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                    <SPLIT distance="100" swimtime="00:01:31.44" />
                    <SPLIT distance="150" swimtime="00:02:21.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-04-08" firstname="Wojciech" gender="M" lastname="Staruch" nation="POL" athleteid="2688">
              <RESULTS>
                <RESULT eventid="1109" points="137" reactiontime="+86" swimtime="00:03:33.30" resultid="2689" heatid="7394" lane="4" entrytime="00:03:33.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:40.49" />
                    <SPLIT distance="150" swimtime="00:02:39.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="178" reactiontime="+82" swimtime="00:03:34.48" resultid="2690" heatid="7474" lane="2" entrytime="00:03:39.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                    <SPLIT distance="100" swimtime="00:01:43.85" />
                    <SPLIT distance="150" swimtime="00:02:40.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="178" reactiontime="+83" swimtime="00:01:30.22" resultid="2691" heatid="7542" lane="3" entrytime="00:01:30.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="198" reactiontime="+81" swimtime="00:01:35.37" resultid="2692" heatid="7597" lane="6" entrytime="00:01:38.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="176" reactiontime="+82" swimtime="00:00:38.87" resultid="2693" heatid="7625" lane="1" entrytime="00:00:46.61" />
                <RESULT eventid="1594" points="144" reactiontime="+89" swimtime="00:01:32.49" resultid="2694" heatid="7740" lane="6" entrytime="00:01:43.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="216" reactiontime="+77" swimtime="00:00:42.05" resultid="2695" heatid="7795" lane="2" entrytime="00:00:42.38" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMT SZCZEC" name="Swimming Masters Team Szczecin" nation="POL" region="ZAC">
          <CONTACT city="Szczecin" email="teczowy.dyndol@gmail.com" name="Brodacki Maciej" />
          <ATHLETES>
            <ATHLETE birthdate="1993-01-20" firstname="Agnieszka" gender="F" lastname="Krzyżostaniak" nation="POL" athleteid="2697">
              <RESULTS>
                <RESULT eventid="1148" points="546" reactiontime="+80" swimtime="00:09:52.48" resultid="2698" heatid="7906" lane="3" entrytime="00:10:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:07.86" />
                    <SPLIT distance="150" swimtime="00:01:43.24" />
                    <SPLIT distance="200" swimtime="00:02:20.20" />
                    <SPLIT distance="250" swimtime="00:02:57.60" />
                    <SPLIT distance="300" swimtime="00:03:35.41" />
                    <SPLIT distance="350" swimtime="00:04:13.15" />
                    <SPLIT distance="400" swimtime="00:04:51.39" />
                    <SPLIT distance="450" swimtime="00:05:29.70" />
                    <SPLIT distance="500" swimtime="00:06:08.00" />
                    <SPLIT distance="550" swimtime="00:06:46.20" />
                    <SPLIT distance="600" swimtime="00:07:23.97" />
                    <SPLIT distance="650" swimtime="00:08:01.19" />
                    <SPLIT distance="700" swimtime="00:08:38.75" />
                    <SPLIT distance="750" swimtime="00:09:16.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="562" reactiontime="+67" swimtime="00:00:31.14" resultid="2699" heatid="7441" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1251" points="549" reactiontime="+81" swimtime="00:01:02.26" resultid="2700" heatid="7497" lane="4" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="532" reactiontime="+77" swimtime="00:01:08.16" resultid="2701" heatid="7658" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="507" reactiontime="+84" swimtime="00:02:19.36" resultid="2702" heatid="7684" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="150" swimtime="00:01:44.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" status="DNS" swimtime="00:00:00.00" resultid="2703" heatid="8025" lane="4" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-09" firstname="Helena" gender="F" lastname="Szulc" nation="POL" athleteid="2704">
              <RESULTS>
                <RESULT eventid="1092" points="312" reactiontime="+95" swimtime="00:03:03.59" resultid="2705" heatid="7386" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:25.13" />
                    <SPLIT distance="150" swimtime="00:02:18.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="323" reactiontime="+88" swimtime="00:01:24.10" resultid="2706" heatid="7532" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="258" reactiontime="+87" swimtime="00:00:38.26" resultid="2707" heatid="7616" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1645" points="270" reactiontime="+91" swimtime="00:00:44.54" resultid="2708" heatid="7781" lane="4" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-15" firstname="Paulina" gender="F" lastname="Kotfica" nation="POL" athleteid="2709">
              <RESULTS>
                <RESULT eventid="1183" status="DNS" swimtime="00:00:00.00" resultid="2711" heatid="7441" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="2712" heatid="7497" lane="5" entrytime="00:01:05.00" />
                <RESULT eventid="1487" status="DNS" swimtime="00:00:00.00" resultid="2713" heatid="7684" lane="5" entrytime="00:02:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-12" firstname="Kamila" gender="F" lastname="Gębka" nation="POL" athleteid="2714">
              <RESULTS>
                <RESULT eventid="1092" points="343" swimtime="00:02:57.86" resultid="2715" heatid="7387" lane="5" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:01:23.96" />
                    <SPLIT distance="150" swimtime="00:02:14.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="324" reactiontime="+90" swimtime="00:03:15.73" resultid="2716" heatid="7468" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                    <SPLIT distance="100" swimtime="00:01:34.49" />
                    <SPLIT distance="150" swimtime="00:02:25.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="360" reactiontime="+87" swimtime="00:01:21.14" resultid="2717" heatid="7532" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="318" reactiontime="+88" swimtime="00:01:31.82" resultid="2718" heatid="7589" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="279" swimtime="00:00:37.27" resultid="2719" heatid="7617" lane="5" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="Brodacki" nation="POL" athleteid="2721">
              <RESULTS>
                <RESULT eventid="1075" points="498" reactiontime="+79" swimtime="00:00:25.60" resultid="2722" heatid="7378" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1109" points="473" reactiontime="+82" swimtime="00:02:21.25" resultid="2723" heatid="7404" lane="3" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="100" swimtime="00:01:05.77" />
                    <SPLIT distance="150" swimtime="00:01:48.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="534" reactiontime="+80" swimtime="00:00:55.37" resultid="2724" heatid="7523" lane="1" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="503" reactiontime="+80" swimtime="00:01:03.79" resultid="2725" heatid="7555" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="483" reactiontime="+82" swimtime="00:02:06.61" resultid="2726" heatid="7702" lane="3" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                    <SPLIT distance="100" swimtime="00:01:00.05" />
                    <SPLIT distance="150" swimtime="00:01:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="380" swimtime="00:00:34.85" resultid="2728" heatid="7788" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="2729" heatid="8054" lane="4" entrytime="00:05:00.00" />
                <RESULT eventid="1559" points="414" reactiontime="+85" swimtime="00:05:15.77" resultid="8003" heatid="7980" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:52.72" />
                    <SPLIT distance="200" swimtime="00:02:32.99" />
                    <SPLIT distance="250" swimtime="00:03:19.17" />
                    <SPLIT distance="300" swimtime="00:04:06.25" />
                    <SPLIT distance="350" swimtime="00:04:42.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-13" firstname="Piotr" gender="M" lastname="Kozłowski" nation="POL" athleteid="2730">
              <RESULTS>
                <RESULT eventid="1165" points="285" swimtime="00:21:31.39" resultid="2731" heatid="7915" lane="5" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:00.64" />
                    <SPLIT distance="200" swimtime="00:02:43.11" />
                    <SPLIT distance="250" swimtime="00:03:25.79" />
                    <SPLIT distance="300" swimtime="00:04:08.78" />
                    <SPLIT distance="350" swimtime="00:04:51.10" />
                    <SPLIT distance="400" swimtime="00:05:33.52" />
                    <SPLIT distance="450" swimtime="00:06:16.38" />
                    <SPLIT distance="500" swimtime="00:06:59.32" />
                    <SPLIT distance="550" swimtime="00:07:42.00" />
                    <SPLIT distance="600" swimtime="00:08:25.01" />
                    <SPLIT distance="650" swimtime="00:09:08.35" />
                    <SPLIT distance="700" swimtime="00:09:51.58" />
                    <SPLIT distance="750" swimtime="00:10:34.58" />
                    <SPLIT distance="800" swimtime="00:11:17.88" />
                    <SPLIT distance="850" swimtime="00:12:01.33" />
                    <SPLIT distance="900" swimtime="00:12:44.88" />
                    <SPLIT distance="950" swimtime="00:13:28.64" />
                    <SPLIT distance="1000" swimtime="00:14:12.39" />
                    <SPLIT distance="1050" swimtime="00:14:56.36" />
                    <SPLIT distance="1100" swimtime="00:15:40.46" />
                    <SPLIT distance="1150" swimtime="00:16:24.52" />
                    <SPLIT distance="1200" swimtime="00:17:08.56" />
                    <SPLIT distance="1250" swimtime="00:17:52.80" />
                    <SPLIT distance="1300" swimtime="00:18:36.65" />
                    <SPLIT distance="1350" swimtime="00:19:20.75" />
                    <SPLIT distance="1400" swimtime="00:20:04.31" />
                    <SPLIT distance="1450" swimtime="00:20:48.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="330" reactiontime="+93" swimtime="00:01:05.03" resultid="2732" heatid="7515" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="295" reactiontime="+93" swimtime="00:02:29.14" resultid="2733" heatid="7698" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                    <SPLIT distance="150" swimtime="00:01:52.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="2734" heatid="8053" lane="1" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-27" firstname="Rafał" gender="M" lastname="Lisiecki" nation="POL" athleteid="2735">
              <RESULTS>
                <RESULT eventid="1075" points="404" reactiontime="+88" swimtime="00:00:27.46" resultid="2736" heatid="7372" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1200" points="394" reactiontime="+71" swimtime="00:00:30.82" resultid="2737" heatid="7457" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1268" points="410" reactiontime="+84" swimtime="00:01:00.46" resultid="2738" heatid="7519" lane="4" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="387" reactiontime="+72" swimtime="00:01:07.13" resultid="2739" heatid="7672" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-20" firstname="Marcin" gender="M" lastname="Łogin" nation="POL" athleteid="2740">
              <RESULTS>
                <RESULT eventid="1075" points="322" reactiontime="+91" swimtime="00:00:29.61" resultid="2741" heatid="7362" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1234" points="290" reactiontime="+97" swimtime="00:03:02.13" resultid="2742" heatid="7479" lane="2" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:01:27.21" />
                    <SPLIT distance="150" swimtime="00:02:16.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="349" reactiontime="+94" swimtime="00:01:18.95" resultid="2743" heatid="7604" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="283" reactiontime="+93" swimtime="00:00:33.17" resultid="2744" heatid="7632" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="2745" heatid="7805" lane="5" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="Roenig" nation="POL" athleteid="2746">
              <RESULTS>
                <RESULT eventid="1075" points="358" swimtime="00:00:28.57" resultid="2747" heatid="7363" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1234" points="343" reactiontime="+94" swimtime="00:02:52.32" resultid="2748" heatid="7479" lane="4" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:08.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="390" reactiontime="+95" swimtime="00:01:16.06" resultid="2749" heatid="7607" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="2750" heatid="7810" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-28" firstname="Hubert" gender="M" lastname="Frączyk" nation="POL" athleteid="2751">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="2752" heatid="7359" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1402" points="165" reactiontime="+89" swimtime="00:01:41.30" resultid="2753" heatid="7596" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="198" reactiontime="+90" swimtime="00:00:43.27" resultid="2754" heatid="7794" lane="3" entrytime="00:00:43.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-05" firstname="Rafał" gender="M" lastname="Dobrowolski" nation="POL" athleteid="2755">
              <RESULTS>
                <RESULT eventid="1075" points="237" reactiontime="+78" swimtime="00:00:32.77" resultid="2756" heatid="7358" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1268" points="196" reactiontime="+78" swimtime="00:01:17.25" resultid="2757" heatid="7505" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="212" swimtime="00:01:33.23" resultid="2758" heatid="7597" lane="5" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="231" reactiontime="+76" swimtime="00:00:41.14" resultid="2759" heatid="7795" lane="3" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-21" firstname="Michał" gender="M" lastname="Krysiak" nation="POL" athleteid="2760">
              <RESULTS>
                <RESULT eventid="1075" points="425" reactiontime="+83" swimtime="00:00:27.00" resultid="2761" heatid="7376" lane="6" entrytime="00:00:26.50" />
                <RESULT eventid="1109" points="318" reactiontime="+84" swimtime="00:02:41.21" resultid="2762" heatid="7404" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:13.39" />
                    <SPLIT distance="150" swimtime="00:02:02.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="393" reactiontime="+79" swimtime="00:01:01.35" resultid="2763" heatid="7522" lane="1" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="358" swimtime="00:02:33.56" resultid="2764" heatid="7570" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="150" swimtime="00:01:54.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="418" reactiontime="+78" swimtime="00:00:29.15" resultid="2765" heatid="7642" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="2766" heatid="7979" lane="1" entrytime="00:06:10.00" />
                <RESULT eventid="1594" points="412" swimtime="00:01:05.10" resultid="2767" heatid="7750" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="345" reactiontime="+72" swimtime="00:02:10.86" resultid="2775" heatid="7928" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:06.93" />
                    <SPLIT distance="150" swimtime="00:01:36.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2735" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2740" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="2760" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2751" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="314" reactiontime="+86" swimtime="00:01:58.79" resultid="2776" heatid="7709" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="100" swimtime="00:01:01.68" />
                    <SPLIT distance="150" swimtime="00:01:31.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2735" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="2740" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2760" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="2751" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1377" points="365" reactiontime="+75" swimtime="00:02:08.38" resultid="2777" heatid="7928" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="150" swimtime="00:01:36.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2721" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="2746" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="2730" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="2755" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="343" reactiontime="+88" swimtime="00:01:55.35" resultid="2778" heatid="7709" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                    <SPLIT distance="100" swimtime="00:00:59.74" />
                    <SPLIT distance="150" swimtime="00:01:29.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2721" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="2746" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2730" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="2755" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1370" status="DNS" swimtime="00:00:00.00" resultid="2773" heatid="7572" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2697" number="1" />
                    <RELAYPOSITION athleteid="2714" number="2" />
                    <RELAYPOSITION athleteid="2704" number="3" />
                    <RELAYPOSITION athleteid="2709" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1521" status="DNS" swimtime="00:00:00.00" resultid="2774" heatid="7707" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2697" number="1" />
                    <RELAYPOSITION athleteid="2714" number="2" />
                    <RELAYPOSITION athleteid="2704" number="3" />
                    <RELAYPOSITION athleteid="2709" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1679" points="344" reactiontime="+69" swimtime="00:02:10.89" resultid="2770" heatid="7815" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="150" swimtime="00:01:45.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2697" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2704" number="2" />
                    <RELAYPOSITION athleteid="2760" number="3" />
                    <RELAYPOSITION athleteid="2721" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1126" points="333" reactiontime="+83" swimtime="00:01:56.43" resultid="2771" heatid="7411" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                    <SPLIT distance="100" swimtime="00:00:55.47" />
                    <SPLIT distance="150" swimtime="00:01:29.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2697" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2704" number="2" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2735" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="2760" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="2772" heatid="7814" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2709" number="1" />
                    <RELAYPOSITION athleteid="2704" number="2" />
                    <RELAYPOSITION athleteid="2721" number="3" />
                    <RELAYPOSITION athleteid="2760" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="WOPR Tczew" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1987-01-01" firstname="Aleksandra" gender="F" lastname="Hebel " nation="POL" athleteid="2780">
              <RESULTS>
                <RESULT eventid="1058" points="356" reactiontime="+96" swimtime="00:00:32.78" resultid="2781" heatid="7340" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1183" points="231" reactiontime="+96" swimtime="00:00:41.86" resultid="2782" heatid="7435" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1251" points="293" swimtime="00:01:16.74" resultid="2783" heatid="7494" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="211" reactiontime="+112" swimtime="00:01:32.71" resultid="2784" heatid="7652" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="271" reactiontime="+105" swimtime="00:02:51.61" resultid="2785" heatid="7680" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:21.17" />
                    <SPLIT distance="150" swimtime="00:02:06.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="250" reactiontime="+95" swimtime="00:03:10.45" resultid="2786" heatid="7756" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:33.01" />
                    <SPLIT distance="150" swimtime="00:02:22.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Andrzej " gender="M" lastname="Gołembiewski" nation="POL" athleteid="2787">
              <RESULTS>
                <RESULT eventid="1075" points="411" reactiontime="+88" swimtime="00:00:27.29" resultid="2788" heatid="7371" lane="2" entrytime="00:00:27.80" />
                <RESULT eventid="1234" points="389" reactiontime="+94" swimtime="00:02:45.21" resultid="2789" heatid="7482" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:16.87" />
                    <SPLIT distance="150" swimtime="00:02:00.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="412" swimtime="00:01:00.35" resultid="2790" heatid="7517" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="459" reactiontime="+89" swimtime="00:01:12.04" resultid="2791" heatid="7608" lane="6" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="401" reactiontime="+89" swimtime="00:02:14.65" resultid="2792" heatid="7700" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:04.27" />
                    <SPLIT distance="150" swimtime="00:01:40.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="436" reactiontime="+91" swimtime="00:00:33.28" resultid="2793" heatid="7807" lane="3" entrytime="00:00:34.80" />
                <RESULT eventid="1710" points="362" reactiontime="+95" swimtime="00:04:58.32" resultid="2794" heatid="8054" lane="6" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                    <SPLIT distance="150" swimtime="00:01:45.76" />
                    <SPLIT distance="200" swimtime="00:02:23.87" />
                    <SPLIT distance="250" swimtime="00:03:02.99" />
                    <SPLIT distance="300" swimtime="00:03:42.24" />
                    <SPLIT distance="350" swimtime="00:04:21.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Marek" gender="M" lastname="Stuczyński " nation="POL" athleteid="2795">
              <RESULTS>
                <RESULT eventid="1075" points="531" reactiontime="+79" swimtime="00:00:25.06" resultid="2796" heatid="7380" lane="6" entrytime="00:00:25.00" />
                <RESULT eventid="1302" points="492" reactiontime="+80" swimtime="00:01:04.28" resultid="2797" heatid="7559" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="526" reactiontime="+81" swimtime="00:01:08.88" resultid="2798" heatid="7610" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="572" reactiontime="+78" swimtime="00:00:30.41" resultid="2799" heatid="7812" lane="2" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Plavecky klub Zabreh" nation="CZE">
          <ATHLETES>
            <ATHLETE birthdate="1973-01-01" firstname="Petr" gender="M" lastname="HORVAT " nation="POL" athleteid="2806">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="2807" heatid="7365" lane="2" entrytime="00:00:29.62" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2808" heatid="7399" lane="3" entrytime="00:02:46.44" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="2809" heatid="7480" lane="2" entrytime="00:02:59.64" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="2810" heatid="7603" lane="3" entrytime="00:01:24.69" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="2811" heatid="7701" lane="5" entrytime="00:02:34.31" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Masters Bialystok" nation="POL">
          <CONTACT email="mbzgloszenia@gmail.com" name="MICHALIK DOMINIKA" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="2813">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1148" points="482" reactiontime="+90" swimtime="00:10:17.70" resultid="2814" heatid="7906" lane="1" entrytime="00:10:30.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:11.65" />
                    <SPLIT distance="150" swimtime="00:01:49.60" />
                    <SPLIT distance="200" swimtime="00:02:28.18" />
                    <SPLIT distance="250" swimtime="00:03:07.24" />
                    <SPLIT distance="300" swimtime="00:03:46.46" />
                    <SPLIT distance="350" swimtime="00:04:25.89" />
                    <SPLIT distance="400" swimtime="00:05:05.22" />
                    <SPLIT distance="450" swimtime="00:05:45.03" />
                    <SPLIT distance="500" swimtime="00:06:24.55" />
                    <SPLIT distance="550" swimtime="00:07:03.80" />
                    <SPLIT distance="600" swimtime="00:07:42.97" />
                    <SPLIT distance="650" swimtime="00:08:22.40" />
                    <SPLIT distance="700" swimtime="00:09:01.88" />
                    <SPLIT distance="750" swimtime="00:09:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="477" reactiontime="+85" swimtime="00:01:05.27" resultid="2815" heatid="7496" lane="2" entrytime="00:01:07.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1487" points="505" reactiontime="+85" swimtime="00:02:19.55" resultid="2816" heatid="7684" lane="1" entrytime="00:02:25.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:08.61" />
                    <SPLIT distance="150" swimtime="00:01:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1693" points="492" reactiontime="+89" swimtime="00:04:57.46" resultid="2817" heatid="8025" lane="2" entrytime="00:05:03.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="150" swimtime="00:01:48.88" />
                    <SPLIT distance="200" swimtime="00:02:27.08" />
                    <SPLIT distance="250" swimtime="00:03:05.42" />
                    <SPLIT distance="300" swimtime="00:03:43.91" />
                    <SPLIT distance="350" swimtime="00:04:21.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Bartosz" gender="M" lastname="Bogdanowicz" nation="POL" athleteid="2818">
              <RESULTS>
                <RESULT eventid="1336" points="283" reactiontime="+80" swimtime="00:02:46.12" resultid="2819" heatid="7569" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:21.12" />
                    <SPLIT distance="150" swimtime="00:02:05.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="315" reactiontime="+72" swimtime="00:02:35.92" resultid="2821" heatid="7772" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="150" swimtime="00:01:57.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Magdalena" gender="F" lastname="Tomaszuk" nation="POL" athleteid="2822">
              <RESULTS>
                <RESULT eventid="1183" points="220" reactiontime="+114" swimtime="00:00:42.52" resultid="2823" heatid="7435" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1251" points="334" reactiontime="+106" swimtime="00:01:13.52" resultid="2824" heatid="7493" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" status="DNS" swimtime="00:00:00.00" resultid="2825" heatid="7615" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="2826" heatid="7651" lane="4" entrytime="00:01:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Elżbieta" gender="F" lastname="Piwowarczyk" nation="POL" athleteid="2827">
              <RESULTS>
                <RESULT eventid="1058" points="326" reactiontime="+81" swimtime="00:00:33.77" resultid="2828" heatid="7340" lane="6" entrytime="00:00:33.80" />
                <RESULT eventid="1092" points="294" reactiontime="+83" swimtime="00:03:07.31" resultid="2829" heatid="7386" lane="1" entrytime="00:03:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="100" swimtime="00:01:29.57" />
                    <SPLIT distance="150" swimtime="00:02:25.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="253" reactiontime="+73" swimtime="00:00:40.61" resultid="2830" heatid="7436" lane="2" entrytime="00:00:40.10" />
                <RESULT eventid="1251" points="307" reactiontime="+77" swimtime="00:01:15.57" resultid="2831" heatid="7494" lane="3" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="256" reactiontime="+71" swimtime="00:01:26.98" resultid="2832" heatid="7652" lane="3" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="289" reactiontime="+85" swimtime="00:02:48.01" resultid="2833" heatid="7681" lane="2" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:01:20.40" />
                    <SPLIT distance="150" swimtime="00:02:04.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="251" reactiontime="+75" swimtime="00:03:10.14" resultid="2834" heatid="7758" lane="6" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                    <SPLIT distance="100" swimtime="00:01:31.79" />
                    <SPLIT distance="150" swimtime="00:02:21.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="267" reactiontime="+87" swimtime="00:06:04.50" resultid="2835" heatid="8022" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:24.16" />
                    <SPLIT distance="150" swimtime="00:02:10.26" />
                    <SPLIT distance="200" swimtime="00:02:57.07" />
                    <SPLIT distance="250" swimtime="00:03:43.84" />
                    <SPLIT distance="300" swimtime="00:04:30.89" />
                    <SPLIT distance="350" swimtime="00:05:18.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Joanna" gender="F" lastname="Wasilewicz" nation="POL" athleteid="2836">
              <RESULTS>
                <RESULT eventid="1058" points="252" swimtime="00:00:36.78" resultid="2837" heatid="7337" lane="5" entrytime="00:00:36.90" />
                <RESULT eventid="1251" points="199" reactiontime="+58" swimtime="00:01:27.24" resultid="2838" heatid="7490" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" status="DNS" swimtime="00:00:00.00" resultid="2839" heatid="7528" lane="5" entrytime="00:01:40.00" />
                <RESULT eventid="1487" points="174" reactiontime="+92" swimtime="00:03:19.06" resultid="2840" heatid="7678" lane="6" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                    <SPLIT distance="100" swimtime="00:01:33.59" />
                    <SPLIT distance="150" swimtime="00:02:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="2841" heatid="7778" lane="6" entrytime="00:00:55.00" />
                <RESULT eventid="1693" status="DNS" swimtime="00:00:00.00" resultid="2842" heatid="8020" lane="3" entrytime="00:06:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosław" gender="M" lastname="Matusik" nation="POL" athleteid="2843">
              <RESULTS>
                <RESULT eventid="1075" points="234" swimtime="00:00:32.90" resultid="2844" heatid="7357" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1165" status="DNF" swimtime="00:00:00.00" resultid="2845" heatid="7911" lane="5" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                    <SPLIT distance="100" swimtime="00:01:27.16" />
                    <SPLIT distance="150" swimtime="00:02:14.31" />
                    <SPLIT distance="200" swimtime="00:03:01.50" />
                    <SPLIT distance="250" swimtime="00:03:49.85" />
                    <SPLIT distance="300" swimtime="00:04:37.67" />
                    <SPLIT distance="350" swimtime="00:05:25.75" />
                    <SPLIT distance="400" swimtime="00:06:15.01" />
                    <SPLIT distance="450" swimtime="00:07:03.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="2846" heatid="7507" lane="4" entrytime="00:01:14.00" />
                <RESULT eventid="1436" points="248" reactiontime="+97" swimtime="00:00:34.68" resultid="2847" heatid="7633" lane="1" entrytime="00:00:33.50" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="2848" heatid="7694" lane="3" entrytime="00:02:40.00" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="2849" heatid="7742" lane="5" entrytime="00:01:24.00" />
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="2850" heatid="8050" lane="1" entrytime="00:05:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="UKS Trójka Oborniki" nation="POL" region="WIE">
          <CONTACT city="Oborniki" email="janwol@poczta,onet.pl" name="Wolniewicz Janusz" phone="791064667" state="WIE" street="Piłsudskiego 49/42" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="2852">
              <RESULTS>
                <RESULT eventid="1075" points="180" swimtime="00:00:35.92" resultid="2853" heatid="7352" lane="5" entrytime="00:00:35.11" entrycourse="SCM" />
                <RESULT eventid="1165" points="111" reactiontime="+104" swimtime="00:29:25.48" resultid="2854" heatid="7909" lane="6" entrytime="00:28:22.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.11" />
                    <SPLIT distance="100" swimtime="00:01:46.24" />
                    <SPLIT distance="150" swimtime="00:02:43.04" />
                    <SPLIT distance="200" swimtime="00:03:41.07" />
                    <SPLIT distance="250" swimtime="00:04:39.48" />
                    <SPLIT distance="300" swimtime="00:05:37.01" />
                    <SPLIT distance="350" swimtime="00:06:34.56" />
                    <SPLIT distance="400" swimtime="00:07:32.58" />
                    <SPLIT distance="450" swimtime="00:08:31.10" />
                    <SPLIT distance="500" swimtime="00:09:30.23" />
                    <SPLIT distance="550" swimtime="00:10:29.06" />
                    <SPLIT distance="600" swimtime="00:11:28.51" />
                    <SPLIT distance="650" swimtime="00:12:27.27" />
                    <SPLIT distance="700" swimtime="00:13:26.41" />
                    <SPLIT distance="750" swimtime="00:14:25.43" />
                    <SPLIT distance="800" swimtime="00:15:24.48" />
                    <SPLIT distance="850" swimtime="00:16:24.36" />
                    <SPLIT distance="900" swimtime="00:17:24.17" />
                    <SPLIT distance="950" swimtime="00:18:22.81" />
                    <SPLIT distance="1000" swimtime="00:19:22.86" />
                    <SPLIT distance="1050" swimtime="00:20:23.02" />
                    <SPLIT distance="1100" swimtime="00:21:24.18" />
                    <SPLIT distance="1150" swimtime="00:22:24.61" />
                    <SPLIT distance="1200" swimtime="00:23:25.94" />
                    <SPLIT distance="1250" swimtime="00:24:25.60" />
                    <SPLIT distance="1300" swimtime="00:25:26.51" />
                    <SPLIT distance="1350" swimtime="00:26:27.35" />
                    <SPLIT distance="1400" swimtime="00:27:27.56" />
                    <SPLIT distance="1450" swimtime="00:28:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="169" reactiontime="+98" swimtime="00:01:21.24" resultid="2855" heatid="7504" lane="2" entrytime="00:01:22.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="133" reactiontime="+95" swimtime="00:03:14.38" resultid="2856" heatid="7689" lane="2" entrytime="00:03:16.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.12" />
                    <SPLIT distance="100" swimtime="00:01:33.53" />
                    <SPLIT distance="150" swimtime="00:02:25.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="125" swimtime="00:07:05.31" resultid="2857" heatid="8046" lane="5" entrytime="00:06:59.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.34" />
                    <SPLIT distance="100" swimtime="00:01:38.79" />
                    <SPLIT distance="150" swimtime="00:02:32.56" />
                    <SPLIT distance="200" swimtime="00:03:26.52" />
                    <SPLIT distance="250" swimtime="00:04:21.16" />
                    <SPLIT distance="300" swimtime="00:05:15.94" />
                    <SPLIT distance="350" swimtime="00:06:11.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="SK Spolchemie Usti nad Labem" nation="CZE">
          <CONTACT email="benova.dana@seznam.cz" name="SK Spolchemie Usti nad Labem" phone="+420728212656" />
          <ATHLETES>
            <ATHLETE birthdate="1956-07-10" firstname="Vaclav" gender="M" lastname="Valtr" nation="CZE" license="560710" athleteid="2863">
              <RESULTS>
                <RESULT eventid="1200" points="266" reactiontime="+79" swimtime="00:00:35.14" resultid="2864" heatid="7449" lane="3" entrytime="00:00:36.20" />
                <RESULT eventid="1302" points="319" reactiontime="+85" swimtime="00:01:14.27" resultid="2865" heatid="7548" lane="4" entrytime="00:01:15.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="272" reactiontime="+87" swimtime="00:01:25.73" resultid="2866" heatid="7602" lane="1" entrytime="00:01:25.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="234" reactiontime="+88" swimtime="00:06:21.63" resultid="2867" heatid="7978" lane="2" entrytime="00:06:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.57" />
                    <SPLIT distance="100" swimtime="00:01:33.65" />
                    <SPLIT distance="150" swimtime="00:02:21.90" />
                    <SPLIT distance="200" swimtime="00:03:10.10" />
                    <SPLIT distance="250" swimtime="00:04:03.45" />
                    <SPLIT distance="300" swimtime="00:04:56.43" />
                    <SPLIT distance="350" swimtime="00:05:40.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="229" reactiontime="+77" swimtime="00:02:53.34" resultid="2868" heatid="7767" lane="4" entrytime="00:02:55.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.63" />
                    <SPLIT distance="100" swimtime="00:01:25.07" />
                    <SPLIT distance="150" swimtime="00:02:10.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="251" reactiontime="+88" swimtime="00:05:37.12" resultid="2869" heatid="8051" lane="6" entrytime="00:05:38.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                    <SPLIT distance="100" swimtime="00:01:19.37" />
                    <SPLIT distance="150" swimtime="00:02:02.05" />
                    <SPLIT distance="200" swimtime="00:02:45.21" />
                    <SPLIT distance="250" swimtime="00:03:28.10" />
                    <SPLIT distance="300" swimtime="00:04:11.69" />
                    <SPLIT distance="350" swimtime="00:04:55.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-26" firstname="Dana" gender="F" lastname="Benova" nation="CZE" license="565126" athleteid="2870">
              <RESULTS>
                <RESULT eventid="1217" points="93" reactiontime="+91" swimtime="00:04:56.94" resultid="2871" heatid="7463" lane="6" entrytime="00:04:50.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.97" />
                    <SPLIT distance="100" swimtime="00:02:24.78" />
                    <SPLIT distance="150" swimtime="00:03:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="23" reactiontime="+97" swimtime="00:07:02.08" resultid="2872" heatid="7561" lane="2" entrytime="00:06:34.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.08" />
                    <SPLIT distance="100" swimtime="00:03:06.22" />
                    <SPLIT distance="150" swimtime="00:05:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="87" swimtime="00:02:21.47" resultid="2873" heatid="7582" lane="5" entrytime="00:02:22.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="77" reactiontime="+92" swimtime="00:04:20.95" resultid="2874" heatid="7675" lane="3" entrytime="00:04:15.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.45" />
                    <SPLIT distance="100" swimtime="00:02:06.14" />
                    <SPLIT distance="150" swimtime="00:03:14.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="89" reactiontime="+80" swimtime="00:04:28.17" resultid="2875" heatid="7754" lane="3" entrytime="00:04:26.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.41" />
                    <SPLIT distance="100" swimtime="00:02:12.71" />
                    <SPLIT distance="150" swimtime="00:03:21.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="83" swimtime="00:08:58.13" resultid="2876" heatid="8019" lane="5" entrytime="00:08:46.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.92" />
                    <SPLIT distance="100" swimtime="00:02:10.43" />
                    <SPLIT distance="150" swimtime="00:03:19.66" />
                    <SPLIT distance="200" swimtime="00:04:28.63" />
                    <SPLIT distance="250" swimtime="00:05:37.47" />
                    <SPLIT distance="300" swimtime="00:06:45.32" />
                    <SPLIT distance="350" swimtime="00:07:52.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKRAS" name="Masterskrasnik" nation="POL" region="LU">
          <CONTACT city="Kraśnik" email="jurek@krasnik.info" name="Michalczyk Jerzy" phone="601698977" state="LUB" street="Żwirki i Wigury 2" zip="23-210" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-04" firstname="Mirosław" gender="M" lastname="Leszczyński" nation="POL" athleteid="2878">
              <RESULTS>
                <RESULT eventid="1234" points="295" reactiontime="+90" swimtime="00:03:01.20" resultid="2879" heatid="7480" lane="4" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:26.95" />
                    <SPLIT distance="150" swimtime="00:02:13.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="307" reactiontime="+93" swimtime="00:01:22.37" resultid="2880" heatid="7604" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MALOD" name="Masters Łódź" nation="POL" region="LO">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="TRUDNOS RAFAŁ" phone="604184311" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Marcin" gender="M" lastname="Strąkowski" nation="POL" athleteid="2882">
              <RESULTS>
                <RESULT eventid="1075" points="343" reactiontime="+84" swimtime="00:00:28.99" resultid="2883" heatid="7370" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1268" points="278" reactiontime="+89" swimtime="00:01:08.85" resultid="2884" heatid="7513" lane="3" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="310" reactiontime="+84" swimtime="00:00:37.27" resultid="2885" heatid="7807" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="2886">
              <RESULTS>
                <RESULT eventid="1075" points="294" reactiontime="+97" swimtime="00:00:30.52" resultid="2887" heatid="7358" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1109" points="215" reactiontime="+97" swimtime="00:03:03.54" resultid="2888" heatid="7397" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:02:19.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="219" swimtime="00:03:19.90" resultid="2889" heatid="7476" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:34.21" />
                    <SPLIT distance="150" swimtime="00:02:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="255" reactiontime="+98" swimtime="00:01:19.96" resultid="2890" heatid="7545" lane="3" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="226" reactiontime="+101" swimtime="00:01:31.24" resultid="2891" heatid="7603" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="2893" heatid="7767" lane="3" entrytime="00:02:55.00" />
                <RESULT eventid="1662" points="269" reactiontime="+93" swimtime="00:00:39.09" resultid="2894" heatid="7799" lane="4" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Jakub" gender="M" lastname="Gryczyński" nation="POL" athleteid="2895">
              <RESULTS>
                <RESULT eventid="1075" points="300" reactiontime="+88" swimtime="00:00:30.30" resultid="2896" heatid="7363" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="2897" heatid="7545" lane="4" entrytime="00:01:22.00" />
                <RESULT eventid="1402" points="265" reactiontime="+84" swimtime="00:01:26.47" resultid="2898" heatid="7601" lane="1" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="280" swimtime="00:00:38.57" resultid="2899" heatid="7800" lane="5" entrytime="00:00:38.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="2900">
              <RESULTS>
                <RESULT eventid="1075" points="431" reactiontime="+95" swimtime="00:00:26.87" resultid="2901" heatid="7377" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1268" points="373" swimtime="00:01:02.41" resultid="2902" heatid="7516" lane="5" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="348" reactiontime="+96" swimtime="00:00:30.98" resultid="2903" heatid="7636" lane="6" entrytime="00:00:31.71" />
                <RESULT eventid="1662" points="388" swimtime="00:00:34.61" resultid="2904" heatid="7807" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Rafał" gender="M" lastname="Trudnos" nation="POL" athleteid="2905">
              <RESULTS>
                <RESULT eventid="1075" points="417" reactiontime="+77" swimtime="00:00:27.17" resultid="2906" heatid="7368" lane="4" entrytime="00:00:28.50" />
                <RESULT eventid="1234" points="393" reactiontime="+79" swimtime="00:02:44.69" resultid="2907" heatid="7482" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="150" swimtime="00:02:01.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="411" swimtime="00:01:14.74" resultid="2908" heatid="7608" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="415" reactiontime="+77" swimtime="00:00:29.21" resultid="2909" heatid="7640" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1662" points="434" swimtime="00:00:33.33" resultid="2910" heatid="7809" lane="5" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" athleteid="2911">
              <RESULTS>
                <RESULT eventid="1075" points="448" reactiontime="+81" swimtime="00:00:26.52" resultid="2912" heatid="7378" lane="4" entrytime="00:00:25.80" />
                <RESULT eventid="1268" points="419" reactiontime="+82" swimtime="00:01:00.03" resultid="2913" heatid="7520" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="382" reactiontime="+76" swimtime="00:00:30.04" resultid="2914" heatid="7643" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="2915" heatid="7702" lane="1" entrytime="00:02:15.00" />
                <RESULT eventid="1594" points="372" reactiontime="+88" swimtime="00:01:07.37" resultid="2916" heatid="7748" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" athleteid="2917">
              <RESULTS>
                <RESULT eventid="1075" points="307" reactiontime="+87" swimtime="00:00:30.07" resultid="2918" heatid="7366" lane="1" entrytime="00:00:29.27" />
                <RESULT eventid="1302" points="254" reactiontime="+82" swimtime="00:01:20.14" resultid="2919" heatid="7546" lane="1" entrytime="00:01:20.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="268" reactiontime="+84" swimtime="00:00:39.13" resultid="2920" heatid="7799" lane="2" entrytime="00:00:39.63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Kornel" gender="M" lastname="Pintara" nation="POL" athleteid="2921">
              <RESULTS>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="2922" heatid="7451" lane="2" entrytime="00:00:34.50" />
                <RESULT eventid="1302" points="342" reactiontime="+88" swimtime="00:01:12.58" resultid="2923" heatid="7553" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="321" reactiontime="+85" swimtime="00:00:31.82" resultid="2924" heatid="7639" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1504" points="310" reactiontime="+86" swimtime="00:02:26.82" resultid="2925" heatid="7699" lane="4" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:47.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="267" reactiontime="+90" swimtime="00:01:15.25" resultid="2926" heatid="7744" lane="6" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="2927" heatid="7800" lane="2" entrytime="00:00:38.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="2928">
              <RESULTS>
                <RESULT eventid="1075" points="355" reactiontime="+84" swimtime="00:00:28.66" resultid="2929" heatid="7364" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1165" points="284" reactiontime="+90" swimtime="00:21:32.03" resultid="2930" heatid="7913" lane="4" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:53.30" />
                    <SPLIT distance="200" swimtime="00:02:33.96" />
                    <SPLIT distance="250" swimtime="00:03:16.36" />
                    <SPLIT distance="300" swimtime="00:03:59.64" />
                    <SPLIT distance="350" swimtime="00:04:42.85" />
                    <SPLIT distance="400" swimtime="00:05:26.85" />
                    <SPLIT distance="450" swimtime="00:06:11.01" />
                    <SPLIT distance="500" swimtime="00:06:54.85" />
                    <SPLIT distance="550" swimtime="00:07:38.99" />
                    <SPLIT distance="600" swimtime="00:08:23.72" />
                    <SPLIT distance="650" swimtime="00:09:07.78" />
                    <SPLIT distance="700" swimtime="00:09:51.78" />
                    <SPLIT distance="750" swimtime="00:10:36.81" />
                    <SPLIT distance="800" swimtime="00:11:20.77" />
                    <SPLIT distance="850" swimtime="00:12:05.14" />
                    <SPLIT distance="900" swimtime="00:12:49.46" />
                    <SPLIT distance="950" swimtime="00:13:33.84" />
                    <SPLIT distance="1000" swimtime="00:14:18.07" />
                    <SPLIT distance="1050" swimtime="00:15:01.99" />
                    <SPLIT distance="1100" swimtime="00:15:46.35" />
                    <SPLIT distance="1150" swimtime="00:16:29.67" />
                    <SPLIT distance="1200" swimtime="00:17:13.38" />
                    <SPLIT distance="1250" swimtime="00:17:57.03" />
                    <SPLIT distance="1300" swimtime="00:18:40.84" />
                    <SPLIT distance="1350" swimtime="00:19:24.57" />
                    <SPLIT distance="1400" swimtime="00:20:08.03" />
                    <SPLIT distance="1450" swimtime="00:20:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="334" reactiontime="+85" swimtime="00:01:04.77" resultid="2931" heatid="7515" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M-12 - Dotkniecie jedną reką sciany nawrotowej w czasie zakonczenia wyścigu" eventid="1436" status="DSQ" swimtime="00:00:31.39" resultid="2932" heatid="7640" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="2933" heatid="7700" lane="3" entrytime="00:02:20.00" />
                <RESULT eventid="1710" points="292" reactiontime="+81" swimtime="00:05:20.37" resultid="2934" heatid="8053" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="150" swimtime="00:01:49.97" />
                    <SPLIT distance="200" swimtime="00:02:30.20" />
                    <SPLIT distance="250" swimtime="00:03:12.19" />
                    <SPLIT distance="300" swimtime="00:03:55.03" />
                    <SPLIT distance="350" swimtime="00:04:38.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="Jakub" gender="M" lastname="Sidorowicz" nation="POL" athleteid="2935">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2936" heatid="7395" lane="5" entrytime="00:03:24.10" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="2937" heatid="7447" lane="4" entrytime="00:00:39.70" />
                <RESULT eventid="1302" points="191" reactiontime="+92" swimtime="00:01:28.03" resultid="2938" heatid="7544" lane="1" entrytime="00:01:27.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="200" reactiontime="+91" swimtime="00:01:34.95" resultid="2939" heatid="7597" lane="4" entrytime="00:01:36.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="2940" heatid="7663" lane="4" entrytime="00:01:29.55" />
                <RESULT eventid="1662" points="229" swimtime="00:00:41.22" resultid="2941" heatid="7799" lane="5" entrytime="00:00:39.95" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Robert" gender="M" lastname="Lesiak" nation="POL" athleteid="2942">
              <RESULTS>
                <RESULT eventid="1075" points="314" reactiontime="+97" swimtime="00:00:29.85" resultid="2943" heatid="7355" lane="3" entrytime="00:00:33.33" />
                <RESULT eventid="1109" points="213" reactiontime="+78" swimtime="00:03:04.15" resultid="2944" heatid="7396" lane="4" entrytime="00:03:05.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="150" swimtime="00:02:22.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="2945" heatid="7449" lane="2" entrytime="00:00:36.84" />
                <RESULT eventid="1302" points="217" reactiontime="+97" swimtime="00:01:24.39" resultid="2946" heatid="7546" lane="6" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="221" reactiontime="+73" swimtime="00:01:20.92" resultid="2947" heatid="7665" lane="2" entrytime="00:01:20.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="2948" heatid="7983" lane="5" entrytime="00:06:59.18" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="2949" heatid="7743" lane="5" entrytime="00:01:20.02" />
                <RESULT eventid="1710" points="190" reactiontime="+106" swimtime="00:06:09.52" resultid="2950" heatid="8047" lane="1" entrytime="00:06:30.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                    <SPLIT distance="150" swimtime="00:02:06.56" />
                    <SPLIT distance="200" swimtime="00:02:53.18" />
                    <SPLIT distance="250" swimtime="00:03:42.14" />
                    <SPLIT distance="300" swimtime="00:04:32.95" />
                    <SPLIT distance="350" swimtime="00:05:23.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="Konrad" gender="M" lastname="Hasik" nation="POL" athleteid="2951">
              <RESULTS>
                <RESULT eventid="1075" points="442" reactiontime="+82" swimtime="00:00:26.64" resultid="2952" heatid="7372" lane="6" entrytime="00:00:27.50" />
                <RESULT eventid="1109" points="392" reactiontime="+89" swimtime="00:02:30.29" resultid="2953" heatid="7403" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:51.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="386" swimtime="00:02:45.71" resultid="2954" heatid="7482" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:20.36" />
                    <SPLIT distance="150" swimtime="00:02:04.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="2955" heatid="7554" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="2956" heatid="7606" lane="2" entrytime="00:01:20.00" />
                <RESULT eventid="1470" points="429" reactiontime="+63" swimtime="00:01:04.87" resultid="2957" heatid="7670" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="353" reactiontime="+63" swimtime="00:02:30.14" resultid="2959" heatid="7772" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:49.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="2960" heatid="7807" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Marcin" gender="M" lastname="Babuchowski" nation="POL" athleteid="2961">
              <RESULTS>
                <RESULT eventid="1075" points="579" swimtime="00:00:24.35" resultid="2962" heatid="7381" lane="5" entrytime="00:00:24.00" />
                <RESULT eventid="1268" points="609" reactiontime="+73" swimtime="00:00:53.00" resultid="2963" heatid="7525" lane="2" entrytime="00:00:51.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="638" reactiontime="+71" swimtime="00:00:25.31" resultid="2964" heatid="7647" lane="4" entrytime="00:00:24.48" />
                <RESULT eventid="1504" points="586" reactiontime="+77" swimtime="00:01:58.74" resultid="2965" heatid="7706" lane="2" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                    <SPLIT distance="100" swimtime="00:00:57.04" />
                    <SPLIT distance="150" swimtime="00:01:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1594" points="643" reactiontime="+74" swimtime="00:00:56.16" resultid="2966" heatid="7752" lane="3" entrytime="00:00:54.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Maciej" gender="M" lastname="Machnicki" nation="POL" athleteid="2967">
              <RESULTS>
                <RESULT eventid="1075" points="275" reactiontime="+91" swimtime="00:00:31.19" resultid="2968" heatid="7361" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="2969" heatid="7450" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1268" points="204" reactiontime="+88" swimtime="00:01:16.31" resultid="2970" heatid="7506" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="2971" heatid="7630" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Łukasz" gender="M" lastname="Maślak" nation="POL" athleteid="2972">
              <RESULTS>
                <RESULT eventid="1075" points="102" reactiontime="+120" swimtime="00:00:43.36" resultid="2973" heatid="7348" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="2974" heatid="7443" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="2975" heatid="7501" lane="5" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Damian" gender="M" lastname="Karkusiński" nation="POL" athleteid="2976">
              <RESULTS>
                <RESULT eventid="1075" points="317" reactiontime="+98" swimtime="00:00:29.76" resultid="2977" heatid="7366" lane="3" entrytime="00:00:29.05" />
                <RESULT eventid="1200" points="264" reactiontime="+61" swimtime="00:00:35.23" resultid="2978" heatid="7452" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1470" points="226" reactiontime="+64" swimtime="00:01:20.26" resultid="2979" heatid="7668" lane="5" entrytime="00:01:14.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Artur" gender="M" lastname="Frąckowiak" nation="POL" athleteid="2980">
              <RESULTS>
                <RESULT eventid="1075" points="351" reactiontime="+93" swimtime="00:00:28.76" resultid="2981" heatid="7364" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1268" points="336" swimtime="00:01:04.62" resultid="2982" heatid="7509" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="325" reactiontime="+88" swimtime="00:01:13.77" resultid="2983" heatid="7545" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="336" reactiontime="+84" swimtime="00:00:31.34" resultid="2984" heatid="7634" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1662" points="333" reactiontime="+76" swimtime="00:00:36.40" resultid="2985" heatid="7798" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-01" firstname="Łukasz" gender="M" lastname="Furman" nation="POL" athleteid="8062">
              <RESULTS>
                <RESULT eventid="1628" points="519" status="EXH" swimtime="00:02:11.99" resultid="8063" heatid="7770" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1528" points="473" reactiontime="+88" swimtime="00:01:43.60" resultid="2986" heatid="7716" lane="1" entrytime="00:01:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.94" />
                    <SPLIT distance="100" swimtime="00:00:53.35" />
                    <SPLIT distance="150" swimtime="00:01:19.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2961" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="2911" number="2" reactiontime="+15" />
                    <RELAYPOSITION athleteid="2900" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="2951" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1528" points="378" reactiontime="+78" swimtime="00:01:51.66" resultid="2987" heatid="7714" lane="3" entrytime="00:01:51.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                    <SPLIT distance="100" swimtime="00:00:56.00" />
                    <SPLIT distance="150" swimtime="00:01:24.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2905" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="2928" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="2980" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="2921" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1528" points="300" reactiontime="+96" swimtime="00:02:00.61" resultid="2988" heatid="7714" lane="2" entrytime="00:01:51.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                    <SPLIT distance="100" swimtime="00:01:01.19" />
                    <SPLIT distance="150" swimtime="00:01:31.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2942" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="2917" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2976" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2882" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1528" points="285" swimtime="00:02:02.66" resultid="2989" heatid="7712" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="100" swimtime="00:01:00.20" />
                    <SPLIT distance="150" swimtime="00:01:31.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2886" number="1" />
                    <RELAYPOSITION athleteid="2895" number="2" />
                    <RELAYPOSITION athleteid="2967" number="3" />
                    <RELAYPOSITION athleteid="2935" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1377" points="525" reactiontime="+64" swimtime="00:01:53.75" resultid="2990" heatid="7934" lane="4" entrytime="00:01:54.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                    <SPLIT distance="100" swimtime="00:01:02.91" />
                    <SPLIT distance="150" swimtime="00:01:27.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2951" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2905" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="2961" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="2911" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1377" points="343" reactiontime="+65" swimtime="00:02:11.13" resultid="2991" heatid="7933" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:12.87" />
                    <SPLIT distance="150" swimtime="00:01:44.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2976" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2895" number="2" />
                    <RELAYPOSITION athleteid="2921" number="3" />
                    <RELAYPOSITION athleteid="2900" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="1377" points="308" reactiontime="+79" swimtime="00:02:15.85" resultid="2992" heatid="7933" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:13.31" />
                    <SPLIT distance="150" swimtime="00:01:44.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2928" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2917" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2942" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2980" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1377" points="248" reactiontime="+72" swimtime="00:02:25.97" resultid="2993" heatid="7931" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:19.01" />
                    <SPLIT distance="150" swimtime="00:01:54.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2935" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2967" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2886" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="2882" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ZKS DRZONK" name="ZKS Drzonków" nation="POL" region="LBS">
          <CONTACT city="Zielona Góra" email="wojtek696@gmail.com" name="Barta Piotr" phone="602347348" state="LUBUS" street="Wyszyńskiego" zip="65-001" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-18" firstname="Piotr" gender="M" lastname="Barta" nation="POL" athleteid="3030">
              <RESULTS>
                <RESULT eventid="1234" points="451" reactiontime="+91" swimtime="00:02:37.34" resultid="3031" heatid="7484" lane="6" entrytime="00:02:40.00" entrycourse="SCY">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:01:55.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="3032" heatid="7553" lane="4" entrytime="00:01:10.00" entrycourse="SCM" />
                <RESULT eventid="1402" points="446" reactiontime="+90" swimtime="00:01:12.74" resultid="3033" heatid="7609" lane="4" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="373" reactiontime="+99" swimtime="00:05:26.97" resultid="3034" heatid="7982" lane="6" entrytime="00:05:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                    <SPLIT distance="150" swimtime="00:01:58.13" />
                    <SPLIT distance="200" swimtime="00:02:43.36" />
                    <SPLIT distance="250" swimtime="00:03:26.70" />
                    <SPLIT distance="300" swimtime="00:04:10.54" />
                    <SPLIT distance="350" swimtime="00:04:49.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="452" reactiontime="+86" swimtime="00:00:32.88" resultid="3035" heatid="7811" lane="1" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1710" points="429" reactiontime="+96" swimtime="00:04:41.98" resultid="3036" heatid="8056" lane="4" entrytime="00:04:44.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                    <SPLIT distance="150" swimtime="00:01:43.34" />
                    <SPLIT distance="200" swimtime="00:02:18.64" />
                    <SPLIT distance="250" swimtime="00:02:53.19" />
                    <SPLIT distance="300" swimtime="00:03:28.74" />
                    <SPLIT distance="350" swimtime="00:04:04.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Start Poznań" nation="POL" region="WIE">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" phone="512111513" street="Os. Batorego 8/67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1967-02-22" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="3038">
              <RESULTS>
                <RESULT eventid="1075" points="460" swimtime="00:00:26.28" resultid="3039" heatid="7375" lane="5" entrytime="00:00:26.80" entrycourse="SCM" />
                <RESULT eventid="1109" points="417" reactiontime="+75" swimtime="00:02:27.33" resultid="3040" heatid="7404" lane="4" entrytime="00:02:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:53.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="478" reactiontime="+56" swimtime="00:00:57.47" resultid="3041" heatid="7522" lane="3" entrytime="00:00:58.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="432" reactiontime="+73" swimtime="00:01:07.12" resultid="3042" heatid="7557" lane="6" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="448" reactiontime="+58" swimtime="00:02:09.81" resultid="3043" heatid="7703" lane="3" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:03.26" />
                    <SPLIT distance="150" swimtime="00:01:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="371" reactiontime="+79" swimtime="00:05:27.54" resultid="3044" heatid="7980" lane="1" entrytime="00:05:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:12.97" />
                    <SPLIT distance="150" swimtime="00:01:55.32" />
                    <SPLIT distance="200" swimtime="00:02:37.89" />
                    <SPLIT distance="250" swimtime="00:03:26.62" />
                    <SPLIT distance="300" swimtime="00:04:14.95" />
                    <SPLIT distance="350" swimtime="00:04:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="438" swimtime="00:04:40.16" resultid="3045" heatid="8056" lane="5" entrytime="00:04:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:44.06" />
                    <SPLIT distance="200" swimtime="00:02:20.51" />
                    <SPLIT distance="250" swimtime="00:02:55.80" />
                    <SPLIT distance="300" swimtime="00:03:30.94" />
                    <SPLIT distance="350" swimtime="00:04:06.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-26" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="3046">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="3047" heatid="7370" lane="6" entrytime="00:00:28.01" entrycourse="SCM" />
                <RESULT eventid="1165" points="351" reactiontime="+109" swimtime="00:20:04.58" resultid="3048" heatid="7913" lane="2" entrytime="00:22:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:52.66" />
                    <SPLIT distance="200" swimtime="00:02:32.83" />
                    <SPLIT distance="250" swimtime="00:03:13.53" />
                    <SPLIT distance="300" swimtime="00:03:54.15" />
                    <SPLIT distance="350" swimtime="00:04:35.64" />
                    <SPLIT distance="400" swimtime="00:05:16.78" />
                    <SPLIT distance="450" swimtime="00:05:57.29" />
                    <SPLIT distance="500" swimtime="00:06:37.52" />
                    <SPLIT distance="550" swimtime="00:07:18.06" />
                    <SPLIT distance="600" swimtime="00:07:58.20" />
                    <SPLIT distance="650" swimtime="00:08:38.76" />
                    <SPLIT distance="700" swimtime="00:09:19.68" />
                    <SPLIT distance="750" swimtime="00:10:00.22" />
                    <SPLIT distance="800" swimtime="00:10:40.77" />
                    <SPLIT distance="850" swimtime="00:11:21.22" />
                    <SPLIT distance="900" swimtime="00:12:01.79" />
                    <SPLIT distance="950" swimtime="00:12:42.14" />
                    <SPLIT distance="1000" swimtime="00:13:22.19" />
                    <SPLIT distance="1050" swimtime="00:14:02.80" />
                    <SPLIT distance="1100" swimtime="00:14:43.31" />
                    <SPLIT distance="1150" swimtime="00:15:23.39" />
                    <SPLIT distance="1200" swimtime="00:16:03.94" />
                    <SPLIT distance="1250" swimtime="00:16:44.47" />
                    <SPLIT distance="1300" swimtime="00:17:24.97" />
                    <SPLIT distance="1350" swimtime="00:18:05.29" />
                    <SPLIT distance="1400" swimtime="00:18:45.85" />
                    <SPLIT distance="1450" swimtime="00:19:26.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="3049" heatid="7454" lane="1" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="3050" heatid="7520" lane="1" entrytime="00:01:01.00" entrycourse="SCM" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="3051" heatid="7670" lane="5" entrytime="00:01:10.00" entrycourse="SCM" />
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="3052" heatid="7771" lane="1" entrytime="00:02:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Takas" nation="LTU">
          <CONTACT city="Kaunas" email="abicka@takas.lt" internet="www.klubastakas.lt" name="Arlandas Juodeska" phone="+37068687934" street="Lentvario g. 19" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1961-12-26" firstname="Arlandas" gender="M" lastname="juodeska" nation="LTU" athleteid="3055">
              <RESULTS>
                <RESULT eventid="1075" points="328" reactiontime="+81" swimtime="00:00:29.42" resultid="3056" heatid="7367" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1302" points="327" reactiontime="+84" swimtime="00:01:13.67" resultid="3058" heatid="7549" lane="3" entrytime="00:01:14.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="313" reactiontime="+81" swimtime="00:01:21.87" resultid="3059" heatid="7605" lane="6" entrytime="00:01:21.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="276" reactiontime="+66" swimtime="00:01:15.12" resultid="3060" heatid="7668" lane="1" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="244" reactiontime="+65" swimtime="00:02:49.64" resultid="3061" heatid="7768" lane="6" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                    <SPLIT distance="100" swimtime="00:01:21.43" />
                    <SPLIT distance="150" swimtime="00:02:05.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="323" reactiontime="+80" swimtime="00:00:36.78" resultid="3062" heatid="7805" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1200" points="328" reactiontime="+67" swimtime="00:00:32.77" resultid="6424" heatid="7453" lane="5" entrytime="00:00:33.28" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-11-16" firstname="Violeta" gender="F" lastname="povilaitiene" nation="LTU" athleteid="6075">
              <RESULTS>
                <RESULT eventid="1058" points="91" swimtime="00:00:51.69" resultid="6076" heatid="7333" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1217" points="103" reactiontime="+125" swimtime="00:04:46.61" resultid="6077" heatid="7463" lane="2" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.04" />
                    <SPLIT distance="100" swimtime="00:03:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="6078" heatid="7583" lane="1" entrytime="00:02:10.00" />
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="6080" heatid="7755" lane="1" entrytime="00:04:15.00" />
                <RESULT eventid="1645" points="114" reactiontime="+117" swimtime="00:00:59.24" resultid="6081" heatid="7778" lane="1" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-14" firstname="Violeta" gender="F" lastname="Penkauskaite" nation="LTU" athleteid="6082">
              <RESULTS>
                <RESULT eventid="1058" points="111" reactiontime="+92" swimtime="00:00:48.34" resultid="6083" heatid="7333" lane="6" entrytime="00:00:59.00" />
                <RESULT eventid="1092" points="124" swimtime="00:04:09.61" resultid="6084" heatid="7383" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.16" />
                    <SPLIT distance="100" swimtime="00:02:01.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="89" swimtime="00:01:53.88" resultid="6085" heatid="7487" lane="5" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="114" reactiontime="+99" swimtime="00:01:59.06" resultid="6086" heatid="7527" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="6087" heatid="7649" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:31.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="104" reactiontime="+71" swimtime="00:04:15.05" resultid="6088" heatid="7754" lane="4" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:05.07" />
                    <SPLIT distance="100" swimtime="00:03:10.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="106" swimtime="00:00:54.20" resultid="7849" heatid="7431" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-10-18" firstname="Ramune" gender="F" lastname="ivanauskaite" nation="LTU" athleteid="6089">
              <RESULTS>
                <RESULT eventid="1092" points="307" reactiontime="+91" swimtime="00:03:04.67" resultid="6090" heatid="7387" lane="1" entrytime="00:03:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                    <SPLIT distance="100" swimtime="00:01:28.52" />
                    <SPLIT distance="150" swimtime="00:02:21.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="247" swimtime="00:00:40.91" resultid="6091" heatid="7437" lane="2" entrytime="00:00:39.70" />
                <RESULT eventid="1217" points="297" reactiontime="+86" swimtime="00:03:21.68" resultid="6092" heatid="7466" lane="6" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                    <SPLIT distance="100" swimtime="00:01:37.80" />
                    <SPLIT distance="150" swimtime="00:02:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="280" reactiontime="+88" swimtime="00:01:35.77" resultid="6093" heatid="7588" lane="2" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="247" reactiontime="+82" swimtime="00:01:27.92" resultid="6094" heatid="7653" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="270" reactiontime="+84" swimtime="00:03:05.53" resultid="6095" heatid="7758" lane="4" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                    <SPLIT distance="100" swimtime="00:01:30.21" />
                    <SPLIT distance="150" swimtime="00:02:18.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-04-12" firstname="Aleksandra" gender="F" lastname="yliene" nation="LTU" athleteid="6096">
              <RESULTS>
                <RESULT eventid="1058" points="141" swimtime="00:00:44.61" resultid="6097" heatid="7334" lane="5" entrytime="00:00:44.00" />
                <RESULT eventid="1183" points="120" swimtime="00:00:52.02" resultid="6098" heatid="7433" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1251" points="116" reactiontime="+125" swimtime="00:01:44.54" resultid="6099" heatid="7488" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="104" reactiontime="+85" swimtime="00:01:57.09" resultid="6100" heatid="7650" lane="1" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="89" reactiontime="+92" swimtime="00:04:27.97" resultid="6101" heatid="7755" lane="2" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.52" />
                    <SPLIT distance="100" swimtime="00:02:11.92" />
                    <SPLIT distance="150" swimtime="00:03:22.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="TKKF Koszalin Masters" nation="POL">
          <CONTACT city="Koszalin" email="jakubkielar3@gmail.com" name="Kielar Jakub" phone="693193137" state="ZACH" street="Holenderska 6" zip="75-430" />
          <ATHLETES>
            <ATHLETE birthdate="1974-01-21" firstname="Jakub" gender="M" lastname="Kielar" nation="POL" athleteid="3071">
              <RESULTS>
                <RESULT eventid="1075" points="423" reactiontime="+74" swimtime="00:00:27.03" resultid="5571" heatid="7375" lane="3" entrytime="00:00:26.50" entrycourse="SCM" />
                <RESULT eventid="1109" points="342" reactiontime="+79" swimtime="00:02:37.36" resultid="5572" heatid="7405" lane="6" entrytime="00:02:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:13.36" />
                    <SPLIT distance="150" swimtime="00:02:01.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="5573" heatid="7500" lane="4" />
                <RESULT eventid="1302" points="430" reactiontime="+78" swimtime="00:01:07.24" resultid="5574" heatid="7556" lane="2" entrytime="00:01:07.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="431" reactiontime="+77" swimtime="00:00:28.86" resultid="5575" heatid="7643" lane="2" entrytime="00:00:28.38" entrycourse="SCM" />
                <RESULT eventid="1594" points="363" reactiontime="+93" swimtime="00:01:07.94" resultid="5577" heatid="7749" lane="4" entrytime="00:01:07.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="375" reactiontime="+87" swimtime="00:00:35.01" resultid="5578" heatid="7808" lane="1" entrytime="00:00:34.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-06-12" firstname="Joanna" gender="F" lastname="Stankiewicz - Majkowska" nation="POL" athleteid="3080">
              <RESULTS>
                <RESULT eventid="1058" points="209" reactiontime="+88" swimtime="00:00:39.12" resultid="5579" heatid="7336" lane="4" entrytime="00:00:37.50" entrycourse="SCM" />
                <RESULT eventid="1092" points="198" reactiontime="+83" swimtime="00:03:33.42" resultid="5580" heatid="7384" lane="3" entrytime="00:03:35.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="100" swimtime="00:01:40.36" />
                    <SPLIT distance="150" swimtime="00:02:39.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="164" reactiontime="+83" swimtime="00:00:46.91" resultid="5581" heatid="7434" lane="5" entrytime="00:00:45.20" entrycourse="SCM" />
                <RESULT eventid="1285" points="208" swimtime="00:01:37.43" resultid="5582" heatid="7529" lane="5" entrytime="00:01:32.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="179" reactiontime="+92" swimtime="00:01:51.11" resultid="5583" heatid="7586" lane="2" entrytime="00:01:42.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="187" reactiontime="+90" swimtime="00:00:50.33" resultid="5584" heatid="7781" lane="2" entrytime="00:00:47.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-02-16" firstname="Katarzyna" gender="F" lastname="Gudaniec" nation="POL" athleteid="3087">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="5585" heatid="7337" lane="6" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1148" points="416" reactiontime="+58" swimtime="00:10:48.76" resultid="5586" heatid="7905" lane="3" entrytime="00:10:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:52.59" />
                    <SPLIT distance="200" swimtime="00:02:32.85" />
                    <SPLIT distance="250" swimtime="00:03:13.32" />
                    <SPLIT distance="300" swimtime="00:03:53.92" />
                    <SPLIT distance="350" swimtime="00:04:34.76" />
                    <SPLIT distance="400" swimtime="00:05:16.01" />
                    <SPLIT distance="450" swimtime="00:05:57.34" />
                    <SPLIT distance="500" swimtime="00:06:39.01" />
                    <SPLIT distance="550" swimtime="00:07:20.50" />
                    <SPLIT distance="600" swimtime="00:08:01.92" />
                    <SPLIT distance="650" swimtime="00:08:43.50" />
                    <SPLIT distance="700" swimtime="00:09:25.53" />
                    <SPLIT distance="750" swimtime="00:10:07.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="382" reactiontime="+52" swimtime="00:01:19.55" resultid="5587" heatid="7531" lane="3" entrytime="00:01:25.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="398" swimtime="00:02:31.02" resultid="5588" heatid="7683" lane="5" entrytime="00:02:31.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:10.38" />
                    <SPLIT distance="150" swimtime="00:01:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="401" swimtime="00:05:18.42" resultid="5589" heatid="8024" lane="5" entrytime="00:05:20.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:13.24" />
                    <SPLIT distance="150" swimtime="00:01:52.45" />
                    <SPLIT distance="200" swimtime="00:02:33.42" />
                    <SPLIT distance="250" swimtime="00:03:14.82" />
                    <SPLIT distance="300" swimtime="00:03:56.55" />
                    <SPLIT distance="350" swimtime="00:04:37.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-21" firstname="Janusz" gender="M" lastname="Dudziński" nation="POL" athleteid="3093">
              <RESULTS>
                <RESULT eventid="1075" points="314" reactiontime="+90" swimtime="00:00:29.85" resultid="5590" heatid="7369" lane="2" entrytime="00:00:28.20" entrycourse="SCM" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="5592" heatid="7481" lane="3" entrytime="00:02:54.00" entrycourse="SCM" />
                <RESULT eventid="1302" points="238" reactiontime="+89" swimtime="00:01:21.80" resultid="5593" heatid="7550" lane="1" entrytime="00:01:14.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="5594" heatid="7637" lane="4" entrytime="00:00:30.95" entrycourse="SCM" />
                <RESULT eventid="1662" points="288" reactiontime="+87" swimtime="00:00:38.21" resultid="5595" heatid="7806" lane="1" entrytime="00:00:35.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-08-26" firstname="Dorota" gender="F" lastname="Gudaniec" nation="POL" athleteid="3100">
              <RESULTS>
                <RESULT eventid="1058" points="236" swimtime="00:00:37.62" resultid="5596" heatid="7336" lane="5" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1148" points="219" reactiontime="+105" swimtime="00:13:22.70" resultid="5597" heatid="7904" lane="1" entrytime="00:12:54.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                    <SPLIT distance="100" swimtime="00:01:31.45" />
                    <SPLIT distance="150" swimtime="00:02:22.03" />
                    <SPLIT distance="200" swimtime="00:03:13.13" />
                    <SPLIT distance="250" swimtime="00:04:04.28" />
                    <SPLIT distance="300" swimtime="00:04:55.33" />
                    <SPLIT distance="350" swimtime="00:05:46.65" />
                    <SPLIT distance="400" swimtime="00:06:37.80" />
                    <SPLIT distance="450" swimtime="00:07:28.64" />
                    <SPLIT distance="500" swimtime="00:08:19.95" />
                    <SPLIT distance="550" swimtime="00:09:11.10" />
                    <SPLIT distance="600" swimtime="00:10:02.28" />
                    <SPLIT distance="650" swimtime="00:10:53.23" />
                    <SPLIT distance="700" swimtime="00:11:43.97" />
                    <SPLIT distance="750" swimtime="00:12:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="206" reactiontime="+101" swimtime="00:03:47.59" resultid="5598" heatid="7465" lane="3" entrytime="00:03:41.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.56" />
                    <SPLIT distance="100" swimtime="00:01:49.71" />
                    <SPLIT distance="150" swimtime="00:02:49.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="232" reactiontime="+92" swimtime="00:01:33.89" resultid="5599" heatid="7529" lane="4" entrytime="00:01:30.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="5600" heatid="7586" lane="1" entrytime="00:01:43.50" entrycourse="SCM" />
                <RESULT eventid="1487" points="193" reactiontime="+94" swimtime="00:03:12.04" resultid="5601" heatid="7678" lane="2" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:30.58" />
                    <SPLIT distance="150" swimtime="00:02:21.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5602" heatid="7780" lane="3" entrytime="00:00:48.30" entrycourse="SCM" />
                <RESULT eventid="1693" points="213" reactiontime="+101" swimtime="00:06:32.90" resultid="5603" heatid="8021" lane="2" entrytime="00:06:24.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:30.32" />
                    <SPLIT distance="150" swimtime="00:02:20.19" />
                    <SPLIT distance="200" swimtime="00:03:10.94" />
                    <SPLIT distance="250" swimtime="00:04:01.67" />
                    <SPLIT distance="300" swimtime="00:04:52.92" />
                    <SPLIT distance="350" swimtime="00:05:43.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-20" firstname="Joanna" gender="F" lastname="Wojciechowska" nation="POL" athleteid="3109">
              <RESULTS>
                <RESULT eventid="1058" points="203" reactiontime="+85" swimtime="00:00:39.56" resultid="5604" heatid="7336" lane="3" entrytime="00:00:37.20" entrycourse="SCM" />
                <RESULT eventid="1251" points="186" reactiontime="+86" swimtime="00:01:29.22" resultid="5605" heatid="7491" lane="3" entrytime="00:01:22.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="5606" heatid="7584" lane="1" entrytime="00:01:53.30" entrycourse="SCM" />
                <RESULT eventid="1487" status="DNS" swimtime="00:00:00.00" resultid="5607" heatid="7678" lane="5" entrytime="00:03:10.00" entrycourse="SCM" />
                <RESULT eventid="1645" points="192" reactiontime="+82" swimtime="00:00:49.89" resultid="5608" heatid="7780" lane="4" entrytime="00:00:48.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-07-05" firstname="Krzysztof" gender="M" lastname="Stefański" nation="POL" athleteid="3115">
              <RESULTS>
                <RESULT eventid="1075" points="354" reactiontime="+87" swimtime="00:00:28.68" resultid="5609" heatid="7373" lane="1" entrytime="00:00:27.10" entrycourse="SCM" />
                <RESULT eventid="1268" points="322" reactiontime="+91" swimtime="00:01:05.50" resultid="5610" heatid="7517" lane="1" entrytime="00:01:03.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="247" reactiontime="+83" swimtime="00:01:28.56" resultid="5611" heatid="7593" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="5612" heatid="7638" lane="6" entrytime="00:00:30.80" entrycourse="SCM" />
                <RESULT eventid="1662" points="272" reactiontime="+86" swimtime="00:00:38.96" resultid="5613" heatid="7806" lane="6" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-08" firstname="Dawid" gender="M" lastname="Borus" nation="POL" athleteid="5614">
              <RESULTS>
                <RESULT eventid="1200" points="321" reactiontime="+77" swimtime="00:00:32.99" resultid="5615" heatid="7453" lane="4" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1302" points="341" reactiontime="+82" swimtime="00:01:12.62" resultid="5616" heatid="7553" lane="1" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="5617" heatid="7602" lane="4" entrytime="00:01:25.00" entrycourse="SCM" />
                <RESULT eventid="1470" points="321" swimtime="00:01:11.46" resultid="5618" heatid="7670" lane="2" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="5619" heatid="7771" lane="2" entrytime="00:02:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="365" reactiontime="+64" swimtime="00:02:08.41" resultid="5625" heatid="7931" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="150" swimtime="00:01:40.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5614" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="3093" number="2" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3071" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3115" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="358" swimtime="00:01:53.73" resultid="5626" heatid="7714" lane="5" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                    <SPLIT distance="100" swimtime="00:00:56.92" />
                    <SPLIT distance="150" swimtime="00:01:26.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5614" number="1" />
                    <RELAYPOSITION athleteid="3093" number="2" />
                    <RELAYPOSITION athleteid="3071" number="3" />
                    <RELAYPOSITION athleteid="3115" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1521" points="239" reactiontime="+84" swimtime="00:02:30.10" resultid="5621" heatid="7707" lane="2" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:18.52" />
                    <SPLIT distance="150" swimtime="00:01:57.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3080" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3109" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3100" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3087" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1370" points="204" reactiontime="+68" swimtime="00:02:54.36" resultid="5622" heatid="7572" lane="2" entrytime="00:02:43.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.45" />
                    <SPLIT distance="100" swimtime="00:01:36.26" />
                    <SPLIT distance="150" swimtime="00:02:22.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3080" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3109" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3100" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3087" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1679" points="246" reactiontime="+71" swimtime="00:02:26.44" resultid="5623" heatid="7817" lane="1" entrytime="00:02:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                    <SPLIT distance="100" swimtime="00:01:29.41" />
                    <SPLIT distance="150" swimtime="00:01:58.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3087" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3100" number="2" reactiontime="+92" />
                    <RELAYPOSITION athleteid="3071" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3115" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1126" points="207" reactiontime="+86" swimtime="00:02:16.49" resultid="5624" heatid="7409" lane="4" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:07.24" />
                    <SPLIT distance="150" swimtime="00:01:48.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3093" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="3109" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="3080" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3115" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AZS PWSZ R" name="AZS PWSZ Racibórz" nation="POL" region="SLA">
          <CONTACT city="Racibórz" email="m,kunicki@" name="Marcin Kunicki" phone="504 233 267" state="ŚLĄSK" street="Słowackiego 55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-04-11" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="3131">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="3132" heatid="7360" lane="5" entrytime="00:00:31.24" entrycourse="SCM" />
                <RESULT eventid="1109" points="227" reactiontime="+91" swimtime="00:03:00.33" resultid="3133" heatid="7397" lane="6" entrytime="00:03:01.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:23.15" />
                    <SPLIT distance="150" swimtime="00:02:17.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="226" reactiontime="+100" swimtime="00:03:17.95" resultid="3134" heatid="7477" lane="1" entrytime="00:03:15.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                    <SPLIT distance="100" swimtime="00:01:37.73" />
                    <SPLIT distance="150" swimtime="00:02:28.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="201" reactiontime="+93" swimtime="00:03:06.13" resultid="3135" heatid="7568" lane="1" entrytime="00:03:10.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                    <SPLIT distance="100" swimtime="00:01:27.61" />
                    <SPLIT distance="150" swimtime="00:02:16.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="239" reactiontime="+74" swimtime="00:01:29.52" resultid="3136" heatid="7601" lane="4" entrytime="00:01:27.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="218" swimtime="00:06:31.14" resultid="3137" heatid="7978" lane="5" entrytime="00:06:26.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.53" />
                    <SPLIT distance="100" swimtime="00:01:38.88" />
                    <SPLIT distance="150" swimtime="00:02:28.86" />
                    <SPLIT distance="200" swimtime="00:03:18.78" />
                    <SPLIT distance="250" swimtime="00:04:12.76" />
                    <SPLIT distance="300" swimtime="00:05:06.63" />
                    <SPLIT distance="350" swimtime="00:05:49.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="197" reactiontime="+92" swimtime="00:01:23.26" resultid="3138" heatid="7742" lane="6" entrytime="00:01:24.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="267" reactiontime="+89" swimtime="00:00:39.17" resultid="3139" heatid="7802" lane="2" entrytime="00:00:37.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Sebastian " gender="M" lastname="Filuś" nation="POL" athleteid="6475">
              <RESULTS>
                <RESULT eventid="1075" points="529" reactiontime="+83" swimtime="00:00:25.09" resultid="6476" heatid="7379" lane="6" entrytime="00:00:25.50" />
                <RESULT comment="M-9 - Niejednoczesne dotkniecie ściany w czasie wykonywania nawrotu" eventid="1109" reactiontime="+89" status="DSQ" swimtime="00:02:25.51" resultid="6477" heatid="7406" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:05.19" />
                    <SPLIT distance="150" swimtime="00:01:51.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="6478" heatid="7459" lane="4" entrytime="00:00:28.40" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="6479" heatid="7524" lane="4" entrytime="00:00:55.00" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="6480" heatid="7674" lane="6" entrytime="00:01:02.00" />
                <RESULT eventid="1628" reactiontime="+73" status="DNS" swimtime="00:00:00.00" resultid="6482" heatid="7774" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:01:04.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Patryk " gender="M" lastname="Suchodolski" nation="POL" athleteid="6483">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="6484" heatid="7379" lane="1" entrytime="00:00:25.50" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="6485" heatid="7406" lane="2" entrytime="00:02:19.00" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="6486" heatid="7485" lane="6" entrytime="00:02:30.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="6487" heatid="7611" lane="1" entrytime="00:01:06.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="6488" heatid="7560" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="6489" heatid="7646" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="6490" heatid="7813" lane="4" entrytime="00:00:29.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="JOKRA" name="KS Masters Jordan Kraków" nation="POL" region="MAL">
          <CONTACT name="mr" />
          <ATHLETES>
            <ATHLETE birthdate="1978-06-10" firstname="Grzegorz" gender="M" lastname="Dadej" nation="POL" license="500106200001" athleteid="3141">
              <RESULTS>
                <RESULT eventid="1200" points="390" reactiontime="+56" swimtime="00:00:30.93" resultid="3142" heatid="7456" lane="3" entrytime="00:00:30.59" />
                <RESULT eventid="1302" points="412" reactiontime="+81" swimtime="00:01:08.18" resultid="3143" heatid="7554" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="402" reactiontime="+63" swimtime="00:01:06.28" resultid="3144" heatid="7672" lane="1" entrytime="00:01:07.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="366" reactiontime="+55" swimtime="00:02:28.24" resultid="3145" heatid="7772" lane="2" entrytime="00:02:30.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:52.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="019/11" name="RMKS Rybnik" nation="POL" region="SLA">
          <CONTACT city="Rybnik" email="aniaduda0511@tlen.pl" name="Duda" phone="792666159" state="SLASK" street="Anna" zip="44-217" />
          <ATHLETES>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="3147">
              <RESULTS>
                <RESULT eventid="1058" points="510" reactiontime="+83" swimtime="00:00:29.09" resultid="3148" heatid="7343" lane="3" entrytime="00:00:28.80" />
                <RESULT eventid="1092" points="428" reactiontime="+93" swimtime="00:02:45.29" resultid="3149" heatid="7388" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:17.28" />
                    <SPLIT distance="150" swimtime="00:02:06.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="497" reactiontime="+85" swimtime="00:01:04.38" resultid="3150" heatid="7497" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="448" reactiontime="+85" swimtime="00:01:15.42" resultid="3151" heatid="7536" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="502" reactiontime="+80" swimtime="00:00:30.67" resultid="3152" heatid="7621" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1487" points="409" reactiontime="+84" swimtime="00:02:29.67" resultid="3153" heatid="7684" lane="6" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:51.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="426" reactiontime="+89" swimtime="00:01:13.15" resultid="3154" heatid="7735" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DELOD" name="DELFIN MASTERS Łódź" nation="POL" region="LOD">
          <CONTACT city="Łódź" email="jblasiak@biol.uni.lodz.pl" internet="http://www.delfinmasters.pl/" name="Błasiak" phone="696 033 013" state="ŁÓDZK" street="Podchorążych 35A m 20" zip="90-234" />
          <ATHLETES>
            <ATHLETE birthdate="1974-04-10" firstname="Grzegorz" gender="M" lastname="Rogalski" nation="POL" athleteid="3156">
              <RESULTS>
                <RESULT eventid="1075" points="398" reactiontime="+88" swimtime="00:00:27.58" resultid="3157" heatid="7371" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1504" points="389" reactiontime="+88" swimtime="00:02:16.11" resultid="3158" heatid="7697" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:04.72" />
                    <SPLIT distance="150" swimtime="00:01:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="361" swimtime="00:01:08.04" resultid="3159" heatid="7745" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-26" firstname="Ewa" gender="F" lastname="Cieplucha" nation="POL" athleteid="3160">
              <RESULTS>
                <RESULT eventid="1183" points="347" reactiontime="+68" swimtime="00:00:36.55" resultid="3161" heatid="7439" lane="4" entrytime="00:00:36.03" />
                <RESULT eventid="1453" points="324" reactiontime="+73" swimtime="00:01:20.38" resultid="3162" heatid="7656" lane="4" entrytime="00:01:18.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" athleteid="3163">
              <RESULTS>
                <RESULT eventid="1109" points="75" reactiontime="+107" swimtime="00:04:20.20" resultid="3164" heatid="7392" lane="1" entrytime="00:04:28.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.47" />
                    <SPLIT distance="100" swimtime="00:02:03.36" />
                    <SPLIT distance="150" swimtime="00:03:23.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="118" reactiontime="+104" swimtime="00:01:31.50" resultid="3165" heatid="7499" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="90" reactiontime="+106" swimtime="00:01:52.93" resultid="3166" heatid="7540" lane="6" entrytime="00:01:54.00" />
                <RESULT eventid="1436" points="64" reactiontime="+89" swimtime="00:00:54.24" resultid="3167" heatid="7624" lane="4" entrytime="00:00:54.51" />
                <RESULT eventid="1470" points="62" reactiontime="+104" swimtime="00:02:03.03" resultid="3168" heatid="7661" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="47" swimtime="00:02:14.01" resultid="3169" heatid="7736" lane="5" entrytime="00:02:04.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="94" reactiontime="+96" swimtime="00:00:55.44" resultid="3170" heatid="7789" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-11" firstname="Rafał" gender="M" lastname="Maciejewski" nation="POL" athleteid="3171">
              <RESULTS>
                <RESULT eventid="1075" points="255" reactiontime="+94" swimtime="00:00:32.01" resultid="3172" heatid="7362" lane="2" entrytime="00:00:30.01" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="3173" heatid="7450" lane="2" entrytime="00:00:35.09" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="3174" heatid="7509" lane="1" entrytime="00:01:10.12" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="3175" heatid="7665" lane="4" entrytime="00:01:20.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-11" firstname="Arkadiusz" gender="M" lastname="Piecyk" nation="POL" athleteid="3176">
              <RESULTS>
                <RESULT eventid="1075" points="337" reactiontime="+90" swimtime="00:00:29.16" resultid="3177" heatid="7354" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1200" points="285" reactiontime="+79" swimtime="00:00:34.33" resultid="3178" heatid="7448" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1470" points="307" reactiontime="+69" swimtime="00:01:12.51" resultid="3179" heatid="7664" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-18" firstname="Adam" gender="M" lastname="Jerzykowski" nation="POL" athleteid="3180">
              <RESULTS>
                <RESULT comment="Przekroczono limit czasu" eventid="1165" reactiontime="+126" status="DSQ" swimtime="00:00:00.00" resultid="3181" heatid="7914" lane="6" entrytime="00:21:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                    <SPLIT distance="150" swimtime="00:01:59.70" />
                    <SPLIT distance="200" swimtime="00:02:43.15" />
                    <SPLIT distance="250" swimtime="00:03:28.88" />
                    <SPLIT distance="300" swimtime="00:04:14.74" />
                    <SPLIT distance="350" swimtime="00:05:02.10" />
                    <SPLIT distance="400" swimtime="00:05:49.23" />
                    <SPLIT distance="450" swimtime="00:06:36.39" />
                    <SPLIT distance="500" swimtime="00:07:24.23" />
                    <SPLIT distance="550" swimtime="00:08:15.46" />
                    <SPLIT distance="600" swimtime="00:09:02.42" />
                    <SPLIT distance="650" swimtime="00:09:50.14" />
                    <SPLIT distance="700" swimtime="00:10:38.09" />
                    <SPLIT distance="750" swimtime="00:11:26.06" />
                    <SPLIT distance="800" swimtime="00:12:14.46" />
                    <SPLIT distance="850" swimtime="00:13:04.05" />
                    <SPLIT distance="900" swimtime="00:13:53.28" />
                    <SPLIT distance="950" swimtime="00:14:42.46" />
                    <SPLIT distance="1000" swimtime="00:15:31.35" />
                    <SPLIT distance="1050" swimtime="00:16:20.74" />
                    <SPLIT distance="1100" swimtime="00:17:08.98" />
                    <SPLIT distance="1150" swimtime="00:17:57.24" />
                    <SPLIT distance="1200" swimtime="00:18:45.30" />
                    <SPLIT distance="1250" swimtime="00:19:39.26" />
                    <SPLIT distance="1300" swimtime="00:20:31.37" />
                    <SPLIT distance="1350" swimtime="00:21:19.59" />
                    <SPLIT distance="1400" swimtime="00:22:08.00" />
                    <SPLIT distance="1450" swimtime="00:23:11.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="126" reactiontime="+74" swimtime="00:00:43.37" resultid="3182" heatid="7622" lane="3" />
                <RESULT eventid="1504" points="230" reactiontime="+81" swimtime="00:02:42.03" resultid="3183" heatid="7687" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:01:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="221" reactiontime="+85" swimtime="00:05:51.66" resultid="3184" heatid="8043" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:01:22.77" />
                    <SPLIT distance="150" swimtime="00:02:06.66" />
                    <SPLIT distance="200" swimtime="00:02:51.98" />
                    <SPLIT distance="250" swimtime="00:04:24.01" />
                    <SPLIT distance="300" swimtime="00:05:09.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-24" firstname="Piotr" gender="M" lastname="Gaede" nation="POL" athleteid="3185">
              <RESULTS>
                <RESULT eventid="1402" points="292" reactiontime="+91" swimtime="00:01:23.75" resultid="3186" heatid="7604" lane="1" entrytime="00:01:23.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="270" reactiontime="+96" swimtime="00:00:39.04" resultid="3187" heatid="7802" lane="4" entrytime="00:00:37.58" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-03" firstname="Tomasz" gender="M" lastname="Wiaderny" nation="POL" athleteid="3188">
              <RESULTS>
                <RESULT eventid="1075" points="231" reactiontime="+89" swimtime="00:00:33.07" resultid="3189" heatid="7359" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1200" points="157" reactiontime="+68" swimtime="00:00:41.85" resultid="3190" heatid="7448" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1268" points="205" reactiontime="+94" swimtime="00:01:16.19" resultid="3191" heatid="7506" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="182" reactiontime="+102" swimtime="00:00:38.43" resultid="3192" heatid="7628" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1504" points="160" swimtime="00:03:02.81" resultid="3193" heatid="7691" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:23.86" />
                    <SPLIT distance="150" swimtime="00:02:13.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="3194" heatid="7740" lane="4" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="299" reactiontime="+68" swimtime="00:02:17.27" resultid="3196" heatid="7929" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:13.07" />
                    <SPLIT distance="150" swimtime="00:01:43.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3176" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3185" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3156" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3188" number="4" reactiontime="+99" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3195" heatid="7710" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3176" number="1" />
                    <RELAYPOSITION athleteid="3180" number="2" />
                    <RELAYPOSITION athleteid="3188" number="3" />
                    <RELAYPOSITION athleteid="3156" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Masters Gorzów Wlkp." nation="POL" region="LBS">
          <CONTACT city="Osiedle Poznańskie" email="stanislaw.kaczmarek@tpv-tech.com" name="Kaczmarek Stanisław" phone="600277732" state="LUBUS" street="Liliowa 9" zip="66-446" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" license="79012614295" athleteid="3205">
              <RESULTS>
                <RESULT eventid="1109" points="459" reactiontime="+79" swimtime="00:02:22.68" resultid="3206" heatid="7406" lane="3" entrytime="00:02:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:08.63" />
                    <SPLIT distance="150" swimtime="00:01:49.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1165" points="511" swimtime="00:17:42.64" resultid="3207" heatid="7917" lane="5" entrytime="00:17:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:07.67" />
                    <SPLIT distance="150" swimtime="00:01:42.97" />
                    <SPLIT distance="200" swimtime="00:02:18.64" />
                    <SPLIT distance="250" swimtime="00:02:54.63" />
                    <SPLIT distance="300" swimtime="00:03:30.52" />
                    <SPLIT distance="350" swimtime="00:04:06.13" />
                    <SPLIT distance="400" swimtime="00:04:41.82" />
                    <SPLIT distance="450" swimtime="00:05:17.76" />
                    <SPLIT distance="500" swimtime="00:05:53.54" />
                    <SPLIT distance="550" swimtime="00:06:28.77" />
                    <SPLIT distance="600" swimtime="00:07:04.42" />
                    <SPLIT distance="650" swimtime="00:07:39.90" />
                    <SPLIT distance="700" swimtime="00:08:15.33" />
                    <SPLIT distance="750" swimtime="00:08:50.69" />
                    <SPLIT distance="800" swimtime="00:09:26.48" />
                    <SPLIT distance="850" swimtime="00:10:02.27" />
                    <SPLIT distance="900" swimtime="00:10:37.82" />
                    <SPLIT distance="950" swimtime="00:11:13.32" />
                    <SPLIT distance="1000" swimtime="00:11:49.11" />
                    <SPLIT distance="1050" swimtime="00:12:24.65" />
                    <SPLIT distance="1100" swimtime="00:13:00.02" />
                    <SPLIT distance="1150" swimtime="00:13:35.50" />
                    <SPLIT distance="1200" swimtime="00:14:11.31" />
                    <SPLIT distance="1250" swimtime="00:14:47.00" />
                    <SPLIT distance="1300" swimtime="00:15:22.52" />
                    <SPLIT distance="1350" swimtime="00:15:57.86" />
                    <SPLIT distance="1400" swimtime="00:16:33.48" />
                    <SPLIT distance="1450" swimtime="00:17:08.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="421" swimtime="00:02:40.92" resultid="3208" heatid="7484" lane="5" entrytime="00:02:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:17.23" />
                    <SPLIT distance="150" swimtime="00:01:59.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="441" reactiontime="+82" swimtime="00:02:23.30" resultid="3209" heatid="7571" lane="4" entrytime="00:02:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="100" swimtime="00:01:06.82" />
                    <SPLIT distance="150" swimtime="00:01:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="480" reactiontime="+80" swimtime="00:02:06.84" resultid="3210" heatid="7706" lane="6" entrytime="00:02:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="100" swimtime="00:01:01.72" />
                    <SPLIT distance="150" swimtime="00:01:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="432" reactiontime="+84" swimtime="00:05:11.48" resultid="3211" heatid="7983" lane="1" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:07.63" />
                    <SPLIT distance="150" swimtime="00:01:51.25" />
                    <SPLIT distance="200" swimtime="00:02:32.67" />
                    <SPLIT distance="250" swimtime="00:03:16.98" />
                    <SPLIT distance="300" swimtime="00:04:01.39" />
                    <SPLIT distance="350" swimtime="00:04:37.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="425" reactiontime="+75" swimtime="00:01:04.44" resultid="3212" heatid="7750" lane="4" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="496" reactiontime="+79" swimtime="00:04:28.70" resultid="3213" heatid="8058" lane="1" entrytime="00:04:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:04.09" />
                    <SPLIT distance="150" swimtime="00:01:37.92" />
                    <SPLIT distance="200" swimtime="00:02:12.22" />
                    <SPLIT distance="250" swimtime="00:02:46.56" />
                    <SPLIT distance="300" swimtime="00:03:20.54" />
                    <SPLIT distance="350" swimtime="00:03:55.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" license="55071506113" athleteid="5251">
              <RESULTS>
                <RESULT eventid="1075" points="137" reactiontime="+112" swimtime="00:00:39.36" resultid="5252" heatid="7350" lane="3" entrytime="00:00:38.20" entrycourse="SCM" />
                <RESULT eventid="1165" points="139" reactiontime="+123" swimtime="00:27:18.13" resultid="5253" heatid="7908" lane="4" entrytime="00:28:30.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.41" />
                    <SPLIT distance="100" swimtime="00:01:37.88" />
                    <SPLIT distance="150" swimtime="00:02:30.46" />
                    <SPLIT distance="200" swimtime="00:03:24.80" />
                    <SPLIT distance="250" swimtime="00:04:18.39" />
                    <SPLIT distance="300" swimtime="00:05:13.49" />
                    <SPLIT distance="350" swimtime="00:06:08.73" />
                    <SPLIT distance="400" swimtime="00:07:04.65" />
                    <SPLIT distance="450" swimtime="00:07:59.64" />
                    <SPLIT distance="500" swimtime="00:08:53.93" />
                    <SPLIT distance="550" swimtime="00:09:48.49" />
                    <SPLIT distance="600" swimtime="00:10:43.41" />
                    <SPLIT distance="650" swimtime="00:11:38.54" />
                    <SPLIT distance="700" swimtime="00:12:34.05" />
                    <SPLIT distance="750" swimtime="00:13:29.58" />
                    <SPLIT distance="800" swimtime="00:14:25.57" />
                    <SPLIT distance="850" swimtime="00:15:21.86" />
                    <SPLIT distance="900" swimtime="00:16:17.85" />
                    <SPLIT distance="950" swimtime="00:17:13.41" />
                    <SPLIT distance="1000" swimtime="00:18:08.88" />
                    <SPLIT distance="1050" swimtime="00:19:04.68" />
                    <SPLIT distance="1100" swimtime="00:19:59.37" />
                    <SPLIT distance="1150" swimtime="00:20:54.20" />
                    <SPLIT distance="1200" swimtime="00:21:49.61" />
                    <SPLIT distance="1250" swimtime="00:22:44.83" />
                    <SPLIT distance="1300" swimtime="00:23:39.39" />
                    <SPLIT distance="1350" swimtime="00:24:34.59" />
                    <SPLIT distance="1400" swimtime="00:25:29.49" />
                    <SPLIT distance="1450" swimtime="00:26:24.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G-3 - Wynurzenie głowy spod lustra wody po starcie poza 15m" eventid="1200" reactiontime="+80" status="DSQ" swimtime="00:00:54.81" resultid="5254" heatid="7444" lane="2" entrytime="00:00:51.90" entrycourse="SCM" />
                <RESULT eventid="1268" points="117" swimtime="00:01:31.66" resultid="5255" heatid="7504" lane="5" entrytime="00:01:24.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="122" reactiontime="+123" swimtime="00:01:51.86" resultid="5256" heatid="7595" lane="2" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="121" reactiontime="+115" swimtime="00:03:20.83" resultid="5257" heatid="7690" lane="6" entrytime="00:03:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                    <SPLIT distance="100" swimtime="00:01:35.58" />
                    <SPLIT distance="150" swimtime="00:02:29.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="129" reactiontime="+124" swimtime="00:00:49.95" resultid="5258" heatid="7791" lane="6" entrytime="00:00:55.00" entrycourse="SCM" />
                <RESULT eventid="1710" points="134" reactiontime="+123" swimtime="00:06:54.91" resultid="5259" heatid="8046" lane="1" entrytime="00:07:05.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:01:31.72" />
                    <SPLIT distance="150" swimtime="00:02:25.31" />
                    <SPLIT distance="200" swimtime="00:03:19.34" />
                    <SPLIT distance="250" swimtime="00:04:13.52" />
                    <SPLIT distance="300" swimtime="00:05:08.25" />
                    <SPLIT distance="350" swimtime="00:06:02.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="TJ Alcedo Vsetín" nation="CZE">
          <ATHLETES>
            <ATHLETE birthdate="1967-01-01" firstname="Pavel" gender="M" lastname="OBR " nation="POL" athleteid="3215">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="3216" heatid="7375" lane="6" entrytime="00:00:26.80" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="3217" heatid="7403" lane="4" entrytime="00:02:33.00" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="3218" heatid="7521" lane="1" entrytime="00:00:59.50" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="3219" heatid="7555" lane="5" entrytime="00:01:08.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="3220" heatid="7607" lane="5" entrytime="00:01:17.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DOL" name="10 Brygada Kawalerii Pancernej Świętoszów" nation="POL" region="DOL" shortname="10 Brygada Kawalerii Pancernej">
          <CONTACT city="Świdnica" email="horbacz.marcin@wp.pl" name="Horbacz Marcin" phone="603672717" state="LUB" street="Buchałów 12c" zip="66-008" />
          <ATHLETES>
            <ATHLETE birthdate="1974-12-15" firstname="Oskar" gender="M" lastname="Bogucki" nation="POL" athleteid="3223">
              <RESULTS>
                <RESULT eventid="1075" points="273" reactiontime="+84" swimtime="00:00:31.26" resultid="3224" heatid="7360" lane="2" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1234" points="236" reactiontime="+90" swimtime="00:03:15.20" resultid="3225" heatid="7477" lane="3" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                    <SPLIT distance="100" swimtime="00:01:32.26" />
                    <SPLIT distance="150" swimtime="00:02:24.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="286" reactiontime="+86" swimtime="00:01:24.36" resultid="3226" heatid="7603" lane="1" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="309" swimtime="00:00:37.31" resultid="3227" heatid="7801" lane="5" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-14" firstname="Jarosław" gender="M" lastname="Druciarek" nation="POL" athleteid="3228">
              <RESULTS>
                <RESULT eventid="1075" points="322" reactiontime="+75" swimtime="00:00:29.60" resultid="3229" heatid="7371" lane="1" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1268" points="288" reactiontime="+88" swimtime="00:01:08.01" resultid="3230" heatid="7515" lane="1" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="3231" heatid="7627" lane="3" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1504" points="238" reactiontime="+95" swimtime="00:02:40.31" resultid="3232" heatid="7697" lane="2" entrytime="00:02:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="150" swimtime="00:02:00.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="202" reactiontime="+93" swimtime="00:06:02.16" resultid="3233" heatid="8049" lane="6" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:22.59" />
                    <SPLIT distance="150" swimtime="00:02:09.28" />
                    <SPLIT distance="200" swimtime="00:02:56.73" />
                    <SPLIT distance="250" swimtime="00:03:44.70" />
                    <SPLIT distance="300" swimtime="00:04:33.14" />
                    <SPLIT distance="350" swimtime="00:05:19.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-16" firstname="Marcin" gender="M" lastname="Horbacz" nation="POL" athleteid="3234">
              <RESULTS>
                <RESULT eventid="1075" points="427" reactiontime="+86" swimtime="00:00:26.95" resultid="3235" heatid="7374" lane="6" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1234" points="415" reactiontime="+86" swimtime="00:02:41.66" resultid="3236" heatid="7473" lane="6" entrytime="00:04:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:16.44" />
                    <SPLIT distance="150" swimtime="00:01:58.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="3237" heatid="7556" lane="3" entrytime="00:01:07.00" entrycourse="SCM" />
                <RESULT eventid="1504" points="492" reactiontime="+87" swimtime="00:02:05.79" resultid="3238" heatid="7705" lane="1" entrytime="00:02:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                    <SPLIT distance="100" swimtime="00:01:01.59" />
                    <SPLIT distance="150" swimtime="00:01:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="427" reactiontime="+73" swimtime="00:00:33.52" resultid="3239" heatid="7809" lane="1" entrytime="00:00:34.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-11-04" firstname="Mariusz" gender="M" lastname="Janowski" nation="POL" athleteid="3240">
              <RESULTS>
                <RESULT eventid="1075" points="317" reactiontime="+88" swimtime="00:00:29.76" resultid="3241" heatid="7360" lane="4" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1234" points="236" reactiontime="+94" swimtime="00:03:15.05" resultid="3242" heatid="7478" lane="6" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:01:31.25" />
                    <SPLIT distance="150" swimtime="00:02:22.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="263" reactiontime="+95" swimtime="00:01:26.71" resultid="3243" heatid="7603" lane="4" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="291" reactiontime="+89" swimtime="00:00:38.07" resultid="3244" heatid="7801" lane="6" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-29" firstname="Radosław" gender="M" lastname="Stępień" nation="POL" athleteid="3245">
              <RESULTS>
                <RESULT eventid="1075" points="360" reactiontime="+77" swimtime="00:00:28.51" resultid="3246" heatid="7370" lane="1" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1268" points="304" reactiontime="+79" swimtime="00:01:06.79" resultid="3247" heatid="7514" lane="3" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="232" swimtime="00:01:30.45" resultid="3248" heatid="7600" lane="5" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="250" reactiontime="+80" swimtime="00:00:40.05" resultid="3249" heatid="7800" lane="6" entrytime="00:00:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-27" firstname="Natalia" gender="F" lastname="Szczęsnowicz" nation="POL" athleteid="3250">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="3251" heatid="7341" lane="3" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1251" points="302" reactiontime="+72" swimtime="00:01:16.02" resultid="3252" heatid="7492" lane="4" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="329" reactiontime="+69" swimtime="00:00:35.30" resultid="3253" heatid="7618" lane="2" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="310" reactiontime="+63" swimtime="00:02:15.52" resultid="3254" heatid="7929" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:02:15.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3234" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="3223" number="2" />
                    <RELAYPOSITION athleteid="3228" number="3" />
                    <RELAYPOSITION athleteid="3245" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1528" points="347" reactiontime="+78" swimtime="00:01:54.85" resultid="3255" heatid="7715" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="100" swimtime="00:00:56.66" />
                    <SPLIT distance="150" swimtime="00:01:26.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3234" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3228" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3240" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3245" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="07614" name="UKS Gos Raszyn" nation="POL" region="14">
          <ATHLETES>
            <ATHLETE birthdate="1968-01-01" firstname="Tomasz" gender="M" lastname="Rozmysłowski" nation="POL" athleteid="3259">
              <RESULTS>
                <RESULT eventid="1075" points="407" reactiontime="+77" swimtime="00:00:27.38" resultid="3260" heatid="7377" lane="1" entrytime="00:00:26.39" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Msc &quot;Euro-Lviv&quot;" nation="UKR">
          <CONTACT city="Lviv" email="riff@mail.lviv.ua" fax="+380322430304" name="Ruslan Friauf" phone="+380676734796" street="Karpincya 18A/3" zip="79012" />
          <ATHLETES>
            <ATHLETE birthdate="1976-02-23" firstname="Oleksandr" gender="M" lastname="Shavrov" nation="UKR" athleteid="5299">
              <RESULTS>
                <RESULT eventid="1234" points="361" reactiontime="+79" swimtime="00:02:49.35" resultid="5300" heatid="7480" lane="6" entrytime="00:03:00.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                    <SPLIT distance="100" swimtime="00:01:20.54" />
                    <SPLIT distance="150" swimtime="00:02:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="398" swimtime="00:01:15.55" resultid="5301" heatid="7606" lane="5" entrytime="00:01:20.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="400" reactiontime="+80" swimtime="00:00:34.25" resultid="5302" heatid="7806" lane="2" entrytime="00:00:35.09" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-08" firstname="Ihor" gender="M" lastname="Rudnyk" nation="UKR" athleteid="5303">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5304" heatid="7355" lane="1" entrytime="00:00:33.60" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="5305" heatid="7795" lane="6" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-06-05" firstname="Mykhailo" gender="M" lastname="Shelest" nation="UKR" athleteid="5306">
              <RESULTS>
                <RESULT eventid="1200" points="211" reactiontime="+76" swimtime="00:00:37.93" resultid="5307" heatid="7448" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1302" points="243" reactiontime="+93" swimtime="00:01:21.29" resultid="5308" heatid="7546" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="256" swimtime="00:01:27.55" resultid="5309" heatid="7602" lane="5" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="5310" heatid="7664" lane="4" entrytime="00:01:25.00" />
                <RESULT eventid="1662" points="279" reactiontime="+103" swimtime="00:00:38.62" resultid="5311" heatid="7801" lane="1" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-22" firstname="Volodymyr" gender="M" lastname="Rybko" nation="UKR" athleteid="5312">
              <RESULTS>
                <RESULT eventid="1109" points="303" reactiontime="+94" swimtime="00:02:43.77" resultid="5313" heatid="7405" lane="3" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:15.25" />
                    <SPLIT distance="150" swimtime="00:02:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="313" reactiontime="+94" swimtime="00:20:51.10" resultid="5314" heatid="7917" lane="2" entrytime="00:17:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:01:57.23" />
                    <SPLIT distance="200" swimtime="00:02:38.34" />
                    <SPLIT distance="250" swimtime="00:03:20.35" />
                    <SPLIT distance="300" swimtime="00:04:02.36" />
                    <SPLIT distance="350" swimtime="00:04:44.54" />
                    <SPLIT distance="400" swimtime="00:05:25.97" />
                    <SPLIT distance="450" swimtime="00:06:08.53" />
                    <SPLIT distance="500" swimtime="00:06:49.51" />
                    <SPLIT distance="550" swimtime="00:07:32.45" />
                    <SPLIT distance="600" swimtime="00:08:15.49" />
                    <SPLIT distance="650" swimtime="00:08:58.84" />
                    <SPLIT distance="700" swimtime="00:09:42.28" />
                    <SPLIT distance="750" swimtime="00:10:24.57" />
                    <SPLIT distance="800" swimtime="00:11:07.00" />
                    <SPLIT distance="850" swimtime="00:11:50.96" />
                    <SPLIT distance="900" swimtime="00:12:33.42" />
                    <SPLIT distance="950" swimtime="00:13:16.33" />
                    <SPLIT distance="1000" swimtime="00:13:59.61" />
                    <SPLIT distance="1050" swimtime="00:14:42.39" />
                    <SPLIT distance="1100" swimtime="00:15:25.82" />
                    <SPLIT distance="1150" swimtime="00:16:07.48" />
                    <SPLIT distance="1200" swimtime="00:16:48.94" />
                    <SPLIT distance="1250" swimtime="00:17:30.63" />
                    <SPLIT distance="1300" swimtime="00:18:12.68" />
                    <SPLIT distance="1350" swimtime="00:18:54.71" />
                    <SPLIT distance="1400" swimtime="00:19:35.73" />
                    <SPLIT distance="1450" swimtime="00:20:15.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="342" reactiontime="+83" swimtime="00:01:04.22" resultid="5315" heatid="7521" lane="3" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="349" reactiontime="+88" swimtime="00:01:12.09" resultid="5316" heatid="7554" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="370" reactiontime="+85" swimtime="00:00:30.34" resultid="5317" heatid="7646" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1559" points="267" reactiontime="+99" swimtime="00:06:05.39" resultid="5318" heatid="7983" lane="2" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:20.18" />
                    <SPLIT distance="150" swimtime="00:02:08.85" />
                    <SPLIT distance="200" swimtime="00:02:56.06" />
                    <SPLIT distance="250" swimtime="00:03:52.73" />
                    <SPLIT distance="300" swimtime="00:04:48.37" />
                    <SPLIT distance="350" swimtime="00:05:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="285" reactiontime="+86" swimtime="00:01:13.62" resultid="5319" heatid="7749" lane="6" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="292" reactiontime="+95" swimtime="00:05:20.36" resultid="5320" heatid="8043" lane="1" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="150" swimtime="00:01:59.14" />
                    <SPLIT distance="200" swimtime="00:02:40.88" />
                    <SPLIT distance="250" swimtime="00:03:23.43" />
                    <SPLIT distance="300" swimtime="00:04:03.82" />
                    <SPLIT distance="350" swimtime="00:04:43.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-05" firstname="Lyudmyla" gender="F" lastname="Khiresh" nation="UKR" athleteid="5321">
              <RESULTS>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1058" reactiontime="+67" status="DSQ" swimtime="00:00:35.48" resultid="5322" heatid="7338" lane="2" entrytime="00:00:35.50" />
                <RESULT eventid="1183" points="294" reactiontime="+73" swimtime="00:00:38.63" resultid="5323" heatid="7437" lane="4" entrytime="00:00:39.50" />
                <RESULT eventid="1285" points="305" reactiontime="+84" swimtime="00:01:25.76" resultid="5324" heatid="7530" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="273" reactiontime="+78" swimtime="00:01:25.08" resultid="5325" heatid="7653" lane="4" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-06-01" firstname="Serhiy" gender="M" lastname="Simankov" nation="UKR" athleteid="5326">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5327" heatid="7349" lane="2" entrytime="00:00:41.66" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="5328" heatid="7502" lane="1" entrytime="00:01:38.65" />
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="5329" heatid="7624" lane="3" entrytime="00:00:48.66" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5330" heatid="7737" lane="3" entrytime="00:02:09.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-10-31" firstname="Dmytro" gender="M" lastname="Ishchenko" nation="UKR" athleteid="5331">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5332" heatid="7365" lane="1" entrytime="00:00:29.80" />
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="5333" heatid="7634" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5334" heatid="7744" lane="1" entrytime="00:01:18.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-11-17" firstname="Iurii" gender="M" lastname="Viiuk" nation="UKR" athleteid="5335">
              <RESULTS>
                <RESULT eventid="1075" points="310" swimtime="00:00:29.98" resultid="5336" heatid="7364" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1402" points="287" reactiontime="+97" swimtime="00:01:24.24" resultid="5337" heatid="7602" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="320" swimtime="00:00:36.88" resultid="5338" heatid="7803" lane="5" entrytime="00:00:37.17" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-08-08" firstname="Andrii" gender="M" lastname="Hertsyk" nation="UKR" athleteid="5339">
              <RESULTS>
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="5340" heatid="7600" lane="1" entrytime="00:01:30.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="5341" heatid="7799" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-11" firstname="Natalya" gender="F" lastname="Hertsyk" nation="UKR" athleteid="5342">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="5343" heatid="7337" lane="2" entrytime="00:00:36.90" />
                <RESULT eventid="1419" status="DNS" swimtime="00:00:00.00" resultid="5344" heatid="7616" lane="6" entrytime="00:00:40.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-05-09" firstname="Lidiya" gender="F" lastname="Tymoshenko" nation="UKR" athleteid="5345">
              <RESULTS>
                <RESULT eventid="1058" points="131" reactiontime="+103" swimtime="00:00:45.75" resultid="5346" heatid="7333" lane="3" entrytime="00:00:49.60" />
                <RESULT eventid="1183" points="71" reactiontime="+77" swimtime="00:01:01.86" resultid="5347" heatid="7432" lane="4" entrytime="00:01:04.83" />
                <RESULT eventid="1251" points="90" reactiontime="+108" swimtime="00:01:53.80" resultid="5348" heatid="7487" lane="2" entrytime="00:01:55.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="119" reactiontime="+122" swimtime="00:02:07.44" resultid="5349" heatid="7583" lane="3" entrytime="00:02:09.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="133" reactiontime="+118" swimtime="00:00:56.34" resultid="5350" heatid="7777" lane="2" entrytime="00:00:58.76" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-11" firstname="Alla" gender="F" lastname="Poniavina" nation="UKR" athleteid="5351">
              <RESULTS>
                <RESULT eventid="1148" points="369" swimtime="00:11:14.97" resultid="5352" heatid="7905" lane="5" entrytime="00:11:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="150" swimtime="00:01:59.60" />
                    <SPLIT distance="200" swimtime="00:02:41.92" />
                    <SPLIT distance="250" swimtime="00:03:24.80" />
                    <SPLIT distance="300" swimtime="00:04:08.02" />
                    <SPLIT distance="350" swimtime="00:04:50.94" />
                    <SPLIT distance="400" swimtime="00:05:33.84" />
                    <SPLIT distance="450" swimtime="00:06:16.46" />
                    <SPLIT distance="500" swimtime="00:06:59.01" />
                    <SPLIT distance="550" swimtime="00:07:41.68" />
                    <SPLIT distance="600" swimtime="00:08:24.00" />
                    <SPLIT distance="650" swimtime="00:09:06.60" />
                    <SPLIT distance="700" swimtime="00:09:49.54" />
                    <SPLIT distance="750" swimtime="00:10:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="409" reactiontime="+90" swimtime="00:01:08.68" resultid="5353" heatid="7496" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="393" reactiontime="+88" swimtime="00:01:18.81" resultid="5354" heatid="7536" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="360" reactiontime="+75" swimtime="00:01:17.63" resultid="5355" heatid="7656" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="378" reactiontime="+86" swimtime="00:02:33.71" resultid="5356" heatid="7682" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:14.01" />
                    <SPLIT distance="150" swimtime="00:01:54.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="363" reactiontime="+78" swimtime="00:02:48.17" resultid="5357" heatid="7756" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:01:21.87" />
                    <SPLIT distance="150" swimtime="00:02:05.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="364" reactiontime="+92" swimtime="00:05:28.85" resultid="5358" heatid="8024" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:16.67" />
                    <SPLIT distance="150" swimtime="00:01:58.60" />
                    <SPLIT distance="200" swimtime="00:02:41.24" />
                    <SPLIT distance="250" swimtime="00:03:23.89" />
                    <SPLIT distance="300" swimtime="00:04:06.74" />
                    <SPLIT distance="350" swimtime="00:04:49.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-18" firstname="Vladyslav" gender="M" lastname="Horovoy" nation="UKR" athleteid="5359">
              <RESULTS>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="5360" heatid="7523" lane="3" entrytime="00:00:57.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="5361" heatid="7705" lane="5" entrytime="00:02:07.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-18" firstname="Igor" gender="M" lastname="Shchotkin" nation="UKR" athleteid="5368">
              <RESULTS>
                <RESULT eventid="1075" points="541" swimtime="00:00:24.91" resultid="5369" heatid="7379" lane="2" entrytime="00:00:24.50" />
                <RESULT eventid="1268" points="506" reactiontime="+76" swimtime="00:00:56.37" resultid="5370" heatid="7524" lane="1" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="517" reactiontime="+69" swimtime="00:00:27.16" resultid="5371" heatid="7646" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1662" points="518" reactiontime="+72" swimtime="00:00:31.42" resultid="5372" heatid="7812" lane="1" entrytime="00:00:31.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-03-29" firstname="Tetyana" gender="F" lastname="Zelikova" nation="UKR" athleteid="5373">
              <RESULTS>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5374" heatid="7782" lane="6" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-08-09" firstname="Igor" gender="M" lastname="Medvediev" nation="UKR" athleteid="5375">
              <RESULTS>
                <RESULT eventid="1234" points="453" reactiontime="+76" swimtime="00:02:37.08" resultid="5376" heatid="7483" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:16.31" />
                    <SPLIT distance="150" swimtime="00:01:56.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="476" reactiontime="+77" swimtime="00:01:11.21" resultid="5377" heatid="7610" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="371" reactiontime="+77" swimtime="00:00:30.32" resultid="5378" heatid="7643" lane="1" entrytime="00:00:28.50" />
                <RESULT eventid="1662" points="478" reactiontime="+78" swimtime="00:00:32.28" resultid="5379" heatid="7811" lane="2" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="Friauf" nation="UKR" athleteid="5380">
              <RESULTS>
                <RESULT eventid="1109" points="225" reactiontime="+83" swimtime="00:03:00.91" resultid="5381" heatid="7398" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="150" swimtime="00:02:16.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="232" reactiontime="+79" swimtime="00:00:36.78" resultid="5382" heatid="7449" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1302" points="274" reactiontime="+82" swimtime="00:01:18.13" resultid="5383" heatid="7546" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-03-11" firstname="Lyudmyla" gender="F" lastname="Maksymiv" nation="UKR" athleteid="5384">
              <RESULTS>
                <RESULT eventid="1217" points="210" reactiontime="+105" swimtime="00:03:46.16" resultid="5385" heatid="7465" lane="4" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.79" />
                    <SPLIT distance="100" swimtime="00:01:52.35" />
                    <SPLIT distance="150" swimtime="00:02:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="196" reactiontime="+104" swimtime="00:01:47.79" resultid="5386" heatid="7585" lane="4" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="161" reactiontime="+81" swimtime="00:01:41.37" resultid="5387" heatid="7650" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="190" swimtime="00:00:50.07" resultid="5388" heatid="7780" lane="5" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-08-05" firstname="Iryna" gender="F" lastname="Ponomarenko" nation="UKR" athleteid="5389">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="5390" heatid="7341" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="5391" heatid="7495" lane="2" entrytime="00:01:12.00" />
                <RESULT eventid="1487" status="DNS" swimtime="00:00:00.00" resultid="5392" heatid="7682" lane="1" entrytime="00:02:45.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5393" heatid="7784" lane="4" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1528" points="405" reactiontime="+69" swimtime="00:01:49.15" resultid="5396" heatid="7716" lane="6" entrytime="00:01:46.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.04" />
                    <SPLIT distance="100" swimtime="00:00:53.97" />
                    <SPLIT distance="150" swimtime="00:01:21.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5299" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="5312" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="5375" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="5368" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1377" status="DNS" swimtime="00:00:00.00" resultid="5397" heatid="7932" lane="2" entrytime="00:02:08.86">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5380" number="1" />
                    <RELAYPOSITION athleteid="5299" number="2" />
                    <RELAYPOSITION athleteid="5312" number="3" />
                    <RELAYPOSITION athleteid="5331" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1377" points="372" reactiontime="+78" swimtime="00:02:07.58" resultid="5399" heatid="7933" lane="3" entrytime="00:02:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:10.13" />
                    <SPLIT distance="150" swimtime="00:01:37.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5306" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="5375" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="5368" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="5335" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="5400" heatid="7712" lane="1" entrytime="00:02:05.30">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5335" number="1" />
                    <RELAYPOSITION athleteid="5331" number="2" />
                    <RELAYPOSITION athleteid="5380" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1521" status="DNS" swimtime="00:00:00.00" resultid="5401" heatid="7708" lane="6" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5389" number="1" />
                    <RELAYPOSITION athleteid="5321" number="2" />
                    <RELAYPOSITION athleteid="5384" number="3" />
                    <RELAYPOSITION athleteid="5351" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="5394" heatid="7819" lane="1" entrytime="00:02:09.20">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5321" number="1" />
                    <RELAYPOSITION athleteid="5368" number="2" />
                    <RELAYPOSITION athleteid="5312" number="3" />
                    <RELAYPOSITION athleteid="5351" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1126" points="310" reactiontime="+93" swimtime="00:01:59.26" resultid="5395" heatid="7411" lane="4" entrytime="00:01:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:00:58.65" />
                    <SPLIT distance="150" swimtime="00:01:34.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5351" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="5312" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="5389" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="5368" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1679" points="154" reactiontime="+83" swimtime="00:02:51.01" resultid="5398" heatid="7816" lane="6" entrytime="00:02:48.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:22.86" />
                    <SPLIT distance="150" swimtime="00:02:09.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5306" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="5373" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5335" number="3" reactiontime="+98" />
                    <RELAYPOSITION athleteid="5345" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Gdynia Masters" nation="POL">
          <CONTACT email="k.mysiak@wpit.am.gdynia.pl" name="Mysiak Katarzyna" />
          <ATHLETES>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="3367">
              <RESULTS>
                <RESULT eventid="1075" points="191" reactiontime="+99" swimtime="00:00:35.21" resultid="3368" heatid="7354" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1234" points="195" reactiontime="+94" swimtime="00:03:27.77" resultid="3369" heatid="7475" lane="2" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:38.18" />
                    <SPLIT distance="150" swimtime="00:02:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="231" swimtime="00:01:30.57" resultid="3370" heatid="7599" lane="5" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="230" reactiontime="+83" swimtime="00:00:41.16" resultid="3371" heatid="7796" lane="6" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="3372">
              <RESULTS>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="3373" heatid="7445" lane="2" entrytime="00:00:48.86" />
                <RESULT comment="Rekord Polski Masters" eventid="1234" points="129" reactiontime="+91" swimtime="00:03:58.81" resultid="3374" heatid="7472" lane="3" entrytime="00:04:11.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.51" />
                    <SPLIT distance="100" swimtime="00:01:53.74" />
                    <SPLIT distance="150" swimtime="00:02:56.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1402" points="135" reactiontime="+100" swimtime="00:01:48.30" resultid="3375" heatid="7595" lane="4" entrytime="00:01:48.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="138" reactiontime="+95" swimtime="00:00:48.77" resultid="3376" heatid="7792" lane="4" entrytime="00:00:48.76" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="Mikołajczyk" nation="POL" athleteid="3377">
              <RESULTS>
                <RESULT eventid="1109" points="109" reactiontime="+93" swimtime="00:03:50.43" resultid="3378" heatid="7394" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.80" />
                    <SPLIT distance="100" swimtime="00:01:55.63" />
                    <SPLIT distance="150" swimtime="00:02:56.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" status="WDR" swimtime="00:00:00.00" resultid="3379" entrytime="00:03:40.00" />
                <RESULT eventid="1336" status="DNS" swimtime="00:00:00.00" resultid="3380" heatid="7566" lane="4" entrytime="00:03:50.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="3381" heatid="7596" lane="4" entrytime="00:01:40.00" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="3383" heatid="7739" lane="2" entrytime="00:01:45.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="3384" heatid="7793" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Barbara" gender="F" lastname="Chomicka" nation="POL" athleteid="3385">
              <RESULTS>
                <RESULT eventid="1092" points="95" reactiontime="+107" swimtime="00:04:33.00" resultid="3386" heatid="7383" lane="3" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.72" />
                    <SPLIT distance="100" swimtime="00:02:13.91" />
                    <SPLIT distance="150" swimtime="00:03:25.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="103" reactiontime="+73" swimtime="00:00:54.73" resultid="3387" heatid="7432" lane="3" entrytime="00:00:55.00" />
                <RESULT eventid="1319" points="57" reactiontime="+112" swimtime="00:05:12.49" resultid="3388" heatid="7561" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.54" />
                    <SPLIT distance="100" swimtime="00:02:29.41" />
                    <SPLIT distance="150" swimtime="00:03:53.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" status="DNS" swimtime="00:00:00.00" resultid="3389" heatid="7613" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="1453" points="97" reactiontime="+76" swimtime="00:01:59.99" resultid="3390" heatid="7649" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="58" reactiontime="+115" swimtime="00:02:21.89" resultid="3391" heatid="7730" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="84" reactiontime="+79" swimtime="00:04:33.89" resultid="3392" heatid="7755" lane="5" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:14.82" />
                    <SPLIT distance="150" swimtime="00:03:26.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Leszek" gender="M" lastname="Kubicki" nation="POL" athleteid="3393">
              <RESULTS>
                <RESULT eventid="1075" points="249" reactiontime="+102" swimtime="00:00:32.24" resultid="3394" heatid="7356" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1165" points="227" reactiontime="+105" swimtime="00:23:13.34" resultid="3395" heatid="7912" lane="2" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                    <SPLIT distance="100" swimtime="00:01:18.94" />
                    <SPLIT distance="150" swimtime="00:02:04.25" />
                    <SPLIT distance="200" swimtime="00:02:50.25" />
                    <SPLIT distance="250" swimtime="00:03:36.59" />
                    <SPLIT distance="300" swimtime="00:04:22.96" />
                    <SPLIT distance="350" swimtime="00:05:09.22" />
                    <SPLIT distance="400" swimtime="00:05:56.09" />
                    <SPLIT distance="450" swimtime="00:06:43.13" />
                    <SPLIT distance="500" swimtime="00:07:29.97" />
                    <SPLIT distance="550" swimtime="00:08:17.34" />
                    <SPLIT distance="600" swimtime="00:09:04.00" />
                    <SPLIT distance="650" swimtime="00:09:50.96" />
                    <SPLIT distance="700" swimtime="00:10:38.22" />
                    <SPLIT distance="750" swimtime="00:11:24.95" />
                    <SPLIT distance="800" swimtime="00:12:12.12" />
                    <SPLIT distance="850" swimtime="00:12:59.14" />
                    <SPLIT distance="900" swimtime="00:13:46.44" />
                    <SPLIT distance="950" swimtime="00:14:33.46" />
                    <SPLIT distance="1000" swimtime="00:15:20.60" />
                    <SPLIT distance="1050" swimtime="00:16:08.17" />
                    <SPLIT distance="1100" swimtime="00:16:56.10" />
                    <SPLIT distance="1150" swimtime="00:17:43.04" />
                    <SPLIT distance="1200" swimtime="00:18:30.30" />
                    <SPLIT distance="1250" swimtime="00:19:17.82" />
                    <SPLIT distance="1300" swimtime="00:20:05.27" />
                    <SPLIT distance="1350" swimtime="00:20:53.18" />
                    <SPLIT distance="1400" swimtime="00:21:40.58" />
                    <SPLIT distance="1450" swimtime="00:22:27.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="229" reactiontime="+103" swimtime="00:01:13.41" resultid="3396" heatid="7507" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="196" reactiontime="+97" swimtime="00:01:27.36" resultid="3397" heatid="7544" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="3398" heatid="7596" lane="6" entrytime="00:01:45.00" />
                <RESULT eventid="1504" points="205" reactiontime="+102" swimtime="00:02:48.47" resultid="3399" heatid="7693" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:17.24" />
                    <SPLIT distance="150" swimtime="00:02:02.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="3400" heatid="7800" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1710" points="209" reactiontime="+105" swimtime="00:05:58.18" resultid="3401" heatid="8050" lane="6" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                    <SPLIT distance="150" swimtime="00:02:05.29" />
                    <SPLIT distance="200" swimtime="00:02:51.46" />
                    <SPLIT distance="250" swimtime="00:03:37.94" />
                    <SPLIT distance="300" swimtime="00:04:24.65" />
                    <SPLIT distance="350" swimtime="00:05:11.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Hanka" gender="F" lastname="Kania" nation="POL" athleteid="3402">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="3403" heatid="7336" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1092" points="172" swimtime="00:03:43.71" resultid="3404" heatid="7384" lane="5" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.84" />
                    <SPLIT distance="100" swimtime="00:01:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="192" reactiontime="+119" swimtime="00:03:53.08" resultid="3405" heatid="7464" lane="4" entrytime="00:04:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.27" />
                    <SPLIT distance="100" swimtime="00:01:51.14" />
                    <SPLIT distance="150" swimtime="00:02:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="189" reactiontime="+113" swimtime="00:01:40.61" resultid="3406" heatid="7528" lane="1" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="180" reactiontime="+109" swimtime="00:01:51.04" resultid="3407" heatid="7584" lane="3" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="133" reactiontime="+120" swimtime="00:00:47.66" resultid="3408" heatid="7614" lane="1" entrytime="00:00:49.00" />
                <RESULT eventid="1577" points="107" reactiontime="+122" swimtime="00:01:55.65" resultid="3409" heatid="7731" lane="3" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="188" reactiontime="+113" swimtime="00:00:50.20" resultid="3410" heatid="7779" lane="2" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="3411">
              <RESULTS>
                <RESULT eventid="1109" points="94" reactiontime="+112" swimtime="00:04:01.26" resultid="3412" heatid="7393" lane="4" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.46" />
                    <SPLIT distance="100" swimtime="00:02:00.47" />
                    <SPLIT distance="150" swimtime="00:03:06.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="97" reactiontime="+113" swimtime="00:04:22.43" resultid="3413" heatid="7473" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.77" />
                    <SPLIT distance="100" swimtime="00:02:04.84" />
                    <SPLIT distance="150" swimtime="00:03:15.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="102" reactiontime="+115" swimtime="00:01:48.35" resultid="3414" heatid="7541" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="117" reactiontime="+110" swimtime="00:01:53.54" resultid="3415" heatid="7596" lane="1" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="63" reactiontime="+107" swimtime="00:02:01.44" resultid="3416" heatid="7739" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="144" reactiontime="+110" swimtime="00:00:48.16" resultid="3417" heatid="7794" lane="2" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Katarzyna" gender="F" lastname="Gąsiorowska  " nation="POL" athleteid="4215">
              <RESULTS>
                <RESULT eventid="1058" points="488" reactiontime="+82" swimtime="00:00:29.52" resultid="4216" heatid="7343" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1148" points="392" reactiontime="+86" swimtime="00:11:01.50" resultid="4217" heatid="7905" lane="2" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:52.59" />
                    <SPLIT distance="200" swimtime="00:02:33.58" />
                    <SPLIT distance="250" swimtime="00:03:15.11" />
                    <SPLIT distance="300" swimtime="00:03:56.99" />
                    <SPLIT distance="350" swimtime="00:04:38.46" />
                    <SPLIT distance="400" swimtime="00:05:20.23" />
                    <SPLIT distance="450" swimtime="00:06:02.46" />
                    <SPLIT distance="500" swimtime="00:06:45.11" />
                    <SPLIT distance="550" swimtime="00:07:28.36" />
                    <SPLIT distance="600" swimtime="00:08:11.41" />
                    <SPLIT distance="650" swimtime="00:08:54.60" />
                    <SPLIT distance="700" swimtime="00:09:38.27" />
                    <SPLIT distance="750" swimtime="00:10:20.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="495" reactiontime="+82" swimtime="00:01:04.47" resultid="4218" heatid="7498" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="244" reactiontime="+88" swimtime="00:03:13.14" resultid="4219" heatid="7563" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:01:27.21" />
                    <SPLIT distance="150" swimtime="00:02:17.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="443" reactiontime="+84" swimtime="00:02:25.74" resultid="4220" heatid="7685" lane="1" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:48.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3420" heatid="7710" lane="3" entrytime="00:03:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3411" number="1" />
                    <RELAYPOSITION athleteid="3372" number="2" />
                    <RELAYPOSITION athleteid="3367" number="3" />
                    <RELAYPOSITION athleteid="3393" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="319" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" status="DNS" swimtime="00:00:00.00" resultid="3421" heatid="7929" lane="3" entrytime="00:03:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3411" number="1" />
                    <RELAYPOSITION athleteid="3372" number="2" />
                    <RELAYPOSITION athleteid="3377" number="3" />
                    <RELAYPOSITION athleteid="3393" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1679" points="344" reactiontime="+69" status="DNS" swimtime="00:02:10.89" resultid="3418" heatid="7816" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="150" swimtime="00:01:45.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3385" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3372" number="2" />
                    <RELAYPOSITION athleteid="3402" number="3" />
                    <RELAYPOSITION athleteid="3367" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="3419" heatid="7408" lane="3" entrytime="00:03:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3372" number="1" />
                    <RELAYPOSITION athleteid="3402" number="2" />
                    <RELAYPOSITION athleteid="3385" number="3" />
                    <RELAYPOSITION athleteid="3367" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AZS" name="AZS AWF Warszawa" nation="POL" region="14">
          <ATHLETES>
            <ATHLETE birthdate="1991-06-23" firstname="Sebastian" gender="M" lastname="Karaś" nation="POL" license="100114200067" athleteid="3428">
              <RESULTS>
                <RESULT eventid="1075" points="513" reactiontime="+73" swimtime="00:00:25.35" resultid="3429" heatid="7381" lane="6" entrytime="00:00:24.50" />
                <RESULT eventid="1165" points="695" reactiontime="+72" swimtime="00:15:59.47" resultid="3430" heatid="7917" lane="4" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="100" swimtime="00:01:01.52" />
                    <SPLIT distance="150" swimtime="00:01:33.72" />
                    <SPLIT distance="200" swimtime="00:02:05.65" />
                    <SPLIT distance="250" swimtime="00:02:37.55" />
                    <SPLIT distance="300" swimtime="00:03:09.46" />
                    <SPLIT distance="350" swimtime="00:03:41.30" />
                    <SPLIT distance="400" swimtime="00:04:13.12" />
                    <SPLIT distance="450" swimtime="00:04:44.96" />
                    <SPLIT distance="500" swimtime="00:05:16.98" />
                    <SPLIT distance="550" swimtime="00:05:48.91" />
                    <SPLIT distance="600" swimtime="00:06:21.08" />
                    <SPLIT distance="650" swimtime="00:06:53.37" />
                    <SPLIT distance="700" swimtime="00:07:25.42" />
                    <SPLIT distance="750" swimtime="00:07:57.50" />
                    <SPLIT distance="800" swimtime="00:08:29.50" />
                    <SPLIT distance="850" swimtime="00:09:01.76" />
                    <SPLIT distance="900" swimtime="00:09:33.94" />
                    <SPLIT distance="950" swimtime="00:10:06.25" />
                    <SPLIT distance="1000" swimtime="00:10:38.23" />
                    <SPLIT distance="1050" swimtime="00:11:10.75" />
                    <SPLIT distance="1100" swimtime="00:11:42.96" />
                    <SPLIT distance="1150" swimtime="00:12:15.06" />
                    <SPLIT distance="1200" swimtime="00:12:47.04" />
                    <SPLIT distance="1250" swimtime="00:13:19.10" />
                    <SPLIT distance="1300" swimtime="00:13:51.15" />
                    <SPLIT distance="1350" swimtime="00:14:23.13" />
                    <SPLIT distance="1400" swimtime="00:14:55.77" />
                    <SPLIT distance="1450" swimtime="00:15:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="570" reactiontime="+60" swimtime="00:00:27.26" resultid="3431" heatid="7460" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="3432" heatid="7560" lane="5" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06614" name="Legia Warszawa" nation="POL" region="WAR">
          <CONTACT email="jasnek@plywanielegia.pl" name="Peńsko" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="3434">
              <RESULTS>
                <RESULT eventid="1200" points="576" reactiontime="+62" swimtime="00:00:27.17" resultid="3435" heatid="7460" lane="1" entrytime="00:00:27.27" />
                <RESULT comment="Rekord Polski Masters" eventid="1436" points="585" reactiontime="+77" swimtime="00:00:26.06" resultid="3436" heatid="7647" lane="1" entrytime="00:00:26.26" />
                <RESULT comment="Rekord Polski Masters" eventid="1470" points="560" reactiontime="+63" swimtime="00:00:59.35" resultid="3437" heatid="7674" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="573" reactiontime="+79" swimtime="00:00:58.34" resultid="3438" heatid="7751" lane="3" entrytime="00:00:59.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="3439" heatid="7774" lane="3" entrytime="00:02:11.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-26" firstname="Tomasz" gender="M" lastname="Wilczęga" nation="POL" athleteid="3440">
              <RESULTS>
                <RESULT eventid="1075" points="460" reactiontime="+73" swimtime="00:00:26.29" resultid="3441" heatid="7376" lane="4" entrytime="00:00:26.43" />
                <RESULT eventid="1436" points="438" reactiontime="+72" swimtime="00:00:28.69" resultid="6444" heatid="7644" lane="3" entrytime="00:00:27.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" athleteid="3442">
              <RESULTS>
                <RESULT eventid="1075" points="414" reactiontime="+76" swimtime="00:00:27.23" resultid="3443" heatid="7376" lane="3" entrytime="00:00:26.43" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-21" firstname="Krzysztof" gender="M" lastname="Spyra" nation="POL" athleteid="3444">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="3445" heatid="7376" lane="2" entrytime="00:00:26.43" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1528" points="480" reactiontime="+80" swimtime="00:01:43.13" resultid="3446" heatid="7716" lane="2" entrytime="00:01:43.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.47" />
                    <SPLIT distance="100" swimtime="00:00:53.23" />
                    <SPLIT distance="150" swimtime="00:01:18.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3444" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3442" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3440" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="3434" number="4" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" name="MKP Szczecin" nation="POL" region="ZAC">
          <CONTACT city="Szczecin" email="windmuhle@wp.pl" name="Kowalczyk Piotr" phone="509758055" street="Kaliny 45/9" zip="71-118" />
          <ATHLETES>
            <ATHLETE birthdate="1974-02-10" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="3451">
              <RESULTS>
                <RESULT eventid="1165" points="372" reactiontime="+90" swimtime="00:19:41.02" resultid="3452" heatid="7916" lane="1" entrytime="00:19:17.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:46.88" />
                    <SPLIT distance="200" swimtime="00:02:24.86" />
                    <SPLIT distance="250" swimtime="00:03:02.75" />
                    <SPLIT distance="300" swimtime="00:03:41.30" />
                    <SPLIT distance="350" swimtime="00:04:20.47" />
                    <SPLIT distance="400" swimtime="00:05:00.03" />
                    <SPLIT distance="450" swimtime="00:05:39.99" />
                    <SPLIT distance="500" swimtime="00:06:19.97" />
                    <SPLIT distance="550" swimtime="00:07:00.23" />
                    <SPLIT distance="600" swimtime="00:07:40.17" />
                    <SPLIT distance="650" swimtime="00:08:20.15" />
                    <SPLIT distance="700" swimtime="00:09:00.38" />
                    <SPLIT distance="750" swimtime="00:09:40.01" />
                    <SPLIT distance="800" swimtime="00:10:20.09" />
                    <SPLIT distance="850" swimtime="00:10:59.78" />
                    <SPLIT distance="900" swimtime="00:11:39.89" />
                    <SPLIT distance="950" swimtime="00:12:20.67" />
                    <SPLIT distance="1000" swimtime="00:13:00.61" />
                    <SPLIT distance="1050" swimtime="00:13:41.24" />
                    <SPLIT distance="1100" swimtime="00:14:21.90" />
                    <SPLIT distance="1150" swimtime="00:15:02.21" />
                    <SPLIT distance="1200" swimtime="00:15:42.90" />
                    <SPLIT distance="1250" swimtime="00:16:23.71" />
                    <SPLIT distance="1300" swimtime="00:17:04.30" />
                    <SPLIT distance="1350" swimtime="00:17:44.36" />
                    <SPLIT distance="1400" swimtime="00:18:24.19" />
                    <SPLIT distance="1450" swimtime="00:19:04.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="396" reactiontime="+87" swimtime="00:01:01.18" resultid="3453" heatid="7519" lane="1" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="348" swimtime="00:02:21.14" resultid="3454" heatid="7702" lane="5" entrytime="00:02:14.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="150" swimtime="00:01:45.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="3455" heatid="7771" lane="5" entrytime="00:02:36.00" />
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="3456" heatid="8055" lane="2" entrytime="00:04:49.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="3457">
              <RESULTS>
                <RESULT eventid="1109" points="182" reactiontime="+93" swimtime="00:03:14.22" resultid="3458" heatid="7395" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:30.58" />
                    <SPLIT distance="150" swimtime="00:02:26.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="197" reactiontime="+94" swimtime="00:03:27.08" resultid="3459" heatid="7476" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:38.71" />
                    <SPLIT distance="150" swimtime="00:02:32.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="227" reactiontime="+82" swimtime="00:01:31.16" resultid="3460" heatid="7599" lane="1" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="232" reactiontime="+81" swimtime="00:00:41.05" resultid="3461" heatid="7798" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="3468">
              <RESULTS>
                <RESULT eventid="1058" points="420" reactiontime="+74" swimtime="00:00:31.04" resultid="3469" heatid="7342" lane="3" entrytime="00:00:30.98" />
                <RESULT eventid="1148" points="409" reactiontime="+75" swimtime="00:10:52.69" resultid="3470" heatid="7906" lane="4" entrytime="00:10:28.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:13.95" />
                    <SPLIT distance="150" swimtime="00:01:53.72" />
                    <SPLIT distance="200" swimtime="00:02:34.00" />
                    <SPLIT distance="250" swimtime="00:03:14.70" />
                    <SPLIT distance="300" swimtime="00:03:55.76" />
                    <SPLIT distance="350" swimtime="00:04:37.05" />
                    <SPLIT distance="400" swimtime="00:05:18.38" />
                    <SPLIT distance="450" swimtime="00:05:59.87" />
                    <SPLIT distance="500" swimtime="00:06:41.51" />
                    <SPLIT distance="550" swimtime="00:07:23.27" />
                    <SPLIT distance="600" swimtime="00:08:05.34" />
                    <SPLIT distance="650" swimtime="00:08:47.31" />
                    <SPLIT distance="700" swimtime="00:09:29.27" />
                    <SPLIT distance="750" swimtime="00:10:11.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="396" reactiontime="+77" swimtime="00:01:09.42" resultid="3471" heatid="7497" lane="6" entrytime="00:01:06.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="319" reactiontime="+81" swimtime="00:01:24.45" resultid="3472" heatid="7534" lane="4" entrytime="00:01:19.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="313" reactiontime="+83" swimtime="00:01:21.26" resultid="3473" heatid="7657" lane="1" entrytime="00:01:17.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="387" reactiontime="+80" swimtime="00:02:32.49" resultid="3474" heatid="7684" lane="2" entrytime="00:02:24.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:01:13.35" />
                    <SPLIT distance="150" swimtime="00:01:53.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="316" reactiontime="+84" swimtime="00:02:56.07" resultid="3475" heatid="7760" lane="1" entrytime="00:02:52.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                    <SPLIT distance="100" swimtime="00:01:25.26" />
                    <SPLIT distance="150" swimtime="00:02:10.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="388" reactiontime="+79" swimtime="00:05:21.94" resultid="3476" heatid="8024" lane="3" entrytime="00:05:12.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="150" swimtime="00:01:55.83" />
                    <SPLIT distance="200" swimtime="00:02:37.23" />
                    <SPLIT distance="250" swimtime="00:03:18.82" />
                    <SPLIT distance="300" swimtime="00:04:00.35" />
                    <SPLIT distance="350" swimtime="00:04:41.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-27" firstname="Szymon" gender="M" lastname="Kluczyk" nation="POL" athleteid="3477">
              <RESULTS>
                <RESULT eventid="1165" points="439" reactiontime="+96" swimtime="00:18:38.23" resultid="3478" heatid="7916" lane="4" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:44.67" />
                    <SPLIT distance="200" swimtime="00:02:21.03" />
                    <SPLIT distance="250" swimtime="00:02:57.62" />
                    <SPLIT distance="300" swimtime="00:03:34.39" />
                    <SPLIT distance="350" swimtime="00:04:11.25" />
                    <SPLIT distance="400" swimtime="00:04:48.38" />
                    <SPLIT distance="450" swimtime="00:05:25.35" />
                    <SPLIT distance="500" swimtime="00:06:02.58" />
                    <SPLIT distance="550" swimtime="00:06:39.72" />
                    <SPLIT distance="600" swimtime="00:07:16.89" />
                    <SPLIT distance="650" swimtime="00:07:54.34" />
                    <SPLIT distance="700" swimtime="00:08:31.94" />
                    <SPLIT distance="750" swimtime="00:09:09.49" />
                    <SPLIT distance="800" swimtime="00:09:47.05" />
                    <SPLIT distance="850" swimtime="00:10:24.93" />
                    <SPLIT distance="900" swimtime="00:11:02.64" />
                    <SPLIT distance="950" swimtime="00:11:40.43" />
                    <SPLIT distance="1000" swimtime="00:12:18.58" />
                    <SPLIT distance="1050" swimtime="00:12:56.89" />
                    <SPLIT distance="1100" swimtime="00:13:34.88" />
                    <SPLIT distance="1150" swimtime="00:14:12.96" />
                    <SPLIT distance="1200" swimtime="00:14:50.66" />
                    <SPLIT distance="1250" swimtime="00:15:28.57" />
                    <SPLIT distance="1300" swimtime="00:16:06.30" />
                    <SPLIT distance="1350" swimtime="00:16:43.92" />
                    <SPLIT distance="1400" swimtime="00:17:22.47" />
                    <SPLIT distance="1450" swimtime="00:18:00.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="382" reactiontime="+89" swimtime="00:02:30.31" resultid="3479" heatid="7570" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:11.12" />
                    <SPLIT distance="150" swimtime="00:01:50.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="403" reactiontime="+91" swimtime="00:05:18.58" resultid="3480" heatid="7982" lane="4" entrytime="00:05:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="150" swimtime="00:01:53.80" />
                    <SPLIT distance="200" swimtime="00:02:33.64" />
                    <SPLIT distance="250" swimtime="00:03:20.22" />
                    <SPLIT distance="300" swimtime="00:04:06.66" />
                    <SPLIT distance="350" swimtime="00:04:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="3481" heatid="7750" lane="2" entrytime="00:01:05.00" />
                <RESULT eventid="1710" points="441" reactiontime="+85" swimtime="00:04:39.33" resultid="3482" heatid="8057" lane="4" entrytime="00:04:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:05.32" />
                    <SPLIT distance="150" swimtime="00:01:40.23" />
                    <SPLIT distance="200" swimtime="00:02:16.14" />
                    <SPLIT distance="250" swimtime="00:02:52.42" />
                    <SPLIT distance="300" swimtime="00:03:28.47" />
                    <SPLIT distance="350" swimtime="00:04:04.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-01-01" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="3483">
              <RESULTS>
                <RESULT eventid="1217" points="103" swimtime="00:04:46.72" resultid="3484" heatid="7462" lane="3" entrytime="00:04:55.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.63" />
                    <SPLIT distance="100" swimtime="00:02:23.22" />
                    <SPLIT distance="150" swimtime="00:03:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="97" swimtime="00:02:16.44" resultid="3485" heatid="7582" lane="4" entrytime="00:02:16.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="94" swimtime="00:01:03.33" resultid="3486" heatid="7776" lane="2" entrytime="00:01:05.72" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MSWIM" name="Mswim Szczecin" nation="POL">
          <CONTACT email="m@mswim.pl" internet="www.mswim.pl" name="kaczanowski" phone="888181234" />
          <ATHLETES>
            <ATHLETE birthdate="1968-05-22" firstname="Miłosz" gender="M" lastname="kaczanowski" nation="POL" athleteid="3488">
              <RESULTS>
                <RESULT eventid="1075" points="429" reactiontime="+82" swimtime="00:00:26.90" resultid="3489" heatid="7347" lane="1" />
                <RESULT eventid="1109" points="433" swimtime="00:02:25.42" resultid="3490" heatid="7405" lane="5" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="462" reactiontime="+77" swimtime="00:00:58.11" resultid="3491" heatid="7499" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="446" swimtime="00:01:06.41" resultid="3492" heatid="7558" lane="5" entrytime="00:01:05.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="396" reactiontime="+83" swimtime="00:01:15.68" resultid="3493" heatid="7592" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="458" reactiontime="+79" swimtime="00:00:28.27" resultid="3494" heatid="7643" lane="4" entrytime="00:00:28.01" />
                <RESULT eventid="1594" points="441" reactiontime="+80" swimtime="00:01:03.67" resultid="3495" heatid="7736" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="410" swimtime="00:00:33.97" resultid="3496" heatid="7810" lane="5" entrytime="00:00:33.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-14" firstname="anna" gender="F" lastname="frankowska" nation="POL" athleteid="3497">
              <RESULTS>
                <RESULT eventid="1217" points="244" reactiontime="+101" swimtime="00:03:35.13" resultid="3498" heatid="7461" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                    <SPLIT distance="100" swimtime="00:01:41.02" />
                    <SPLIT distance="150" swimtime="00:02:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="271" reactiontime="+100" swimtime="00:01:29.14" resultid="3499" heatid="7532" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="258" reactiontime="+93" swimtime="00:01:38.44" resultid="3500" heatid="7590" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" reactiontime="+100" status="DNF" swimtime="00:00:00.00" resultid="3501" heatid="7683" lane="6" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:23.43" />
                    <SPLIT distance="150" swimtime="00:02:10.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="257" reactiontime="+87" swimtime="00:00:45.28" resultid="3502" heatid="7785" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="jadwiga" gender="F" lastname="weber" nation="POL" athleteid="3503">
              <RESULTS>
                <RESULT eventid="1183" points="251" reactiontime="+84" swimtime="00:00:40.73" resultid="3504" heatid="7435" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="1251" points="256" swimtime="00:01:20.33" resultid="3505" heatid="7491" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="255" reactiontime="+85" swimtime="00:01:27.08" resultid="3506" heatid="7653" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="263" reactiontime="+95" swimtime="00:03:07.29" resultid="3507" heatid="7758" lane="2" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:29.60" />
                    <SPLIT distance="150" swimtime="00:02:18.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORSOPOLE" name="Odrzańskie Ratownictwo Specjalistyczne Opole" nation="POL" region="OPO" shortname="Odrzańskie Ratownictwo Specjal">
          <CONTACT email="wkania62@gmail.com" name="Kania" />
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Waldemar" gender="M" lastname="Kania" nation="POL" athleteid="3509">
              <RESULTS>
                <RESULT eventid="1165" points="262" reactiontime="+103" swimtime="00:22:08.49" resultid="3510" heatid="7913" lane="3" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:21.79" />
                    <SPLIT distance="150" swimtime="00:02:06.25" />
                    <SPLIT distance="200" swimtime="00:02:51.16" />
                    <SPLIT distance="250" swimtime="00:03:36.05" />
                    <SPLIT distance="300" swimtime="00:04:20.55" />
                    <SPLIT distance="350" swimtime="00:05:04.87" />
                    <SPLIT distance="400" swimtime="00:05:49.12" />
                    <SPLIT distance="450" swimtime="00:06:33.36" />
                    <SPLIT distance="500" swimtime="00:07:17.20" />
                    <SPLIT distance="550" swimtime="00:08:00.72" />
                    <SPLIT distance="600" swimtime="00:08:45.15" />
                    <SPLIT distance="650" swimtime="00:09:29.23" />
                    <SPLIT distance="700" swimtime="00:10:14.01" />
                    <SPLIT distance="750" swimtime="00:10:59.01" />
                    <SPLIT distance="800" swimtime="00:11:44.41" />
                    <SPLIT distance="850" swimtime="00:12:29.57" />
                    <SPLIT distance="900" swimtime="00:13:14.72" />
                    <SPLIT distance="950" swimtime="00:13:59.77" />
                    <SPLIT distance="1000" swimtime="00:14:44.63" />
                    <SPLIT distance="1050" swimtime="00:15:30.34" />
                    <SPLIT distance="1100" swimtime="00:16:15.35" />
                    <SPLIT distance="1150" swimtime="00:17:00.45" />
                    <SPLIT distance="1200" swimtime="00:17:45.18" />
                    <SPLIT distance="1250" swimtime="00:18:30.20" />
                    <SPLIT distance="1300" swimtime="00:19:14.99" />
                    <SPLIT distance="1350" swimtime="00:19:59.74" />
                    <SPLIT distance="1400" swimtime="00:20:44.40" />
                    <SPLIT distance="1450" swimtime="00:21:26.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="258" reactiontime="+95" swimtime="00:02:36.06" resultid="3511" heatid="7696" lane="4" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:14.34" />
                    <SPLIT distance="150" swimtime="00:01:55.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="3512" heatid="7765" lane="4" entrytime="00:03:25.00" />
                <RESULT eventid="1710" points="260" reactiontime="+97" swimtime="00:05:33.17" resultid="3513" heatid="8051" lane="2" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                    <SPLIT distance="150" swimtime="00:02:00.40" />
                    <SPLIT distance="200" swimtime="00:02:42.92" />
                    <SPLIT distance="250" swimtime="00:03:24.98" />
                    <SPLIT distance="300" swimtime="00:04:07.49" />
                    <SPLIT distance="350" swimtime="00:04:50.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Grzegorz" gender="M" lastname="Stanek" nation="POL" athleteid="3514">
              <RESULTS>
                <RESULT eventid="1268" points="458" swimtime="00:00:58.28" resultid="3515" heatid="7522" lane="5" entrytime="00:00:58.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="3516" heatid="7705" lane="2" entrytime="00:02:06.55" />
                <RESULT comment="Rekord Polski Masters" eventid="1710" points="455" reactiontime="+79" swimtime="00:04:36.51" resultid="3517" heatid="8057" lane="1" entrytime="00:04:39.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:07.59" />
                    <SPLIT distance="150" swimtime="00:01:42.69" />
                    <SPLIT distance="200" swimtime="00:02:17.95" />
                    <SPLIT distance="250" swimtime="00:02:52.81" />
                    <SPLIT distance="300" swimtime="00:03:27.89" />
                    <SPLIT distance="350" swimtime="00:04:02.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="3518">
              <RESULTS>
                <RESULT eventid="1092" points="383" swimtime="00:02:51.53" resultid="3519" heatid="7389" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="100" swimtime="00:01:20.43" />
                    <SPLIT distance="150" swimtime="00:02:13.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="410" reactiontime="+87" swimtime="00:01:17.69" resultid="3520" heatid="7532" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="358" reactiontime="+80" swimtime="00:01:17.75" resultid="3521" heatid="7656" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="320" swimtime="00:06:21.26" resultid="3522" heatid="7717" lane="5" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:01:33.81" />
                    <SPLIT distance="150" swimtime="00:03:10.17" />
                    <SPLIT distance="200" swimtime="00:04:04.95" />
                    <SPLIT distance="250" swimtime="00:04:59.25" />
                    <SPLIT distance="300" swimtime="00:05:41.86" />
                    <SPLIT distance="350" swimtime="00:06:21.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="326" reactiontime="+87" swimtime="00:01:19.91" resultid="3523" heatid="7733" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="333" reactiontime="+86" swimtime="00:02:53.13" resultid="3524" heatid="7759" lane="6" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:26.83" />
                    <SPLIT distance="150" swimtime="00:02:12.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="3525">
              <RESULTS>
                <RESULT eventid="1092" points="298" reactiontime="+92" swimtime="00:03:06.40" resultid="3526" heatid="7387" lane="2" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:01:26.77" />
                    <SPLIT distance="150" swimtime="00:02:22.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="262" reactiontime="+77" swimtime="00:00:40.16" resultid="3527" heatid="7437" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1285" points="312" reactiontime="+96" swimtime="00:01:25.08" resultid="3528" heatid="7533" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="268" reactiontime="+74" swimtime="00:01:25.64" resultid="3529" heatid="7654" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="288" reactiontime="+77" swimtime="00:03:01.68" resultid="3530" heatid="7758" lane="3" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:28.25" />
                    <SPLIT distance="150" swimtime="00:02:15.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Mariusz" gender="M" lastname="Kowalczyk" nation="POL" athleteid="3531">
              <RESULTS>
                <RESULT eventid="1710" points="219" reactiontime="+95" swimtime="00:05:52.56" resultid="3532" heatid="8050" lane="3" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:18.77" />
                    <SPLIT distance="150" swimtime="00:02:03.13" />
                    <SPLIT distance="200" swimtime="00:02:49.03" />
                    <SPLIT distance="250" swimtime="00:03:36.10" />
                    <SPLIT distance="300" swimtime="00:04:23.57" />
                    <SPLIT distance="350" swimtime="00:05:11.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="3533">
              <RESULTS>
                <RESULT eventid="1336" status="DNS" swimtime="00:00:00.00" resultid="3534" heatid="7570" lane="4" entrytime="00:02:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" name="KS Masters Polkowice" nation="POL" region="DOL">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="ul.Kolejowa 6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1952-05-30" firstname="Grażyna" gender="F" lastname="Grzegorzewska" nation="POL" athleteid="3537">
              <RESULTS>
                <RESULT eventid="1058" points="186" reactiontime="+89" swimtime="00:00:40.72" resultid="3538" heatid="7334" lane="3" entrytime="00:00:40.80" entrycourse="SCM" />
                <RESULT eventid="1148" points="147" reactiontime="+94" swimtime="00:15:18.00" resultid="3539" heatid="7902" lane="3" entrytime="00:15:02.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                    <SPLIT distance="100" swimtime="00:01:45.46" />
                    <SPLIT distance="150" swimtime="00:02:43.67" />
                    <SPLIT distance="200" swimtime="00:03:42.07" />
                    <SPLIT distance="250" swimtime="00:04:39.48" />
                    <SPLIT distance="300" swimtime="00:05:38.15" />
                    <SPLIT distance="350" swimtime="00:06:37.06" />
                    <SPLIT distance="400" swimtime="00:07:35.38" />
                    <SPLIT distance="450" swimtime="00:08:33.89" />
                    <SPLIT distance="500" swimtime="00:09:32.33" />
                    <SPLIT distance="550" swimtime="00:10:30.96" />
                    <SPLIT distance="600" swimtime="00:11:29.73" />
                    <SPLIT distance="650" swimtime="00:12:28.03" />
                    <SPLIT distance="700" swimtime="00:13:26.12" />
                    <SPLIT distance="750" swimtime="00:14:25.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="136" reactiontime="+90" swimtime="00:01:39.19" resultid="3540" heatid="7489" lane="4" entrytime="00:01:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="113" swimtime="00:01:59.27" resultid="3541" heatid="7527" lane="5" entrytime="00:01:56.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="89" reactiontime="+87" swimtime="00:00:54.42" resultid="3542" heatid="7613" lane="4" entrytime="00:00:53.70" entrycourse="SCM" />
                <RESULT eventid="1487" points="137" reactiontime="+90" swimtime="00:03:35.34" resultid="3543" heatid="7677" lane="1" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.57" />
                    <SPLIT distance="100" swimtime="00:01:42.34" />
                    <SPLIT distance="150" swimtime="00:02:39.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="90" swimtime="00:02:02.41" resultid="3544" heatid="7731" lane="5" entrytime="00:02:03.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="148" reactiontime="+89" swimtime="00:07:23.42" resultid="3545" heatid="8020" lane="1" entrytime="00:07:21.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                    <SPLIT distance="100" swimtime="00:01:42.91" />
                    <SPLIT distance="150" swimtime="00:02:40.00" />
                    <SPLIT distance="200" swimtime="00:03:37.25" />
                    <SPLIT distance="250" swimtime="00:04:34.49" />
                    <SPLIT distance="300" swimtime="00:05:31.97" />
                    <SPLIT distance="350" swimtime="00:06:29.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-10-02" firstname="Emilia" gender="F" lastname="Kawula" nation="POL" athleteid="3546">
              <RESULTS>
                <RESULT eventid="1058" points="17" swimtime="00:01:29.31" resultid="3547" heatid="7331" lane="4" />
                <RESULT eventid="1217" points="27" swimtime="00:07:28.15" resultid="3548" heatid="7461" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.73" />
                    <SPLIT distance="100" swimtime="00:03:42.77" />
                    <SPLIT distance="150" swimtime="00:05:36.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="12" swimtime="00:03:38.64" resultid="3549" heatid="7486" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:44.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="22" swimtime="00:03:41.32" resultid="3550" heatid="7582" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="25" swimtime="00:01:38.34" resultid="3551" heatid="7775" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-10-10" firstname="Zdzisława" gender="F" lastname="Pachom" nation="POL" athleteid="3552">
              <RESULTS>
                <RESULT eventid="1058" points="20" reactiontime="+139" swimtime="00:01:25.41" resultid="3553" heatid="7331" lane="1" />
                <RESULT eventid="1251" points="21" reactiontime="+147" swimtime="00:03:02.51" resultid="3554" heatid="7486" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="24" reactiontime="+88" swimtime="00:03:18.61" resultid="3555" heatid="7526" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="22" reactiontime="+145" swimtime="00:03:42.78" resultid="3556" heatid="7581" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:46.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="15" reactiontime="+95" swimtime="00:01:36.81" resultid="3557" heatid="7612" lane="4" />
                <RESULT eventid="1645" points="25" reactiontime="+112" swimtime="00:01:37.99" resultid="3558" heatid="7775" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-23" firstname="Józefa" gender="F" lastname="Wołoszczuk" nation="POL" athleteid="3559">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="3560" heatid="7332" lane="5" />
                <RESULT eventid="1183" status="DNS" swimtime="00:00:00.00" resultid="3561" heatid="7431" lane="2" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="3562" heatid="7486" lane="6" />
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="3563" heatid="7648" lane="4" />
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="3564" heatid="7753" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-11-28" firstname="Hanna" gender="F" lastname="Świder" nation="POL" athleteid="3565">
              <RESULTS>
                <RESULT eventid="1058" points="28" swimtime="00:01:16.26" resultid="3566" heatid="7331" lane="2" />
                <RESULT eventid="1217" points="72" swimtime="00:05:22.46" resultid="3567" heatid="7461" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.18" />
                    <SPLIT distance="100" swimtime="00:02:34.85" />
                    <SPLIT distance="150" swimtime="00:03:57.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="33" swimtime="00:02:39.01" resultid="3568" heatid="7486" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="65" swimtime="00:02:35.85" resultid="3569" heatid="7581" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="59" swimtime="00:01:13.64" resultid="3570" heatid="7775" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-15" firstname="Regina" gender="F" lastname="Mładszew" nation="POL" athleteid="3571">
              <RESULTS>
                <RESULT eventid="1058" points="40" reactiontime="+96" swimtime="00:01:07.69" resultid="3572" heatid="7331" lane="3" />
                <RESULT eventid="1183" points="51" reactiontime="+161" swimtime="00:01:09.28" resultid="3573" heatid="7431" lane="4" />
                <RESULT eventid="1285" points="38" swimtime="00:02:51.17" resultid="3574" heatid="7526" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="43" reactiontime="+161" swimtime="00:02:36.59" resultid="3575" heatid="7648" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="48" reactiontime="+183" swimtime="00:05:29.38" resultid="3576" heatid="7754" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.32" />
                    <SPLIT distance="100" swimtime="00:02:43.14" />
                    <SPLIT distance="150" swimtime="00:04:08.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="28" swimtime="00:01:34.16" resultid="3577" heatid="7775" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-02" firstname="Pavlo" gender="M" lastname="Vechirko" nation="POL" athleteid="3578">
              <RESULTS>
                <RESULT eventid="1234" points="291" reactiontime="+100" swimtime="00:03:01.96" resultid="3579" heatid="7481" lane="1" entrytime="00:02:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:01:29.00" />
                    <SPLIT distance="150" swimtime="00:02:15.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="296" reactiontime="+81" swimtime="00:01:23.41" resultid="3580" heatid="7606" lane="4" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="267" reactiontime="+80" swimtime="00:01:15.91" resultid="3581" heatid="7669" lane="1" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="279" reactiontime="+80" swimtime="00:02:42.24" resultid="3582" heatid="7770" lane="5" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                    <SPLIT distance="150" swimtime="00:02:01.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-07-27" firstname="Czesław" gender="M" lastname="Kawałko" nation="POL" athleteid="3583">
              <RESULTS>
                <RESULT eventid="1075" points="34" reactiontime="+131" swimtime="00:01:02.30" resultid="3584" heatid="7346" lane="2" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="3585" heatid="7390" lane="4" />
                <RESULT eventid="1234" points="22" reactiontime="+118" swimtime="00:07:06.23" resultid="3586" heatid="7470" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:32.07" />
                    <SPLIT distance="100" swimtime="00:03:20.92" />
                    <SPLIT distance="150" swimtime="00:05:11.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="16" swimtime="00:03:20.73" resultid="3587" heatid="7538" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="13" reactiontime="+126" swimtime="00:03:26.63" resultid="3588" heatid="7659" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="16" reactiontime="+116" swimtime="00:06:54.63" resultid="3589" heatid="7763" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:40.51" />
                    <SPLIT distance="100" swimtime="00:03:24.19" />
                    <SPLIT distance="150" swimtime="00:05:10.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="22" swimtime="00:01:28.96" resultid="3590" heatid="7789" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-04-23" firstname="Bogdan" gender="M" lastname="Jawor" nation="POL" athleteid="3591">
              <RESULTS>
                <RESULT eventid="1075" points="101" reactiontime="+94" swimtime="00:00:43.56" resultid="3592" heatid="7349" lane="1" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="1109" points="76" swimtime="00:04:19.29" resultid="3593" heatid="7392" lane="5" entrytime="00:04:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.52" />
                    <SPLIT distance="100" swimtime="00:02:08.72" />
                    <SPLIT distance="150" swimtime="00:03:20.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="99" reactiontime="+91" swimtime="00:04:20.76" resultid="3594" heatid="7472" lane="1" entrytime="00:04:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.13" />
                    <SPLIT distance="100" swimtime="00:02:04.75" />
                    <SPLIT distance="150" swimtime="00:03:14.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="76" reactiontime="+92" swimtime="00:01:59.59" resultid="3595" heatid="7539" lane="3" entrytime="00:01:57.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="97" reactiontime="+98" swimtime="00:02:00.63" resultid="3596" heatid="7594" lane="3" entrytime="00:01:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="69" reactiontime="+97" swimtime="00:09:33.00" resultid="3597" heatid="7975" lane="6" entrytime="00:09:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.95" />
                    <SPLIT distance="100" swimtime="00:02:29.99" />
                    <SPLIT distance="150" swimtime="00:03:45.92" />
                    <SPLIT distance="200" swimtime="00:04:57.32" />
                    <SPLIT distance="250" swimtime="00:06:12.41" />
                    <SPLIT distance="300" swimtime="00:07:25.69" />
                    <SPLIT distance="350" swimtime="00:08:29.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="68" reactiontime="+76" swimtime="00:04:19.63" resultid="3598" heatid="7764" lane="6" entrytime="00:04:34.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.65" />
                    <SPLIT distance="100" swimtime="00:02:08.96" />
                    <SPLIT distance="150" swimtime="00:03:15.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="107" reactiontime="+97" swimtime="00:00:53.16" resultid="3599" heatid="7791" lane="3" entrytime="00:00:51.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Rydułtowska Akademia Aktywnego Seniora 60+" nation="POL" region="SLA" shortname="Rydułtowska Akademia Aktywnego">
          <CONTACT email="zurekt@poczta.onet.pl" name="Żurczak Tomasz" phone="504152136" />
          <ATHLETES>
            <ATHLETE birthdate="1951-09-07" firstname="Leon" gender="M" lastname="Irczyk" nation="POL" athleteid="3601">
              <RESULTS>
                <RESULT eventid="1109" points="95" swimtime="00:04:00.79" resultid="3602" heatid="7393" lane="5" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.61" />
                    <SPLIT distance="100" swimtime="00:02:10.74" />
                    <SPLIT distance="150" swimtime="00:03:07.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="3603" heatid="7908" lane="5" entrytime="00:31:05.00" />
                <RESULT eventid="1234" points="155" reactiontime="+117" swimtime="00:03:44.35" resultid="3604" heatid="7473" lane="2" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.13" />
                    <SPLIT distance="100" swimtime="00:01:47.97" />
                    <SPLIT distance="150" swimtime="00:02:46.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="67" reactiontime="+112" swimtime="00:04:28.59" resultid="3605" heatid="7566" lane="6" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.13" />
                    <SPLIT distance="100" swimtime="00:02:08.21" />
                    <SPLIT distance="150" swimtime="00:03:18.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="143" swimtime="00:01:46.25" resultid="3606" heatid="7596" lane="5" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="94" reactiontime="+111" swimtime="00:08:36.61" resultid="3607" heatid="7975" lane="4" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.04" />
                    <SPLIT distance="100" swimtime="00:02:07.85" />
                    <SPLIT distance="150" swimtime="00:03:25.14" />
                    <SPLIT distance="200" swimtime="00:04:38.78" />
                    <SPLIT distance="250" swimtime="00:05:40.20" />
                    <SPLIT distance="300" swimtime="00:06:40.70" />
                    <SPLIT distance="350" swimtime="00:07:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="151" reactiontime="+101" swimtime="00:00:47.39" resultid="3608" heatid="7792" lane="3" entrytime="00:00:47.25" />
                <RESULT eventid="1710" points="102" reactiontime="+134" swimtime="00:07:35.04" resultid="3609" heatid="8045" lane="2" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.96" />
                    <SPLIT distance="100" swimtime="00:01:51.21" />
                    <SPLIT distance="150" swimtime="00:02:49.51" />
                    <SPLIT distance="200" swimtime="00:03:47.45" />
                    <SPLIT distance="250" swimtime="00:04:44.77" />
                    <SPLIT distance="300" swimtime="00:05:42.62" />
                    <SPLIT distance="350" swimtime="00:06:40.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="3610">
              <RESULTS>
                <RESULT eventid="1075" points="84" reactiontime="+103" swimtime="00:00:46.29" resultid="3611" heatid="7350" lane="6" entrytime="00:00:40.05" />
                <RESULT eventid="1109" points="77" reactiontime="+112" swimtime="00:04:18.12" resultid="3612" heatid="7392" lane="3" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.20" />
                    <SPLIT distance="100" swimtime="00:02:07.48" />
                    <SPLIT distance="150" swimtime="00:03:16.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="68" reactiontime="+79" swimtime="00:00:55.26" resultid="3613" heatid="7443" lane="4" entrytime="00:00:56.05" />
                <RESULT eventid="1336" points="59" reactiontime="+119" swimtime="00:04:39.04" resultid="3614" heatid="7566" lane="1" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.71" />
                    <SPLIT distance="100" swimtime="00:02:13.42" />
                    <SPLIT distance="150" swimtime="00:03:25.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="3615" heatid="7625" lane="6" entrytime="00:00:48.00" />
                <RESULT eventid="1559" points="75" reactiontime="+110" swimtime="00:09:18.05" resultid="3616" heatid="7975" lane="2" entrytime="00:09:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.42" />
                    <SPLIT distance="100" swimtime="00:02:10.15" />
                    <SPLIT distance="150" swimtime="00:03:23.73" />
                    <SPLIT distance="200" swimtime="00:04:38.49" />
                    <SPLIT distance="250" swimtime="00:05:50.99" />
                    <SPLIT distance="300" swimtime="00:07:02.22" />
                    <SPLIT distance="350" swimtime="00:08:10.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="55" reactiontime="+106" swimtime="00:02:06.76" resultid="3617" heatid="7738" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="101" reactiontime="+103" swimtime="00:00:54.09" resultid="3618" heatid="7791" lane="2" entrytime="00:00:52.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-02-02" firstname="Maria" gender="F" lastname="Lippa" nation="POL" athleteid="3619">
              <RESULTS>
                <RESULT comment="Przekroczony limit czasu. (19:45.00)" eventid="1148" status="DSQ" swimtime="00:00:00.00" resultid="3620" heatid="7902" lane="5" entrytime="00:19:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.15" />
                    <SPLIT distance="100" swimtime="00:02:41.69" />
                    <SPLIT distance="150" swimtime="00:04:06.79" />
                    <SPLIT distance="200" swimtime="00:05:33.67" />
                    <SPLIT distance="250" swimtime="00:06:59.73" />
                    <SPLIT distance="300" swimtime="00:08:26.31" />
                    <SPLIT distance="350" swimtime="00:09:52.79" />
                    <SPLIT distance="400" swimtime="00:11:21.14" />
                    <SPLIT distance="450" swimtime="00:12:50.19" />
                    <SPLIT distance="500" swimtime="00:14:16.32" />
                    <SPLIT distance="550" swimtime="00:15:43.27" />
                    <SPLIT distance="600" swimtime="00:17:07.96" />
                    <SPLIT distance="650" swimtime="00:18:37.26" />
                    <SPLIT distance="700" swimtime="00:20:04.21" />
                    <SPLIT distance="750" swimtime="00:21:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="30" reactiontime="+139" swimtime="00:05:55.42" resultid="3621" heatid="7675" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.90" />
                    <SPLIT distance="100" swimtime="00:02:49.91" />
                    <SPLIT distance="150" swimtime="00:04:23.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="37" reactiontime="+151" swimtime="00:11:39.57" resultid="3622" heatid="8018" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.10" />
                    <SPLIT distance="100" swimtime="00:02:41.60" />
                    <SPLIT distance="150" swimtime="00:04:12.13" />
                    <SPLIT distance="200" swimtime="00:05:39.34" />
                    <SPLIT distance="250" swimtime="00:07:10.58" />
                    <SPLIT distance="300" swimtime="00:08:40.19" />
                    <SPLIT distance="350" swimtime="00:10:10.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-26" firstname="Władysław" gender="M" lastname="Szurek" nation="POL" athleteid="3623">
              <RESULTS>
                <RESULT eventid="1075" points="28" reactiontime="+188" swimtime="00:01:06.57" resultid="3624" heatid="7346" lane="4" />
                <RESULT eventid="1268" points="22" swimtime="00:02:38.91" resultid="3625" heatid="7500" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="3626" heatid="7687" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-08-10" firstname="Jan" gender="M" lastname="Klapsia" nation="POL" athleteid="3627">
              <RESULTS>
                <RESULT eventid="1075" points="21" swimtime="00:01:13.09" resultid="3628" heatid="7347" lane="5" />
                <RESULT eventid="1200" points="21" swimtime="00:01:21.00" resultid="3629" heatid="7442" lane="2" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="3630" heatid="7500" lane="2" />
                <RESULT comment="K-16 - Brak wynurzenia części głowy w czacie każdego pełnego cyklu ruchu (ramion i nóg)" eventid="1402" reactiontime="+124" status="DSQ" swimtime="00:03:26.16" resultid="3631" heatid="7592" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="3632" heatid="7659" lane="3" />
                <RESULT eventid="1662" points="28" reactiontime="+113" swimtime="00:01:23.15" resultid="3633" heatid="7789" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-08" firstname="Marian" gender="M" lastname="Otlik" nation="POL" athleteid="3634">
              <RESULTS>
                <RESULT eventid="1075" points="323" reactiontime="+71" swimtime="00:00:29.56" resultid="3635" heatid="7362" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="3636" heatid="7395" lane="6" entrytime="00:03:30.00" />
                <RESULT eventid="1268" points="301" reactiontime="+73" swimtime="00:01:06.99" resultid="3637" heatid="7509" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="233" reactiontime="+80" swimtime="00:01:22.43" resultid="3638" heatid="7543" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="227" reactiontime="+79" swimtime="00:00:35.72" resultid="3639" heatid="7630" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1504" points="235" reactiontime="+86" swimtime="00:02:40.85" resultid="3640" heatid="7694" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:01:16.73" />
                    <SPLIT distance="150" swimtime="00:02:00.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="164" reactiontime="+95" swimtime="00:01:28.56" resultid="3641" heatid="7741" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="210" reactiontime="+95" swimtime="00:05:57.54" resultid="3642" heatid="8048" lane="3" entrytime="00:06:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:20.09" />
                    <SPLIT distance="150" swimtime="00:02:03.95" />
                    <SPLIT distance="200" swimtime="00:02:50.04" />
                    <SPLIT distance="250" swimtime="00:03:37.05" />
                    <SPLIT distance="300" swimtime="00:04:25.25" />
                    <SPLIT distance="350" swimtime="00:05:13.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="3643">
              <RESULTS>
                <RESULT eventid="1109" points="181" reactiontime="+87" swimtime="00:03:14.41" resultid="3644" heatid="7396" lane="6" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="150" swimtime="00:02:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="199" reactiontime="+95" swimtime="00:24:15.22" resultid="3645" heatid="7911" lane="1" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:01:26.38" />
                    <SPLIT distance="150" swimtime="00:02:13.91" />
                    <SPLIT distance="200" swimtime="00:03:01.86" />
                    <SPLIT distance="250" swimtime="00:03:50.11" />
                    <SPLIT distance="300" swimtime="00:04:38.24" />
                    <SPLIT distance="350" swimtime="00:05:27.14" />
                    <SPLIT distance="400" swimtime="00:06:15.77" />
                    <SPLIT distance="450" swimtime="00:07:05.06" />
                    <SPLIT distance="500" swimtime="00:07:53.71" />
                    <SPLIT distance="550" swimtime="00:08:43.07" />
                    <SPLIT distance="600" swimtime="00:09:31.90" />
                    <SPLIT distance="650" swimtime="00:10:21.00" />
                    <SPLIT distance="700" swimtime="00:11:09.52" />
                    <SPLIT distance="750" swimtime="00:11:58.43" />
                    <SPLIT distance="800" swimtime="00:12:47.74" />
                    <SPLIT distance="850" swimtime="00:13:37.01" />
                    <SPLIT distance="900" swimtime="00:14:26.22" />
                    <SPLIT distance="950" swimtime="00:15:15.48" />
                    <SPLIT distance="1000" swimtime="00:16:04.31" />
                    <SPLIT distance="1050" swimtime="00:16:53.54" />
                    <SPLIT distance="1100" swimtime="00:17:42.47" />
                    <SPLIT distance="1150" swimtime="00:18:31.49" />
                    <SPLIT distance="1200" swimtime="00:19:20.67" />
                    <SPLIT distance="1250" swimtime="00:20:10.05" />
                    <SPLIT distance="1300" swimtime="00:20:59.57" />
                    <SPLIT distance="1350" swimtime="00:21:48.53" />
                    <SPLIT distance="1400" swimtime="00:22:37.53" />
                    <SPLIT distance="1450" swimtime="00:23:26.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="168" reactiontime="+70" swimtime="00:00:40.95" resultid="3646" heatid="7447" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1336" points="113" reactiontime="+100" swimtime="00:03:45.58" resultid="3647" heatid="7567" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                    <SPLIT distance="100" swimtime="00:01:43.19" />
                    <SPLIT distance="150" swimtime="00:02:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="198" reactiontime="+85" swimtime="00:00:37.36" resultid="3648" heatid="7628" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1470" points="163" reactiontime="+77" swimtime="00:01:29.44" resultid="3649" heatid="7663" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="159" reactiontime="+88" swimtime="00:01:29.44" resultid="3650" heatid="7741" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="151" reactiontime="+88" swimtime="00:03:19.12" resultid="3651" heatid="7766" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                    <SPLIT distance="100" swimtime="00:01:36.32" />
                    <SPLIT distance="150" swimtime="00:02:28.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="133" reactiontime="+82" swimtime="00:02:59.56" resultid="3652" heatid="7928" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.54" />
                    <SPLIT distance="100" swimtime="00:01:48.38" />
                    <SPLIT distance="150" swimtime="00:02:27.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3610" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3601" number="2" />
                    <RELAYPOSITION athleteid="3643" number="3" />
                    <RELAYPOSITION athleteid="3634" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Sikret Gliwice" nation="POL">
          <CONTACT city="Gliwice" email="joannaeco@wp.pl" internet="www.sikret-plywanie.pl" name="ZAGAŁA JOANNA" phone="601427257" state="ŚLĄSK" street="Jagielońska 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1978-08-11" firstname="Agnieszka" gender="F" lastname="Drejka" nation="POL" athleteid="3657">
              <RESULTS>
                <RESULT eventid="1251" points="177" swimtime="00:01:30.75" resultid="3658" heatid="7490" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="182" reactiontime="+98" swimtime="00:01:50.46" resultid="3659" heatid="7585" lane="6" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="161" reactiontime="+96" swimtime="00:03:23.99" resultid="3660" heatid="7677" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:35.86" />
                    <SPLIT distance="150" swimtime="00:02:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="175" swimtime="00:00:51.40" resultid="3661" heatid="7779" lane="5" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="3662">
              <RESULTS>
                <RESULT eventid="1217" points="158" reactiontime="+87" swimtime="00:04:08.78" resultid="3663" heatid="7464" lane="1" entrytime="00:04:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.35" />
                    <SPLIT distance="100" swimtime="00:01:58.39" />
                    <SPLIT distance="150" swimtime="00:03:04.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="75" reactiontime="+96" swimtime="00:04:45.51" resultid="3664" heatid="7561" lane="3" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.01" />
                    <SPLIT distance="100" swimtime="00:02:10.41" />
                    <SPLIT distance="150" swimtime="00:03:25.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="170" reactiontime="+93" swimtime="00:01:53.10" resultid="3665" heatid="7584" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="110" reactiontime="+106" swimtime="00:00:50.74" resultid="3666" heatid="7614" lane="4" entrytime="00:00:48.00" />
                <RESULT eventid="1577" points="92" reactiontime="+92" swimtime="00:02:01.63" resultid="3667" heatid="7731" lane="2" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="187" reactiontime="+89" swimtime="00:00:50.34" resultid="3668" heatid="7780" lane="1" entrytime="00:00:49.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="3669">
              <RESULTS>
                <RESULT eventid="1058" points="241" reactiontime="+76" swimtime="00:00:37.36" resultid="3670" heatid="7332" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1092" points="162" reactiontime="+88" swimtime="00:03:48.34" resultid="3671" heatid="7383" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.34" />
                    <SPLIT distance="100" swimtime="00:01:48.57" />
                    <SPLIT distance="150" swimtime="00:02:52.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="166" reactiontime="+86" swimtime="00:04:04.52" resultid="3672" heatid="7463" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.81" />
                    <SPLIT distance="100" swimtime="00:01:57.02" />
                    <SPLIT distance="150" swimtime="00:03:01.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="185" reactiontime="+84" swimtime="00:01:41.26" resultid="3673" heatid="7527" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="3674" heatid="7583" lane="4" entrytime="00:02:10.00" />
                <RESULT eventid="1487" status="DNS" swimtime="00:00:00.00" resultid="3675" heatid="7676" lane="5" entrytime="00:03:50.00" />
                <RESULT eventid="1611" points="148" reactiontime="+76" swimtime="00:03:46.63" resultid="3676" heatid="7755" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="204" swimtime="00:00:48.90" resultid="3677" heatid="7776" lane="5" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-15" firstname="Mieczysław" gender="M" lastname="Mydłowski" nation="POL" athleteid="3678">
              <RESULTS>
                <RESULT eventid="1075" points="288" reactiontime="+92" swimtime="00:00:30.73" resultid="3679" heatid="7357" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1200" points="212" reactiontime="+75" swimtime="00:00:37.88" resultid="3680" heatid="7447" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1268" points="276" swimtime="00:01:09.01" resultid="3681" heatid="7511" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K-14 - Praca nóg w płaszczyźnie pionowej." eventid="1402" reactiontime="+92" status="DSQ" swimtime="00:01:27.83" resultid="3682" heatid="7601" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="192" reactiontime="+79" swimtime="00:01:24.81" resultid="3683" heatid="7666" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="252" reactiontime="+100" swimtime="00:00:39.95" resultid="3684" heatid="7798" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-10-06" firstname="Arkadiusz" gender="M" lastname="Bednarek" nation="POL" athleteid="3685">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="3686" heatid="7352" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1268" points="169" reactiontime="+102" swimtime="00:01:21.16" resultid="3687" heatid="7505" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="173" reactiontime="+100" swimtime="00:00:39.10" resultid="3688" heatid="7625" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1504" points="141" reactiontime="+99" swimtime="00:03:10.59" resultid="3689" heatid="7689" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:01:29.19" />
                    <SPLIT distance="150" swimtime="00:02:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K-4" eventid="1662" reactiontime="+105" status="DSQ" swimtime="00:00:43.81" resultid="3690" heatid="7794" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-10-21" firstname="Krystian" gender="M" lastname="Kapias" nation="POL" athleteid="3691">
              <RESULTS>
                <RESULT eventid="1075" points="195" swimtime="00:00:34.98" resultid="3692" heatid="7354" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1268" points="158" reactiontime="+85" swimtime="00:01:22.99" resultid="3693" heatid="7506" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-04" firstname="Paweł" gender="M" lastname="Bomastyk" nation="POL" athleteid="3694">
              <RESULTS>
                <RESULT eventid="1075" points="165" reactiontime="+83" swimtime="00:00:36.96" resultid="3695" heatid="7356" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1662" points="181" reactiontime="+103" swimtime="00:00:44.62" resultid="3696" heatid="7796" lane="1" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="206" reactiontime="+77" swimtime="00:02:35.22" resultid="3699" heatid="7930" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:21.01" />
                    <SPLIT distance="150" swimtime="00:01:59.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3678" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3694" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3685" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="3691" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="215" reactiontime="+77" swimtime="00:02:14.77" resultid="3700" heatid="7711" lane="2" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:44.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3678" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3694" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3691" number="3" reactiontime="+10" />
                    <RELAYPOSITION athleteid="3685" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1679" points="147" reactiontime="+75" swimtime="00:02:53.59" resultid="3697" heatid="7815" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="150" swimtime="00:02:20.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3678" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3669" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3662" number="3" />
                    <RELAYPOSITION athleteid="3694" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1126" points="172" swimtime="00:02:25.05" resultid="3698" heatid="7409" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:01:42.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3662" number="1" />
                    <RELAYPOSITION athleteid="3678" number="2" />
                    <RELAYPOSITION athleteid="3669" number="3" />
                    <RELAYPOSITION athleteid="3691" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00408" name="Uks Delfin Masters Tarnobrzeg" nation="POL" region="RZ">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1977-04-24" firstname="Renata" gender="F" lastname="Osmala" nation="POL" athleteid="3707">
              <RESULTS>
                <RESULT eventid="1148" points="377" reactiontime="+87" swimtime="00:11:10.64" resultid="3708" heatid="7905" lane="1" entrytime="00:11:25.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                    <SPLIT distance="150" swimtime="00:01:57.93" />
                    <SPLIT distance="200" swimtime="00:02:39.87" />
                    <SPLIT distance="250" swimtime="00:03:22.43" />
                    <SPLIT distance="300" swimtime="00:04:04.81" />
                    <SPLIT distance="350" swimtime="00:04:47.18" />
                    <SPLIT distance="400" swimtime="00:05:29.88" />
                    <SPLIT distance="450" swimtime="00:06:12.69" />
                    <SPLIT distance="500" swimtime="00:06:55.76" />
                    <SPLIT distance="550" swimtime="00:07:38.55" />
                    <SPLIT distance="600" swimtime="00:08:21.44" />
                    <SPLIT distance="650" swimtime="00:09:03.79" />
                    <SPLIT distance="700" swimtime="00:09:47.04" />
                    <SPLIT distance="750" swimtime="00:10:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="302" reactiontime="+72" swimtime="00:00:38.30" resultid="3709" heatid="7439" lane="1" entrytime="00:00:36.89" />
                <RESULT eventid="1285" points="360" reactiontime="+84" swimtime="00:01:21.10" resultid="3710" heatid="7534" lane="3" entrytime="00:01:19.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="358" reactiontime="+90" swimtime="00:01:28.29" resultid="3711" heatid="7590" lane="2" entrytime="00:01:26.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="302" reactiontime="+71" swimtime="00:01:22.28" resultid="3712" heatid="7656" lane="5" entrytime="00:01:19.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="349" reactiontime="+69" swimtime="00:02:50.33" resultid="3713" heatid="7760" lane="5" entrytime="00:02:50.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                    <SPLIT distance="100" swimtime="00:01:23.61" />
                    <SPLIT distance="150" swimtime="00:02:07.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="363" reactiontime="+89" swimtime="00:00:40.34" resultid="3714" heatid="7785" lane="3" entrytime="00:00:39.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="3715">
              <RESULTS>
                <RESULT eventid="1058" points="402" reactiontime="+87" swimtime="00:00:31.49" resultid="3716" heatid="7341" lane="6" entrytime="00:00:32.06" />
                <RESULT eventid="1251" points="398" reactiontime="+91" swimtime="00:01:09.29" resultid="3717" heatid="7495" lane="4" entrytime="00:01:10.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="360" reactiontime="+91" swimtime="00:01:21.16" resultid="3718" heatid="7534" lane="6" entrytime="00:01:21.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="290" reactiontime="+96" swimtime="00:00:36.82" resultid="3719" heatid="7618" lane="6" entrytime="00:00:37.60" />
                <RESULT eventid="1487" points="330" reactiontime="+99" swimtime="00:02:40.79" resultid="3720" heatid="7682" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="150" swimtime="00:02:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="326" reactiontime="+97" swimtime="00:05:41.31" resultid="3721" heatid="8023" lane="3" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:22.41" />
                    <SPLIT distance="150" swimtime="00:02:06.69" />
                    <SPLIT distance="200" swimtime="00:02:51.24" />
                    <SPLIT distance="250" swimtime="00:03:35.41" />
                    <SPLIT distance="300" swimtime="00:04:19.15" />
                    <SPLIT distance="350" swimtime="00:05:01.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-08-01" firstname="Monika" gender="F" lastname="Maciąg" nation="POL" athleteid="3722">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="3723" heatid="7387" lane="3" entrytime="00:03:01.40" />
                <RESULT eventid="1148" points="263" reactiontime="+106" swimtime="00:12:36.01" resultid="3724" heatid="7904" lane="4" entrytime="00:12:10.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:27.60" />
                    <SPLIT distance="150" swimtime="00:02:14.40" />
                    <SPLIT distance="200" swimtime="00:03:00.76" />
                    <SPLIT distance="250" swimtime="00:03:48.00" />
                    <SPLIT distance="300" swimtime="00:04:34.95" />
                    <SPLIT distance="350" swimtime="00:05:22.28" />
                    <SPLIT distance="400" swimtime="00:06:09.82" />
                    <SPLIT distance="450" swimtime="00:06:58.79" />
                    <SPLIT distance="500" swimtime="00:07:47.98" />
                    <SPLIT distance="550" swimtime="00:08:36.04" />
                    <SPLIT distance="600" swimtime="00:09:24.39" />
                    <SPLIT distance="650" swimtime="00:10:12.97" />
                    <SPLIT distance="700" swimtime="00:11:01.61" />
                    <SPLIT distance="750" swimtime="00:11:49.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="258" reactiontime="+67" swimtime="00:00:40.32" resultid="3725" heatid="7436" lane="5" entrytime="00:00:40.21" />
                <RESULT eventid="1285" points="284" reactiontime="+96" swimtime="00:01:27.77" resultid="3726" heatid="7531" lane="2" entrytime="00:01:25.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="264" reactiontime="+76" swimtime="00:01:26.08" resultid="3727" heatid="7654" lane="6" entrytime="00:01:26.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="276" reactiontime="+97" swimtime="00:02:50.64" resultid="3728" heatid="7681" lane="3" entrytime="00:02:47.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                    <SPLIT distance="100" swimtime="00:01:22.70" />
                    <SPLIT distance="150" swimtime="00:02:06.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="274" reactiontime="+67" swimtime="00:03:04.70" resultid="3729" heatid="7759" lane="5" entrytime="00:03:01.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                    <SPLIT distance="100" swimtime="00:01:30.31" />
                    <SPLIT distance="150" swimtime="00:02:17.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="262" reactiontime="+98" swimtime="00:06:06.96" resultid="3730" heatid="8022" lane="2" entrytime="00:05:55.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                    <SPLIT distance="100" swimtime="00:01:25.70" />
                    <SPLIT distance="150" swimtime="00:03:46.26" />
                    <SPLIT distance="200" swimtime="00:04:33.66" />
                    <SPLIT distance="250" swimtime="00:05:20.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Beata" gender="F" lastname="Kaczmarczyk" nation="POL" athleteid="3731">
              <RESULTS>
                <RESULT eventid="1058" points="280" swimtime="00:00:35.51" resultid="3732" heatid="7339" lane="5" entrytime="00:00:34.70" />
                <RESULT eventid="1183" points="246" reactiontime="+80" swimtime="00:00:40.99" resultid="3733" heatid="7436" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1251" points="281" reactiontime="+88" swimtime="00:01:17.79" resultid="3734" heatid="7493" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="248" reactiontime="+75" swimtime="00:01:27.86" resultid="3735" heatid="7652" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="259" reactiontime="+91" swimtime="00:02:54.29" resultid="3736" heatid="7680" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                    <SPLIT distance="150" swimtime="00:02:10.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="261" reactiontime="+80" swimtime="00:03:07.80" resultid="3737" heatid="7757" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                    <SPLIT distance="100" swimtime="00:01:33.52" />
                    <SPLIT distance="150" swimtime="00:02:21.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="247" reactiontime="+96" swimtime="00:06:14.29" resultid="3738" heatid="8022" lane="6" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                    <SPLIT distance="100" swimtime="00:01:26.76" />
                    <SPLIT distance="150" swimtime="00:02:14.42" />
                    <SPLIT distance="200" swimtime="00:03:02.16" />
                    <SPLIT distance="250" swimtime="00:03:50.27" />
                    <SPLIT distance="300" swimtime="00:04:38.58" />
                    <SPLIT distance="350" swimtime="00:05:26.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-17" firstname="Sławomir" gender="M" lastname="Kowalski" nation="POL" athleteid="3739">
              <RESULTS>
                <RESULT eventid="1075" points="359" swimtime="00:00:28.55" resultid="3740" heatid="7361" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1109" points="321" reactiontime="+82" swimtime="00:02:40.72" resultid="3741" heatid="7398" lane="2" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                    <SPLIT distance="150" swimtime="00:02:02.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="334" reactiontime="+77" swimtime="00:02:53.92" resultid="3742" heatid="7478" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:21.04" />
                    <SPLIT distance="150" swimtime="00:02:07.89" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1302" reactiontime="+65" status="DSQ" swimtime="00:01:12.55" resultid="3743" heatid="7547" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="368" reactiontime="+90" swimtime="00:01:17.58" resultid="3744" heatid="7605" lane="4" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="3745" heatid="7630" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1662" points="385" reactiontime="+88" swimtime="00:00:34.68" resultid="3746" heatid="7802" lane="3" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="Szklarz" nation="POL" athleteid="3747">
              <RESULTS>
                <RESULT eventid="1075" points="322" swimtime="00:00:29.59" resultid="3748" heatid="7367" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1302" points="295" swimtime="00:01:16.19" resultid="3749" heatid="7548" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="322" reactiontime="+75" swimtime="00:00:31.78" resultid="3750" heatid="7636" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="3751" heatid="7745" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1662" points="306" reactiontime="+76" swimtime="00:00:37.47" resultid="3752" heatid="7803" lane="6" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-04-09" firstname="Zbigniew" gender="M" lastname="Ramos" nation="POL" athleteid="3753">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="3754" heatid="7363" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="3755" heatid="7509" lane="6" entrytime="00:01:11.00" />
                <RESULT eventid="1402" points="310" swimtime="00:01:22.08" resultid="3756" heatid="7603" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="280" reactiontime="+92" swimtime="00:00:33.32" resultid="3757" heatid="7632" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1662" points="317" reactiontime="+90" swimtime="00:00:37.00" resultid="3758" heatid="7808" lane="4" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="3759">
              <RESULTS>
                <RESULT eventid="1075" points="414" reactiontime="+81" swimtime="00:00:27.22" resultid="3760" heatid="7367" lane="3" entrytime="00:00:28.54" />
                <RESULT eventid="1268" points="420" reactiontime="+81" swimtime="00:00:59.99" resultid="3761" heatid="7517" lane="6" entrytime="00:01:03.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="385" reactiontime="+79" swimtime="00:01:09.75" resultid="3762" heatid="7550" lane="6" entrytime="00:01:14.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="366" reactiontime="+80" swimtime="00:00:30.47" resultid="3763" heatid="7633" lane="3" entrytime="00:00:32.84" />
                <RESULT eventid="1504" points="384" reactiontime="+86" swimtime="00:02:16.62" resultid="3764" heatid="7699" lane="6" entrytime="00:02:24.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                    <SPLIT distance="150" swimtime="00:01:42.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="298" reactiontime="+83" swimtime="00:01:12.56" resultid="3765" heatid="7745" lane="4" entrytime="00:01:14.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="376" reactiontime="+80" swimtime="00:00:34.98" resultid="3766" heatid="7805" lane="3" entrytime="00:00:35.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="3767">
              <RESULTS>
                <RESULT eventid="1075" points="289" swimtime="00:00:30.68" resultid="3768" heatid="7362" lane="5" entrytime="00:00:30.25" />
                <RESULT eventid="1165" points="251" reactiontime="+86" swimtime="00:22:25.95" resultid="3769" heatid="7911" lane="3" entrytime="00:23:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="150" swimtime="00:02:01.93" />
                    <SPLIT distance="200" swimtime="00:02:44.59" />
                    <SPLIT distance="250" swimtime="00:03:27.55" />
                    <SPLIT distance="300" swimtime="00:04:10.25" />
                    <SPLIT distance="350" swimtime="00:04:53.22" />
                    <SPLIT distance="400" swimtime="00:05:36.66" />
                    <SPLIT distance="450" swimtime="00:06:20.24" />
                    <SPLIT distance="500" swimtime="00:07:04.62" />
                    <SPLIT distance="550" swimtime="00:07:49.81" />
                    <SPLIT distance="600" swimtime="00:08:34.50" />
                    <SPLIT distance="650" swimtime="00:09:19.58" />
                    <SPLIT distance="700" swimtime="00:10:05.63" />
                    <SPLIT distance="750" swimtime="00:10:51.93" />
                    <SPLIT distance="800" swimtime="00:11:38.87" />
                    <SPLIT distance="850" swimtime="00:12:25.42" />
                    <SPLIT distance="900" swimtime="00:13:11.93" />
                    <SPLIT distance="950" swimtime="00:13:58.31" />
                    <SPLIT distance="1000" swimtime="00:14:45.26" />
                    <SPLIT distance="1050" swimtime="00:15:31.15" />
                    <SPLIT distance="1100" swimtime="00:16:18.23" />
                    <SPLIT distance="1150" swimtime="00:17:04.62" />
                    <SPLIT distance="1200" swimtime="00:17:51.97" />
                    <SPLIT distance="1250" swimtime="00:18:37.89" />
                    <SPLIT distance="1300" swimtime="00:19:25.32" />
                    <SPLIT distance="1350" swimtime="00:20:11.49" />
                    <SPLIT distance="1400" swimtime="00:20:58.64" />
                    <SPLIT distance="1450" swimtime="00:21:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="294" reactiontime="+77" swimtime="00:01:07.53" resultid="3770" heatid="7510" lane="3" entrytime="00:01:09.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="248" reactiontime="+84" swimtime="00:00:34.66" resultid="3771" heatid="7629" lane="1" entrytime="00:00:36.25" />
                <RESULT eventid="1504" points="278" reactiontime="+80" swimtime="00:02:32.19" resultid="3772" heatid="7696" lane="2" entrytime="00:02:33.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:14.25" />
                    <SPLIT distance="150" swimtime="00:01:54.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="284" reactiontime="+78" swimtime="00:05:23.63" resultid="3773" heatid="8051" lane="3" entrytime="00:05:29.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:16.28" />
                    <SPLIT distance="150" swimtime="00:01:57.58" />
                    <SPLIT distance="200" swimtime="00:02:38.82" />
                    <SPLIT distance="250" swimtime="00:03:19.82" />
                    <SPLIT distance="300" swimtime="00:04:01.53" />
                    <SPLIT distance="350" swimtime="00:04:44.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-15" firstname="Andrzej" gender="M" lastname="Brożyna" nation="POL" athleteid="3774">
              <RESULTS>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1075" reactiontime="+72" status="DSQ" swimtime="00:00:28.28" resultid="3775" heatid="7371" lane="4" entrytime="00:00:27.74" />
                <RESULT eventid="1200" points="262" reactiontime="+61" swimtime="00:00:35.29" resultid="3776" heatid="7453" lane="1" entrytime="00:00:33.44" />
                <RESULT eventid="1268" points="288" swimtime="00:01:08.05" resultid="3777" heatid="7513" lane="5" entrytime="00:01:06.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="226" reactiontime="+60" swimtime="00:01:20.25" resultid="3778" heatid="7666" lane="2" entrytime="00:01:19.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="364" reactiontime="+70" swimtime="00:02:08.50" resultid="3784" heatid="7932" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:09.00" />
                    <SPLIT distance="150" swimtime="00:01:41.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3774" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="3739" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="3753" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3759" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="360" reactiontime="+87" swimtime="00:01:53.45" resultid="3785" heatid="7715" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="100" swimtime="00:00:58.88" />
                    <SPLIT distance="150" swimtime="00:01:26.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3739" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3753" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3774" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3759" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1370" points="301" reactiontime="+70" swimtime="00:02:33.15" resultid="3779" heatid="7573" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                    <SPLIT distance="100" swimtime="00:01:20.99" />
                    <SPLIT distance="150" swimtime="00:01:58.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3722" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="3707" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3715" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3731" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1521" points="318" swimtime="00:02:16.57" resultid="3780" heatid="7708" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="150" swimtime="00:01:44.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3707" number="1" />
                    <RELAYPOSITION athleteid="3722" number="2" />
                    <RELAYPOSITION athleteid="3731" number="3" />
                    <RELAYPOSITION athleteid="3715" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1126" points="317" reactiontime="+80" swimtime="00:01:58.42" resultid="3781" heatid="7410" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:00.87" />
                    <SPLIT distance="150" swimtime="00:01:31.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3707" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3774" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="3715" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3759" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1679" points="275" reactiontime="+73" swimtime="00:02:21.08" resultid="3783" heatid="7817" lane="2" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="150" swimtime="00:01:51.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3722" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3739" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="3715" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="3767" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1126" points="259" reactiontime="+76" swimtime="00:02:06.65" resultid="3782" heatid="7410" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                    <SPLIT distance="100" swimtime="00:01:03.22" />
                    <SPLIT distance="150" swimtime="00:01:37.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3747" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3722" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="3731" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3739" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Zhytomyr Aqua Masters" nation="UKR" region="ZHTM">
          <CONTACT city="ZHYTOMYR" email="reservation007@mail.ru" fax="+380412418911" name="IGOR KUKHARYEV" phone="+380412418900" street="MOSKOVSKA str. 35, apt.4" zip="10029" />
          <ATHLETES>
            <ATHLETE birthdate="1966-11-25" firstname="Igor" gender="M" lastname="Kukharyev" nation="UKR" athleteid="3799">
              <RESULTS>
                <RESULT eventid="1109" points="293" reactiontime="+93" swimtime="00:02:45.73" resultid="3800" heatid="7400" lane="2" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="100" swimtime="00:01:16.58" />
                    <SPLIT distance="150" swimtime="00:02:09.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="321" reactiontime="+96" swimtime="00:20:40.56" resultid="3801" heatid="7916" lane="6" entrytime="00:19:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:51.36" />
                    <SPLIT distance="200" swimtime="00:02:30.54" />
                    <SPLIT distance="250" swimtime="00:03:10.09" />
                    <SPLIT distance="300" swimtime="00:03:49.69" />
                    <SPLIT distance="350" swimtime="00:04:29.56" />
                    <SPLIT distance="400" swimtime="00:05:09.74" />
                    <SPLIT distance="450" swimtime="00:05:50.54" />
                    <SPLIT distance="500" swimtime="00:06:31.33" />
                    <SPLIT distance="550" swimtime="00:07:13.12" />
                    <SPLIT distance="600" swimtime="00:07:55.19" />
                    <SPLIT distance="650" swimtime="00:08:36.44" />
                    <SPLIT distance="700" swimtime="00:09:18.45" />
                    <SPLIT distance="750" swimtime="00:10:00.56" />
                    <SPLIT distance="800" swimtime="00:10:42.68" />
                    <SPLIT distance="850" swimtime="00:11:25.48" />
                    <SPLIT distance="900" swimtime="00:12:07.82" />
                    <SPLIT distance="950" swimtime="00:12:50.69" />
                    <SPLIT distance="1000" swimtime="00:13:33.57" />
                    <SPLIT distance="1050" swimtime="00:14:16.43" />
                    <SPLIT distance="1100" swimtime="00:14:59.25" />
                    <SPLIT distance="1150" swimtime="00:15:41.91" />
                    <SPLIT distance="1200" swimtime="00:16:25.30" />
                    <SPLIT distance="1250" swimtime="00:17:08.63" />
                    <SPLIT distance="1300" swimtime="00:17:51.59" />
                    <SPLIT distance="1350" swimtime="00:18:34.78" />
                    <SPLIT distance="1400" swimtime="00:19:18.02" />
                    <SPLIT distance="1450" swimtime="00:20:00.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="271" reactiontime="+73" swimtime="00:02:43.85" resultid="3802" heatid="7769" lane="1" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                    <SPLIT distance="150" swimtime="00:02:02.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-08-01" firstname="Mykola" gender="M" lastname="Kulyk" nation="UKR" athleteid="3804">
              <RESULTS>
                <RESULT eventid="1075" points="307" reactiontime="+81" swimtime="00:00:30.09" resultid="3805" heatid="7363" lane="6" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1268" points="302" reactiontime="+84" swimtime="00:01:06.93" resultid="3806" heatid="7513" lane="6" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-10-10" firstname="Nataliia" gender="F" lastname="Ivanova" nation="UKR" athleteid="3807">
              <RESULTS>
                <RESULT eventid="1058" points="240" reactiontime="+82" swimtime="00:00:37.37" resultid="3808" heatid="7337" lane="3" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="3809" heatid="7491" lane="4" entrytime="00:01:23.00" entrycourse="SCM" />
                <RESULT eventid="1487" status="DNS" swimtime="00:00:00.00" resultid="3810" heatid="7679" lane="4" entrytime="00:02:59.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-10-10" firstname="Iryna" gender="F" lastname="Kovalchuk" nation="UKR" athleteid="3811">
              <RESULTS>
                <RESULT eventid="1217" points="225" reactiontime="+105" swimtime="00:03:41.06" resultid="3812" heatid="7465" lane="2" entrytime="00:03:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.91" />
                    <SPLIT distance="100" swimtime="00:01:49.53" />
                    <SPLIT distance="150" swimtime="00:02:46.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="224" reactiontime="+97" swimtime="00:01:43.09" resultid="3813" heatid="7586" lane="4" entrytime="00:01:42.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="230" swimtime="00:00:46.94" resultid="3814" heatid="7784" lane="5" entrytime="00:00:43.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-28" firstname="Yuriy" gender="M" lastname="Ovsiyenko" nation="UKR" athleteid="3815">
              <RESULTS>
                <RESULT eventid="1234" points="254" reactiontime="+101" swimtime="00:03:10.47" resultid="3816" heatid="7477" lane="4" entrytime="00:03:11.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:29.58" />
                    <SPLIT distance="150" swimtime="00:02:20.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="270" reactiontime="+88" swimtime="00:01:25.99" resultid="3817" heatid="7602" lane="6" entrytime="00:01:25.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="327" swimtime="00:00:36.62" resultid="3818" heatid="7804" lane="5" entrytime="00:00:36.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" name="Masters Unia Oświęcim" nation="POL" region="06">
          <ATHLETES>
            <ATHLETE birthdate="1961-03-16" firstname="Tomasz" gender="M" lastname="Dorywalski" nation="POL" athleteid="3820">
              <RESULTS>
                <RESULT eventid="1200" points="229" reactiontime="+67" swimtime="00:00:36.95" resultid="3821" heatid="7448" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1470" points="215" reactiontime="+87" swimtime="00:01:21.67" resultid="3822" heatid="7667" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="219" reactiontime="+69" swimtime="00:02:56.00" resultid="3823" heatid="7766" lane="3" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:01:24.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-11-05" firstname="Sławomir" gender="M" lastname="Formas" nation="POL" athleteid="3824">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1234" points="441" reactiontime="+90" swimtime="00:02:38.51" resultid="3825" heatid="7483" lane="2" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:01:58.55" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1402" points="481" reactiontime="+87" swimtime="00:01:10.94" resultid="3826" heatid="7609" lane="2" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1662" points="509" reactiontime="+82" swimtime="00:00:31.62" resultid="3827" heatid="7811" lane="4" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-27" firstname="Robert" gender="M" lastname="Krulikowski" nation="POL" athleteid="3828">
              <RESULTS>
                <RESULT eventid="1200" points="310" reactiontime="+73" swimtime="00:00:33.38" resultid="3829" heatid="7452" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1302" points="383" swimtime="00:01:09.86" resultid="3830" heatid="7553" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="3831" heatid="7637" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1470" points="295" reactiontime="+70" swimtime="00:01:13.47" resultid="3832" heatid="7671" lane="1" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="324" reactiontime="+70" swimtime="00:01:10.54" resultid="3833" heatid="7748" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-10" firstname="Jolanta" gender="F" lastname="Płatek" nation="POL" athleteid="3834">
              <RESULTS>
                <RESULT eventid="1183" points="326" reactiontime="+73" swimtime="00:00:37.34" resultid="3835" heatid="7439" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1453" points="308" reactiontime="+75" swimtime="00:01:21.76" resultid="3836" heatid="7654" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="307" reactiontime="+80" swimtime="00:02:57.80" resultid="3837" heatid="7759" lane="1" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="100" swimtime="00:01:27.94" />
                    <SPLIT distance="150" swimtime="00:02:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="293" reactiontime="+102" swimtime="00:05:53.30" resultid="3838" heatid="8022" lane="3" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:21.71" />
                    <SPLIT distance="150" swimtime="00:02:06.01" />
                    <SPLIT distance="200" swimtime="00:02:50.77" />
                    <SPLIT distance="250" swimtime="00:03:36.02" />
                    <SPLIT distance="300" swimtime="00:04:21.50" />
                    <SPLIT distance="350" swimtime="00:05:07.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-03" firstname="Ilona" gender="F" lastname="Szkudlarz" nation="POL" athleteid="3839">
              <RESULTS>
                <RESULT eventid="1183" points="242" reactiontime="+68" swimtime="00:00:41.20" resultid="3840" heatid="7436" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1251" points="300" reactiontime="+83" swimtime="00:01:16.17" resultid="3841" heatid="7492" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="298" swimtime="00:01:33.77" resultid="3842" heatid="7587" lane="5" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="291" reactiontime="+93" swimtime="00:02:47.67" resultid="3843" heatid="7679" lane="2" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:21.33" />
                    <SPLIT distance="150" swimtime="00:02:05.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="296" reactiontime="+90" swimtime="00:00:43.19" resultid="3844" heatid="7785" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-05" firstname="Krzysztof" gender="M" lastname="Szpara" nation="POL" athleteid="3845">
              <RESULTS>
                <RESULT eventid="1268" points="396" reactiontime="+82" swimtime="00:01:01.19" resultid="3846" heatid="7514" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="359" reactiontime="+89" swimtime="00:01:11.41" resultid="3847" heatid="7551" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="306" reactiontime="+64" swimtime="00:01:12.61" resultid="3848" heatid="7668" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="311" reactiontime="+88" swimtime="00:02:26.65" resultid="3849" heatid="7695" lane="6" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:09.78" />
                    <SPLIT distance="150" swimtime="00:01:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="307" reactiontime="+73" swimtime="00:02:37.21" resultid="3850" heatid="7768" lane="4" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:55.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="394" reactiontime="+69" swimtime="00:02:05.16" resultid="3851" heatid="7932" lane="4" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:01:07.00" />
                    <SPLIT distance="150" swimtime="00:01:37.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3820" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3824" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="3828" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="3845" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="337" reactiontime="+87" swimtime="00:01:56.04" resultid="3852" heatid="7713" lane="3" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.88" />
                    <SPLIT distance="100" swimtime="00:00:59.76" />
                    <SPLIT distance="150" swimtime="00:01:28.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3845" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3828" number="2" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3820" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3824" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1679" points="331" reactiontime="+80" swimtime="00:02:12.63" resultid="3853" heatid="7818" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:08.76" />
                    <SPLIT distance="150" swimtime="00:01:39.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3834" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3839" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3828" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3845" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Masters Wisła Kraków" nation="POL">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/" name="Wojciech Wolski" phone="791126323" />
          <ATHLETES>
            <ATHLETE birthdate="1951-09-10" firstname="Janusz" gender="M" lastname="Mrozik" nation="POL" athleteid="3861">
              <RESULTS>
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="3862" heatid="7471" lane="1" entrytime="00:05:31.40" />
                <RESULT eventid="1402" points="48" reactiontime="+114" swimtime="00:02:32.08" resultid="3863" heatid="7594" lane="1" entrytime="00:02:33.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="42" reactiontime="+117" swimtime="00:02:20.76" resultid="3864" heatid="7659" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-15 - brak kontaktu ze ścianą." eventid="1628" reactiontime="+114" status="DSQ" swimtime="00:05:19.18" resultid="3865" heatid="7763" lane="5" entrytime="00:05:06.23" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="3866">
              <RESULTS>
                <RESULT eventid="1075" points="126" reactiontime="+100" swimtime="00:00:40.46" resultid="3867" heatid="7349" lane="3" entrytime="00:00:40.33" />
                <RESULT eventid="1109" points="92" reactiontime="+119" swimtime="00:04:03.49" resultid="3868" heatid="7392" lane="4" entrytime="00:04:11.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.62" />
                    <SPLIT distance="100" swimtime="00:02:04.72" />
                    <SPLIT distance="150" swimtime="00:03:13.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="79" reactiontime="+78" swimtime="00:00:52.69" resultid="3869" heatid="7444" lane="4" entrytime="00:00:51.77" />
                <RESULT eventid="1302" points="92" reactiontime="+122" swimtime="00:01:52.37" resultid="3870" heatid="7540" lane="1" entrytime="00:01:51.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="41" swimtime="00:01:02.86" resultid="3871" heatid="7624" lane="5" entrytime="00:00:58.73" />
                <RESULT eventid="1504" points="102" reactiontime="+127" swimtime="00:03:32.24" resultid="3872" heatid="7688" lane="3" entrytime="00:03:34.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.74" />
                    <SPLIT distance="100" swimtime="00:01:40.70" />
                    <SPLIT distance="150" swimtime="00:02:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="93" reactiontime="+128" swimtime="00:00:55.70" resultid="3873" heatid="7791" lane="1" entrytime="00:00:53.83" />
                <RESULT eventid="1710" points="98" reactiontime="+120" swimtime="00:07:41.24" resultid="3874" heatid="8045" lane="4" entrytime="00:07:26.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.41" />
                    <SPLIT distance="100" swimtime="00:01:48.58" />
                    <SPLIT distance="150" swimtime="00:02:47.70" />
                    <SPLIT distance="200" swimtime="00:03:46.73" />
                    <SPLIT distance="250" swimtime="00:04:46.42" />
                    <SPLIT distance="300" swimtime="00:05:44.17" />
                    <SPLIT distance="350" swimtime="00:06:44.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-22" firstname="Mateusz" gender="M" lastname="Dybek" nation="POL" athleteid="3875">
              <RESULTS>
                <RESULT eventid="1075" points="454" reactiontime="+81" swimtime="00:00:26.40" resultid="3876" heatid="7377" lane="6" entrytime="00:00:26.40" />
                <RESULT eventid="1109" points="393" reactiontime="+89" swimtime="00:02:30.28" resultid="3877" heatid="7401" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:12.12" />
                    <SPLIT distance="150" swimtime="00:01:55.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="490" reactiontime="+69" swimtime="00:00:56.99" resultid="3878" heatid="7522" lane="4" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="403" reactiontime="+85" swimtime="00:02:14.42" resultid="3879" heatid="7703" lane="1" entrytime="00:02:12.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:04.01" />
                    <SPLIT distance="150" swimtime="00:01:39.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-19" firstname="Paulina" gender="F" lastname="Palka" nation="POL" athleteid="3880">
              <RESULTS>
                <RESULT eventid="1183" points="415" reactiontime="+59" swimtime="00:00:34.43" resultid="3881" heatid="7441" lane="6" entrytime="00:00:33.79" />
                <RESULT eventid="1453" points="418" reactiontime="+62" swimtime="00:01:13.85" resultid="3882" heatid="7658" lane="1" entrytime="00:01:12.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="3883" heatid="7761" lane="1" entrytime="00:02:40.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-28" firstname="Wojciech" gender="M" lastname="Wolski" nation="POL" athleteid="3884">
              <RESULTS>
                <RESULT eventid="1075" points="253" reactiontime="+96" swimtime="00:00:32.09" resultid="3885" heatid="7347" lane="2" entrytime="00:03:05.47" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="3886" heatid="7477" lane="5" entrytime="00:03:14.79" />
                <RESULT eventid="1336" points="157" reactiontime="+101" swimtime="00:03:22.20" resultid="3887" heatid="7567" lane="3" entrytime="00:03:16.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:01:30.39" />
                    <SPLIT distance="150" swimtime="00:02:26.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="231" reactiontime="+93" swimtime="00:00:35.48" resultid="3888" heatid="7629" lane="2" entrytime="00:00:36.09" />
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="3889" heatid="7974" lane="4" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="3890" heatid="7741" lane="4" entrytime="00:01:25.72" />
                <RESULT eventid="1662" points="277" reactiontime="+91" swimtime="00:00:38.71" resultid="3891" heatid="7800" lane="3" entrytime="00:00:38.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="3892">
              <RESULTS>
                <RESULT eventid="1183" points="114" swimtime="00:00:52.99" resultid="3893" heatid="7433" lane="5" entrytime="00:00:53.71" />
                <RESULT eventid="1217" points="122" reactiontime="+122" swimtime="00:04:30.79" resultid="3894" heatid="7463" lane="3" entrytime="00:04:29.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.24" />
                    <SPLIT distance="100" swimtime="00:02:10.91" />
                    <SPLIT distance="150" swimtime="00:03:21.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="119" reactiontime="+124" swimtime="00:02:07.17" resultid="3895" heatid="7583" lane="6" entrytime="00:02:10.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="100" swimtime="00:01:58.63" resultid="3896" heatid="7650" lane="5" entrytime="00:01:57.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="109" reactiontime="+83" swimtime="00:04:11.22" resultid="3897" heatid="7755" lane="3" entrytime="00:04:08.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.09" />
                    <SPLIT distance="100" swimtime="00:02:00.76" />
                    <SPLIT distance="150" swimtime="00:03:06.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="114" swimtime="00:00:59.31" resultid="3898" heatid="7777" lane="5" entrytime="00:00:58.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-16" firstname="Tomasz" gender="M" lastname="Doniec" nation="POL" athleteid="3899">
              <RESULTS>
                <RESULT eventid="1109" reactiontime="+112" status="DNS" swimtime="00:00:00.00" resultid="3900" heatid="7391" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                    <SPLIT distance="100" swimtime="00:01:55.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="3901" heatid="7474" lane="3" entrytime="00:03:35.73" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="3902" heatid="7538" lane="4" />
                <RESULT eventid="1402" points="228" reactiontime="+102" swimtime="00:01:30.98" resultid="3903" heatid="7599" lane="2" entrytime="00:01:30.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="3904" heatid="7974" lane="2" />
                <RESULT eventid="1594" reactiontime="+135" status="DNS" swimtime="00:00:00.00" resultid="3905" heatid="7736" lane="2" />
                <RESULT eventid="1662" points="253" reactiontime="+100" swimtime="00:00:39.88" resultid="3906" heatid="7797" lane="3" entrytime="00:00:40.48" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-04" firstname="Małgorzata" gender="F" lastname="Skalska" nation="POL" athleteid="3907">
              <RESULTS>
                <RESULT eventid="1058" points="202" reactiontime="+88" swimtime="00:00:39.57" resultid="3908" heatid="7335" lane="1" entrytime="00:00:40.03" />
                <RESULT eventid="1183" points="137" reactiontime="+68" swimtime="00:00:49.78" resultid="3909" heatid="7433" lane="2" entrytime="00:00:52.03" />
                <RESULT eventid="1217" points="242" swimtime="00:03:35.74" resultid="3910" heatid="7465" lane="5" entrytime="00:03:50.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                    <SPLIT distance="100" swimtime="00:01:46.63" />
                    <SPLIT distance="150" swimtime="00:02:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="254" swimtime="00:01:38.90" resultid="3911" heatid="7586" lane="5" entrytime="00:01:43.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="121" reactiontime="+72" swimtime="00:01:51.36" resultid="3912" heatid="7648" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="234" reactiontime="+79" swimtime="00:00:46.72" resultid="3913" heatid="7781" lane="1" entrytime="00:00:48.05" />
                <RESULT eventid="1693" points="179" reactiontime="+83" swimtime="00:06:56.31" resultid="3914" heatid="8018" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.56" />
                    <SPLIT distance="100" swimtime="00:01:39.90" />
                    <SPLIT distance="150" swimtime="00:02:33.27" />
                    <SPLIT distance="200" swimtime="00:03:26.90" />
                    <SPLIT distance="250" swimtime="00:04:20.31" />
                    <SPLIT distance="300" swimtime="00:05:14.44" />
                    <SPLIT distance="350" swimtime="00:06:07.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-10-29" firstname="Ewa" gender="F" lastname="Macierzewska" nation="POL" athleteid="3915">
              <RESULTS>
                <RESULT eventid="1058" points="22" reactiontime="+168" swimtime="00:01:21.84" resultid="3916" heatid="7332" lane="4" entrytime="00:01:15.75" />
                <RESULT eventid="1183" points="36" reactiontime="+120" swimtime="00:01:17.66" resultid="3917" heatid="7432" lane="2" entrytime="00:01:17.10" />
                <RESULT eventid="1251" points="27" swimtime="00:02:50.00" resultid="3918" heatid="7486" lane="3" entrytime="00:02:44.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="40" reactiontime="+141" swimtime="00:03:03.00" resultid="3919" heatid="7582" lane="1" entrytime="00:02:55.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="35" reactiontime="+90" swimtime="00:02:47.96" resultid="3920" heatid="7649" lane="1" entrytime="00:02:44.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="45" reactiontime="+143" swimtime="00:01:20.96" resultid="3921" heatid="7776" lane="1" entrytime="00:01:17.39" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-10" firstname="Dariusz" gender="M" lastname="Wesołowski" nation="POL" athleteid="3922">
              <RESULTS>
                <RESULT eventid="1268" points="295" reactiontime="+91" swimtime="00:01:07.50" resultid="3923" heatid="7512" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="242" reactiontime="+89" swimtime="00:02:39.42" resultid="3924" heatid="7696" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:15.35" />
                    <SPLIT distance="150" swimtime="00:01:58.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="3925" heatid="8050" lane="4" entrytime="00:05:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-02-11" firstname="Agnieszka" gender="F" lastname="Figuła" nation="POL" athleteid="3926">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="3927" heatid="7342" lane="2" entrytime="00:00:31.02" />
                <RESULT eventid="1251" points="409" reactiontime="+79" swimtime="00:01:08.69" resultid="3928" heatid="7496" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="410" reactiontime="+83" swimtime="00:01:17.71" resultid="3929" heatid="7535" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="416" reactiontime="+80" swimtime="00:01:23.93" resultid="3930" heatid="7590" lane="3" entrytime="00:01:25.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="350" reactiontime="+76" swimtime="00:00:34.59" resultid="3931" heatid="7619" lane="2" entrytime="00:00:34.04" />
                <RESULT eventid="1645" points="416" reactiontime="+77" swimtime="00:00:38.55" resultid="3932" heatid="7786" lane="2" entrytime="00:00:39.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-25" firstname="Jerzy" gender="M" lastname="Korba" nation="POL" athleteid="3933">
              <RESULTS>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1075" status="DSQ" swimtime="00:00:28.10" resultid="3934" heatid="7370" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1109" points="296" reactiontime="+91" swimtime="00:02:45.02" resultid="3935" heatid="7400" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:17.85" />
                    <SPLIT distance="150" swimtime="00:02:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="385" reactiontime="+89" swimtime="00:01:01.76" resultid="3936" heatid="7517" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="301" reactiontime="+75" swimtime="00:00:32.50" resultid="3937" heatid="7635" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1504" points="342" reactiontime="+87" swimtime="00:02:22.03" resultid="3938" heatid="7701" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:09.19" />
                    <SPLIT distance="150" swimtime="00:01:46.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="YMCA Kraków" nation="POL" region="MAL">
          <CONTACT city="Kraków" email="jackwi@poczta.onet.pl" name="Kwiatkowski Jacek" phone="601648456" street="Łuzycka" zip="30658" />
          <ATHLETES>
            <ATHLETE birthdate="1957-03-25" firstname="Jacek" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="3940">
              <RESULTS>
                <RESULT eventid="1075" points="230" reactiontime="+84" swimtime="00:00:33.11" resultid="3941" heatid="7359" lane="2" entrytime="00:00:31.58" entrycourse="SCM" />
                <RESULT eventid="1165" points="201" reactiontime="+97" swimtime="00:24:09.01" resultid="3942" heatid="7910" lane="3" entrytime="00:24:47.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:26.21" />
                    <SPLIT distance="150" swimtime="00:02:14.31" />
                    <SPLIT distance="200" swimtime="00:03:02.84" />
                    <SPLIT distance="250" swimtime="00:03:51.49" />
                    <SPLIT distance="300" swimtime="00:04:40.17" />
                    <SPLIT distance="350" swimtime="00:05:28.98" />
                    <SPLIT distance="400" swimtime="00:06:17.34" />
                    <SPLIT distance="450" swimtime="00:07:06.42" />
                    <SPLIT distance="500" swimtime="00:07:55.10" />
                    <SPLIT distance="550" swimtime="00:08:43.87" />
                    <SPLIT distance="600" swimtime="00:09:32.67" />
                    <SPLIT distance="650" swimtime="00:10:21.45" />
                    <SPLIT distance="700" swimtime="00:11:10.31" />
                    <SPLIT distance="750" swimtime="00:11:59.05" />
                    <SPLIT distance="800" swimtime="00:12:48.07" />
                    <SPLIT distance="850" swimtime="00:13:36.66" />
                    <SPLIT distance="900" swimtime="00:14:25.12" />
                    <SPLIT distance="950" swimtime="00:15:14.55" />
                    <SPLIT distance="1000" swimtime="00:16:03.15" />
                    <SPLIT distance="1050" swimtime="00:16:51.60" />
                    <SPLIT distance="1100" swimtime="00:17:41.24" />
                    <SPLIT distance="1150" swimtime="00:18:29.64" />
                    <SPLIT distance="1200" swimtime="00:19:18.83" />
                    <SPLIT distance="1250" swimtime="00:20:07.76" />
                    <SPLIT distance="1300" swimtime="00:20:56.81" />
                    <SPLIT distance="1350" swimtime="00:21:45.09" />
                    <SPLIT distance="1400" swimtime="00:22:35.07" />
                    <SPLIT distance="1450" swimtime="00:23:23.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="3943" heatid="7508" lane="3" entrytime="00:01:11.80" entrycourse="SCM" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="3944" heatid="7692" lane="4" entrytime="00:02:45.50" entrycourse="SCM" />
                <RESULT eventid="1710" points="200" reactiontime="+95" swimtime="00:06:03.46" resultid="8072" heatid="8043" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:23.07" />
                    <SPLIT distance="150" swimtime="00:02:09.05" />
                    <SPLIT distance="200" swimtime="00:02:56.25" />
                    <SPLIT distance="250" swimtime="00:03:43.81" />
                    <SPLIT distance="300" swimtime="00:04:31.66" />
                    <SPLIT distance="350" swimtime="00:05:19.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00111" name="UKS &quot;TRÓJKA&quot;  Częstochowa" nation="POL" region="SLA">
          <CONTACT city="Częstochowa" email="trojkaczestochowa@poczta.onet.pl" name="Gawda Jacek" phone="511181791" state="ŚL" street="Schillera 5" zip="42-200" />
          <ATHLETES>
            <ATHLETE birthdate="1991-09-11" firstname="Karolina" gender="F" lastname="Wawrzyńczak" nation="POL" license="100111100007" athleteid="3947">
              <RESULTS>
                <RESULT eventid="1183" points="383" swimtime="00:00:35.38" resultid="3948" heatid="7440" lane="2" entrytime="00:00:34.40" />
                <RESULT eventid="1285" points="379" swimtime="00:01:19.74" resultid="3949" heatid="7535" lane="5" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="366" swimtime="00:00:34.07" resultid="3950" heatid="7619" lane="5" entrytime="00:00:34.10" />
                <RESULT eventid="1453" points="372" reactiontime="+74" swimtime="00:01:16.77" resultid="3951" heatid="7657" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="327" reactiontime="+94" swimtime="00:01:19.87" resultid="3952" heatid="7734" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OMDDZ" name="OSiR MASTERS Dzierżoniów" nation="POL" region="DOL">
          <CONTACT city="Dzierżoniów" email="serhetabat@wp.pl" name="Kuszka Piotr" phone="604-22-66-49" state="DOL" street="os. Błękitne 11a/12" zip="58-200" />
          <ATHLETES>
            <ATHLETE birthdate="1983-05-03" firstname="Krzysztof" gender="M" lastname="Pawlaczek" nation="POL" athleteid="3960">
              <RESULTS>
                <RESULT eventid="1234" points="322" reactiontime="+80" swimtime="00:02:55.93" resultid="3961" heatid="7484" lane="4" entrytime="00:02:35.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                    <SPLIT distance="150" swimtime="00:02:04.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="377" reactiontime="+76" swimtime="00:01:10.22" resultid="3962" heatid="7557" lane="2" entrytime="00:01:06.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="376" reactiontime="+78" swimtime="00:01:16.98" resultid="3963" heatid="7610" lane="6" entrytime="00:01:10.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="392" swimtime="00:00:29.78" resultid="3964" heatid="7643" lane="5" entrytime="00:00:28.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-04-14" firstname="Piotr" gender="M" lastname="Kuszka" nation="POL" athleteid="3965">
              <RESULTS>
                <RESULT eventid="1234" points="207" reactiontime="+86" swimtime="00:03:23.81" resultid="3966" heatid="7476" lane="1" entrytime="00:03:21.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                    <SPLIT distance="100" swimtime="00:01:38.35" />
                    <SPLIT distance="150" swimtime="00:02:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="156" reactiontime="+88" swimtime="00:01:34.11" resultid="3967" heatid="7541" lane="6" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="219" reactiontime="+91" swimtime="00:01:32.19" resultid="3968" heatid="7598" lane="3" entrytime="00:01:32.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="152" swimtime="00:00:40.77" resultid="3969" heatid="7627" lane="5" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02914" name="UKS Victoria Józefów" nation="POL" region="MAZ">
          <CONTACT email="ali90@o2.pl" name="kowalczyk alicja" />
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Jan" gender="M" lastname="Kośmider" nation="POL" athleteid="3971">
              <RESULTS>
                <RESULT eventid="1234" points="317" reactiontime="+70" swimtime="00:02:56.79" resultid="3972" heatid="7482" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:21.51" />
                    <SPLIT distance="150" swimtime="00:02:07.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="362" reactiontime="+64" swimtime="00:01:18.01" resultid="3973" heatid="7607" lane="3" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="378" reactiontime="+77" swimtime="00:00:34.92" resultid="3975" heatid="7810" lane="6" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Ukraine Kharkiv" nation="UKR">
          <ATHLETES>
            <ATHLETE birthdate="1975-01-01" firstname="ANDRIY " gender="M" lastname="KHOMENKO" nation="POL" athleteid="3986">
              <RESULTS>
                <RESULT eventid="1109" points="322" reactiontime="+86" swimtime="00:02:40.57" resultid="3988" heatid="7402" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="150" swimtime="00:02:02.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="3989" heatid="7453" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1302" points="360" reactiontime="+81" swimtime="00:01:11.34" resultid="3990" heatid="7549" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="306" reactiontime="+76" swimtime="00:01:12.55" resultid="3991" heatid="7669" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="365" reactiontime="+84" swimtime="00:02:19.03" resultid="3992" heatid="7699" lane="2" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="150" swimtime="00:01:44.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="290" reactiontime="+81" swimtime="00:02:40.23" resultid="3993" heatid="7770" lane="6" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:17.99" />
                    <SPLIT distance="150" swimtime="00:01:59.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="ANDRIY " gender="M" lastname="ZURGALIDZE" nation="UKR" athleteid="3995">
              <RESULTS>
                <RESULT eventid="1109" points="536" reactiontime="+93" swimtime="00:02:15.46" resultid="3996" heatid="7402" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:05.67" />
                    <SPLIT distance="150" swimtime="00:01:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="555" reactiontime="+93" swimtime="00:02:26.76" resultid="3997" heatid="7484" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:11.12" />
                    <SPLIT distance="150" swimtime="00:01:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="546" reactiontime="+88" swimtime="00:01:02.07" resultid="3998" heatid="7559" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="3999" heatid="7671" lane="3" entrytime="00:01:08.00" />
                <RESULT eventid="1559" points="484" reactiontime="+90" status="EXH" swimtime="00:04:59.74" resultid="4000" heatid="7980" lane="3" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:08.17" />
                    <SPLIT distance="150" swimtime="00:01:48.73" />
                    <SPLIT distance="200" swimtime="00:02:29.10" />
                    <SPLIT distance="250" swimtime="00:03:10.20" />
                    <SPLIT distance="300" swimtime="00:03:51.47" />
                    <SPLIT distance="350" swimtime="00:04:27.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="567" reactiontime="+86" swimtime="00:00:30.50" resultid="4001" heatid="7812" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1402" points="568" swimtime="00:01:07.12" resultid="7959" heatid="7592" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="SERGII " gender="M" lastname="BABKIN" nation="UKR" athleteid="4064">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4065" heatid="7374" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4066" heatid="7404" lane="6" entrytime="00:02:30.00" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="4067" heatid="7457" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="4068" heatid="7520" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="4069" heatid="7672" lane="5" entrytime="00:01:07.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="4070" heatid="7703" lane="6" entrytime="00:02:13.00" />
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="4071" heatid="7772" lane="5" entrytime="00:02:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="UKS ORLIK" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1963-01-01" firstname="Lechosław " gender="M" lastname="Jacyszyn" nation="POL" athleteid="4007">
              <RESULTS>
                <RESULT eventid="1302" points="115" reactiontime="+98" swimtime="00:01:44.09" resultid="4008" heatid="7539" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="126" reactiontime="+100" swimtime="00:01:29.41" resultid="4009" heatid="7502" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="87" reactiontime="+104" swimtime="00:00:49.10" resultid="4010" heatid="7624" lane="6" entrytime="00:01:00.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4011" heatid="7392" lane="2" entrytime="00:04:20.00" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="4012" heatid="7737" lane="2" entrytime="00:02:20.00" />
                <RESULT eventid="1710" points="105" reactiontime="+109" swimtime="00:07:30.12" resultid="4013" heatid="8045" lane="1" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                    <SPLIT distance="100" swimtime="00:01:41.12" />
                    <SPLIT distance="150" swimtime="00:03:37.19" />
                    <SPLIT distance="200" swimtime="00:04:35.77" />
                    <SPLIT distance="250" swimtime="00:05:34.13" />
                    <SPLIT distance="300" swimtime="00:06:32.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04211" name="KS Delfin Gliwice" nation="POL" region="11">
          <CONTACT email="ksdelfin@op,pl" name="Cupiał Jarosław" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Teodozja" gender="F" lastname="Gdula" nation="POL" athleteid="4015">
              <RESULTS>
                <RESULT eventid="1217" points="93" swimtime="00:04:57.01" resultid="4016" heatid="7463" lane="5" entrytime="00:04:44.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.23" />
                    <SPLIT distance="100" swimtime="00:02:27.22" />
                    <SPLIT distance="150" swimtime="00:03:43.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="91" reactiontime="+101" swimtime="00:02:18.99" resultid="4017" heatid="7582" lane="3" entrytime="00:02:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="92" reactiontime="+117" swimtime="00:01:03.69" resultid="4018" heatid="7776" lane="3" entrytime="00:01:00.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-10" firstname="Barbara" gender="F" lastname="Lipowska" nation="POL" athleteid="4019">
              <RESULTS>
                <RESULT eventid="1217" points="89" reactiontime="+93" swimtime="00:05:00.95" resultid="4020" heatid="7462" lane="4" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.63" />
                    <SPLIT distance="100" swimtime="00:02:25.00" />
                    <SPLIT distance="150" swimtime="00:03:44.60" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1251" reactiontime="+76" status="DSQ" swimtime="00:02:02.21" resultid="4021" heatid="7487" lane="1" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-11-23" firstname="Jerzy" gender="M" lastname="Marciniszko" nation="POL" athleteid="4022">
              <RESULTS>
                <RESULT eventid="1075" points="32" reactiontime="+97" swimtime="00:01:03.37" resultid="4023" heatid="7347" lane="4" entrytime="00:01:00.75" entrycourse="SCM" />
                <RESULT eventid="1200" points="34" reactiontime="+92" swimtime="00:01:09.21" resultid="4024" heatid="7443" lane="6" entrytime="00:01:11.20" entrycourse="SCM" />
                <RESULT eventid="1234" points="49" swimtime="00:05:29.33" resultid="4025" heatid="7471" lane="5" entrytime="00:05:23.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.11" />
                    <SPLIT distance="100" swimtime="00:02:43.25" />
                    <SPLIT distance="150" swimtime="00:04:11.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="55" swimtime="00:02:25.47" resultid="4026" heatid="7594" lane="5" entrytime="00:02:24.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="22" reactiontime="+97" swimtime="00:02:52.65" resultid="4027" heatid="7660" lane="4" entrytime="00:02:45.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="4028" heatid="7762" lane="2" entrytime="00:05:54.60" entrycourse="SCM" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="4029" heatid="7790" lane="2" entrytime="00:01:00.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="031/05" name="UTW &quot;Masters&quot; Zgierz" nation="POL" region="LOD">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105200002" athleteid="5423">
              <RESULTS>
                <RESULT eventid="1234" points="230" reactiontime="+87" swimtime="00:03:16.95" resultid="5424" heatid="7473" lane="3" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                    <SPLIT distance="150" swimtime="00:02:26.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="5425" heatid="7541" lane="3" entrytime="00:01:35.00" entrycourse="SCM" />
                <RESULT eventid="1402" points="250" reactiontime="+101" swimtime="00:01:28.18" resultid="5426" heatid="7597" lane="1" entrytime="00:01:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="275" swimtime="00:00:38.79" resultid="5427" heatid="7798" lane="5" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1922-01-04" firstname="Kazimierz" gender="M" lastname="Mrówczyński" nation="POL" license="503105200015" athleteid="5428">
              <RESULTS>
                <RESULT eventid="1075" points="44" reactiontime="+123" swimtime="00:00:57.11" resultid="5429" heatid="7347" lane="3" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="1268" points="32" reactiontime="+111" swimtime="00:02:20.81" resultid="5430" heatid="7501" lane="6" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="31" reactiontime="+109" swimtime="00:05:16.01" resultid="5431" heatid="7687" lane="4" entrytime="00:04:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.23" />
                    <SPLIT distance="100" swimtime="00:02:26.72" />
                    <SPLIT distance="150" swimtime="00:03:51.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1662" points="44" reactiontime="+116" swimtime="00:01:11.29" resultid="5432" heatid="7790" lane="1" entrytime="00:01:16.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105100003" athleteid="5433">
              <RESULTS>
                <RESULT eventid="1058" points="336" swimtime="00:00:33.42" resultid="5434" heatid="7340" lane="5" entrytime="00:00:33.50" entrycourse="SCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1183" points="323" reactiontime="+76" swimtime="00:00:37.42" resultid="5435" heatid="7438" lane="2" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1319" points="211" reactiontime="+92" swimtime="00:03:22.60" resultid="5436" heatid="7562" lane="3" entrytime="00:03:22.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="100" swimtime="00:01:33.97" />
                    <SPLIT distance="150" swimtime="00:02:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="312" reactiontime="+86" swimtime="00:00:35.94" resultid="5437" heatid="7618" lane="1" entrytime="00:00:37.50" entrycourse="SCM" />
                <RESULT eventid="1453" points="284" reactiontime="+75" swimtime="00:01:23.99" resultid="5438" heatid="7653" lane="3" entrytime="00:01:26.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="259" reactiontime="+90" swimtime="00:01:26.34" resultid="5439" heatid="7733" lane="4" entrytime="00:01:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="233" reactiontime="+73" swimtime="00:03:14.81" resultid="5440" heatid="7757" lane="3" entrytime="00:03:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                    <SPLIT distance="100" swimtime="00:01:36.97" />
                    <SPLIT distance="150" swimtime="00:02:28.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-07-18" firstname="Tomasz" gender="M" lastname="Niedzwiedz" nation="POL" license="503105200009" athleteid="5441">
              <RESULTS>
                <RESULT comment="K-1 - Stanie" eventid="1109" reactiontime="+111" status="DSQ" swimtime="00:03:32.05" resultid="5442" heatid="7395" lane="1" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                    <SPLIT distance="100" swimtime="00:01:46.84" />
                    <SPLIT distance="150" swimtime="00:02:44.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="5443" heatid="7542" lane="6" entrytime="00:01:35.00" entrycourse="SCM" />
                <RESULT eventid="1336" points="113" reactiontime="+109" swimtime="00:03:45.54" resultid="5444" heatid="7566" lane="3" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.49" />
                    <SPLIT distance="100" swimtime="00:01:48.02" />
                    <SPLIT distance="150" swimtime="00:02:46.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="5445" heatid="7627" lane="6" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="1559" points="140" reactiontime="+114" swimtime="00:07:32.90" resultid="5446" heatid="7977" lane="6" entrytime="00:07:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.01" />
                    <SPLIT distance="100" swimtime="00:01:49.75" />
                    <SPLIT distance="150" swimtime="00:02:50.67" />
                    <SPLIT distance="200" swimtime="00:03:51.76" />
                    <SPLIT distance="250" swimtime="00:04:52.33" />
                    <SPLIT distance="300" swimtime="00:05:53.46" />
                    <SPLIT distance="350" swimtime="00:06:42.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5447" heatid="7739" lane="4" entrytime="00:01:45.00" entrycourse="SCM" />
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="5448" heatid="7764" lane="5" entrytime="00:04:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105200011" athleteid="5449">
              <RESULTS>
                <RESULT eventid="1075" points="181" reactiontime="+95" swimtime="00:00:35.83" resultid="5450" heatid="7357" lane="1" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1109" points="148" swimtime="00:03:27.73" resultid="5451" heatid="7394" lane="5" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                    <SPLIT distance="100" swimtime="00:01:41.96" />
                    <SPLIT distance="150" swimtime="00:02:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="162" reactiontime="+92" swimtime="00:03:41.00" resultid="5452" heatid="7475" lane="4" entrytime="00:03:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                    <SPLIT distance="100" swimtime="00:01:43.51" />
                    <SPLIT distance="150" swimtime="00:02:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="180" reactiontime="+93" swimtime="00:01:29.82" resultid="5453" heatid="7542" lane="4" entrytime="00:01:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="208" reactiontime="+87" swimtime="00:01:33.79" resultid="5454" heatid="7598" lane="4" entrytime="00:01:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="240" swimtime="00:00:40.61" resultid="5455" heatid="7797" lane="5" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-08" firstname="Ewa" gender="F" lastname="Zimna-Walendzik" nation="POL" license="503105100001" athleteid="5456">
              <RESULTS>
                <RESULT eventid="1251" points="159" reactiontime="+92" swimtime="00:01:34.12" resultid="5457" heatid="7490" lane="6" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="159" reactiontime="+98" swimtime="00:01:46.56" resultid="5458" heatid="7528" lane="6" entrytime="00:01:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="128" swimtime="00:00:48.26" resultid="5459" heatid="7614" lane="5" entrytime="00:00:49.00" entrycourse="SCM" />
                <RESULT eventid="1487" points="137" reactiontime="+99" swimtime="00:03:35.22" resultid="5460" heatid="7677" lane="2" entrytime="00:03:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                    <SPLIT distance="100" swimtime="00:01:41.64" />
                    <SPLIT distance="150" swimtime="00:02:38.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="5461" heatid="7731" lane="4" entrytime="00:01:57.00" entrycourse="SCM" />
                <RESULT eventid="1693" points="137" reactiontime="+90" swimtime="00:07:35.08" resultid="5462" heatid="8019" lane="3" entrytime="00:07:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="100" swimtime="00:01:37.75" />
                    <SPLIT distance="150" swimtime="00:02:34.13" />
                    <SPLIT distance="200" swimtime="00:03:33.42" />
                    <SPLIT distance="250" swimtime="00:04:33.95" />
                    <SPLIT distance="300" swimtime="00:05:35.50" />
                    <SPLIT distance="350" swimtime="00:06:36.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-02-07" firstname="Krzysztof" gender="M" lastname="Wojciechowski" nation="POL" license="503105200008" athleteid="5463">
              <RESULTS>
                <RESULT eventid="1075" points="213" reactiontime="+103" swimtime="00:00:33.94" resultid="5464" heatid="7352" lane="2" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1234" points="200" reactiontime="+99" swimtime="00:03:26.22" resultid="5465" heatid="7474" lane="1" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                    <SPLIT distance="100" swimtime="00:01:37.21" />
                    <SPLIT distance="150" swimtime="00:02:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="224" reactiontime="+105" swimtime="00:01:31.56" resultid="5466" heatid="7598" lane="2" entrytime="00:01:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="239" reactiontime="+94" swimtime="00:00:40.65" resultid="5467" heatid="7797" lane="2" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="53105200" athleteid="5473">
              <RESULTS>
                <RESULT eventid="1075" points="471" swimtime="00:00:26.08" resultid="5474" heatid="7376" lane="5" entrytime="00:00:26.50" entrycourse="SCM" />
                <RESULT eventid="1109" points="345" swimtime="00:02:36.84" resultid="5475" heatid="7402" lane="5" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="150" swimtime="00:01:57.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="396" reactiontime="+74" swimtime="00:00:30.78" resultid="5476" heatid="7455" lane="6" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1302" points="403" reactiontime="+93" swimtime="00:01:08.72" resultid="5477" heatid="7555" lane="4" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="396" reactiontime="+89" swimtime="00:00:29.68" resultid="5478" heatid="7642" lane="4" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="5479" heatid="7704" lane="4" entrytime="00:02:09.00" entrycourse="SCM" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5480" heatid="7750" lane="1" entrytime="00:01:05.00" entrycourse="SCM" />
                <RESULT eventid="1662" points="405" reactiontime="+94" swimtime="00:00:34.12" resultid="5481" heatid="7809" lane="2" entrytime="00:00:34.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" license="503105100004" athleteid="5482">
              <RESULTS>
                <RESULT eventid="1058" points="370" reactiontime="+80" swimtime="00:00:32.37" resultid="5483" heatid="7341" lane="2" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1092" points="326" reactiontime="+78" swimtime="00:03:01.01" resultid="5484" heatid="7387" lane="4" entrytime="00:03:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:28.68" />
                    <SPLIT distance="150" swimtime="00:02:18.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="341" reactiontime="+77" swimtime="00:01:12.99" resultid="5485" heatid="7495" lane="6" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="362" swimtime="00:01:20.99" resultid="5486" heatid="7531" lane="5" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="372" reactiontime="+79" swimtime="00:01:27.11" resultid="5487" heatid="7589" lane="3" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="303" reactiontime="+79" swimtime="00:02:45.40" resultid="5488" heatid="7680" lane="4" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:19.47" />
                    <SPLIT distance="150" swimtime="00:02:03.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="393" reactiontime="+78" swimtime="00:00:39.29" resultid="5489" heatid="7786" lane="6" entrytime="00:00:39.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105200001" athleteid="5490">
              <RESULTS>
                <RESULT eventid="1075" points="223" swimtime="00:00:33.47" resultid="5491" heatid="7353" lane="5" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1109" points="129" reactiontime="+102" swimtime="00:03:37.84" resultid="5492" heatid="7393" lane="6" entrytime="00:04:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.98" />
                    <SPLIT distance="100" swimtime="00:01:49.00" />
                    <SPLIT distance="150" swimtime="00:02:55.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="197" reactiontime="+98" swimtime="00:01:17.17" resultid="5493" heatid="7505" lane="3" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="78" reactiontime="+115" swimtime="00:04:14.84" resultid="5494" heatid="7565" lane="3" entrytime="00:04:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.49" />
                    <SPLIT distance="100" swimtime="00:02:05.40" />
                    <SPLIT distance="150" swimtime="00:03:14.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="177" swimtime="00:00:38.77" resultid="5495" heatid="7628" lane="5" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5496" heatid="7739" lane="1" entrytime="00:01:47.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-11-08" firstname="Piotr" gender="M" lastname="Kapczyński" nation="POL" license="503105200017" athleteid="5497">
              <RESULTS>
                <RESULT eventid="1234" points="296" reactiontime="+89" swimtime="00:03:01.04" resultid="5498" heatid="7479" lane="1" entrytime="00:03:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                    <SPLIT distance="100" swimtime="00:01:25.47" />
                    <SPLIT distance="150" swimtime="00:02:14.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="326" reactiontime="+98" swimtime="00:01:20.75" resultid="5499" heatid="7605" lane="2" entrytime="00:01:21.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="340" reactiontime="+101" swimtime="00:00:36.17" resultid="5500" heatid="7809" lane="3" entrytime="00:00:34.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105100006" athleteid="5501">
              <RESULTS>
                <RESULT eventid="1058" points="486" reactiontime="+91" swimtime="00:00:29.57" resultid="5502" heatid="7343" lane="1" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1092" points="445" reactiontime="+91" swimtime="00:02:43.13" resultid="5503" heatid="7389" lane="4" entrytime="00:02:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:02:02.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="437" reactiontime="+67" swimtime="00:00:33.86" resultid="5504" heatid="7440" lane="3" entrytime="00:00:33.90" entrycourse="SCM" />
                <RESULT eventid="1285" points="483" swimtime="00:01:13.56" resultid="5505" heatid="7537" lane="1" entrytime="00:01:13.00" entrycourse="SCM" />
                <RESULT eventid="1453" points="422" reactiontime="+68" swimtime="00:01:13.58" resultid="5506" heatid="7657" lane="2" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="408" reactiontime="+72" swimtime="00:02:41.77" resultid="5507" heatid="7760" lane="3" entrytime="00:02:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:01:58.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105100005" athleteid="5508">
              <RESULTS>
                <RESULT eventid="1092" points="484" reactiontime="+92" swimtime="00:02:38.67" resultid="5509" heatid="7389" lane="1" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:14.37" />
                    <SPLIT distance="150" swimtime="00:02:00.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="386" reactiontime="+73" swimtime="00:00:35.28" resultid="5510" heatid="7440" lane="1" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1285" points="499" reactiontime="+91" swimtime="00:01:12.75" resultid="5511" heatid="7536" lane="3" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="442" reactiontime="+90" swimtime="00:00:32.00" resultid="5512" heatid="7620" lane="2" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1577" points="477" reactiontime="+78" swimtime="00:01:10.45" resultid="5513" heatid="7735" lane="4" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-09-03" firstname="Arkadiusz" gender="M" lastname="Bilski" nation="POL" license="503105200013" athleteid="5514">
              <RESULTS>
                <RESULT eventid="1075" points="394" reactiontime="+79" swimtime="00:00:27.67" resultid="5515" heatid="7353" lane="1" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1234" points="371" reactiontime="+80" swimtime="00:02:47.86" resultid="5516" heatid="7476" lane="3" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:19.73" />
                    <SPLIT distance="150" swimtime="00:02:03.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="5517" heatid="7548" lane="6" entrytime="00:01:17.00" entrycourse="SCM" />
                <RESULT eventid="1402" points="412" reactiontime="+78" swimtime="00:01:14.72" resultid="5518" heatid="7600" lane="3" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="5519" heatid="7633" lane="5" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1662" points="421" reactiontime="+76" swimtime="00:00:33.67" resultid="5520" heatid="7794" lane="6" entrytime="00:00:45.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-23" firstname="Tomasz" gender="M" lastname="Cajdler" nation="POL" license="503105200007" athleteid="5521">
              <RESULTS>
                <RESULT eventid="1075" points="256" reactiontime="+88" swimtime="00:00:31.97" resultid="5522" heatid="7359" lane="3" entrytime="00:00:31.50" entrycourse="SCM" />
                <RESULT eventid="1268" points="232" swimtime="00:01:13.06" resultid="5523" heatid="7508" lane="5" entrytime="00:01:12.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="133" reactiontime="+98" swimtime="00:00:42.70" resultid="5524" heatid="7627" lane="4" entrytime="00:00:38.50" entrycourse="SCM" />
                <RESULT eventid="1662" points="178" reactiontime="+97" swimtime="00:00:44.83" resultid="5525" heatid="7797" lane="6" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-03" firstname="Agata" gender="F" lastname="Głowacka" nation="POL" license="503105100007" athleteid="5526">
              <RESULTS>
                <RESULT eventid="1058" points="269" reactiontime="+104" swimtime="00:00:35.99" resultid="5527" heatid="7337" lane="1" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1183" points="221" reactiontime="+85" swimtime="00:00:42.45" resultid="5528" heatid="7436" lane="3" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1251" points="214" reactiontime="+101" swimtime="00:01:25.15" resultid="5529" heatid="7490" lane="1" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" status="DNS" swimtime="00:00:00.00" resultid="5530" heatid="7530" lane="1" entrytime="00:01:30.00" entrycourse="SCM" />
                <RESULT eventid="1419" points="153" reactiontime="+109" swimtime="00:00:45.56" resultid="5531" heatid="7616" lane="1" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105200006" athleteid="5532">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5533" heatid="7363" lane="1" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1109" points="266" swimtime="00:02:51.16" resultid="5534" heatid="7398" lane="5" entrytime="00:02:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:20.14" />
                    <SPLIT distance="150" swimtime="00:02:12.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="5535" heatid="7514" lane="1" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="231" reactiontime="+82" swimtime="00:02:57.78" resultid="5536" heatid="7569" lane="6" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                    <SPLIT distance="100" swimtime="00:01:24.52" />
                    <SPLIT distance="150" swimtime="00:02:11.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="213" reactiontime="+74" swimtime="00:01:21.91" resultid="5537" heatid="7666" lane="1" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="243" reactiontime="+72" swimtime="00:06:17.11" resultid="5538" heatid="7978" lane="3" entrytime="00:06:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:27.13" />
                    <SPLIT distance="150" swimtime="00:02:16.00" />
                    <SPLIT distance="200" swimtime="00:03:03.23" />
                    <SPLIT distance="250" swimtime="00:04:00.91" />
                    <SPLIT distance="300" swimtime="00:04:58.72" />
                    <SPLIT distance="350" swimtime="00:05:39.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5539" heatid="7744" lane="2" entrytime="00:01:17.00" entrycourse="SCM" />
                <RESULT eventid="1628" reactiontime="+79" status="DNS" swimtime="00:00:00.00" resultid="5540" heatid="7767" lane="1" entrytime="00:02:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-20" firstname="Bogdan" gender="M" lastname="Wąsik" nation="POL" athleteid="7058">
              <RESULTS>
                <RESULT eventid="1234" points="222" reactiontime="+97" swimtime="00:03:19.19" resultid="7059" heatid="7477" lane="2" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.37" />
                    <SPLIT distance="100" swimtime="00:01:35.94" />
                    <SPLIT distance="150" swimtime="00:02:26.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="213" swimtime="00:01:32.98" resultid="7060" heatid="7601" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="7061" heatid="7799" lane="3" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="327" reactiontime="+73" swimtime="00:02:13.21" resultid="5547" heatid="7932" lane="6" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:06.70" />
                    <SPLIT distance="150" swimtime="00:01:38.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5473" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="5497" number="2" reactiontime="+3" />
                    <RELAYPOSITION athleteid="5532" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5463" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="310" swimtime="00:01:59.30" resultid="5548" heatid="7713" lane="5" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                    <SPLIT distance="100" swimtime="00:00:54.47" />
                    <SPLIT distance="150" swimtime="00:01:28.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5473" number="1" />
                    <RELAYPOSITION athleteid="5497" number="2" />
                    <RELAYPOSITION athleteid="5463" number="3" />
                    <RELAYPOSITION athleteid="5532" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1377" points="182" reactiontime="+70" swimtime="00:02:41.77" resultid="5549" heatid="7930" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:26.19" />
                    <SPLIT distance="150" swimtime="00:02:13.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5449" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="5423" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5490" number="3" reactiontime="+87" />
                    <RELAYPOSITION athleteid="5521" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="194" swimtime="00:02:19.46" resultid="5550" heatid="7711" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:48.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5449" number="1" />
                    <RELAYPOSITION athleteid="5423" number="2" />
                    <RELAYPOSITION athleteid="5490" number="3" />
                    <RELAYPOSITION athleteid="5521" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1370" points="392" reactiontime="+70" swimtime="00:02:20.21" resultid="5545" heatid="7573" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:13.94" />
                    <SPLIT distance="150" swimtime="00:01:46.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5501" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="5482" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5508" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5433" number="4" reactiontime="+73" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1521" points="398" reactiontime="+88" swimtime="00:02:06.75" resultid="5546" heatid="7708" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="150" swimtime="00:01:37.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5508" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="5433" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="5482" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5501" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1126" points="332" reactiontime="+80" swimtime="00:01:56.64" resultid="5541" heatid="7411" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="150" swimtime="00:01:30.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5514" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5433" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="5501" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5473" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" points="347" reactiontime="+71" swimtime="00:02:10.58" resultid="5542" heatid="7819" lane="5" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="100" swimtime="00:01:07.60" />
                    <SPLIT distance="150" swimtime="00:01:37.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5501" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5514" number="2" />
                    <RELAYPOSITION athleteid="5473" number="3" />
                    <RELAYPOSITION athleteid="5433" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1126" points="285" reactiontime="+93" swimtime="00:02:02.70" resultid="5543" heatid="7411" lane="6" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:01.49" />
                    <SPLIT distance="150" swimtime="00:01:32.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5497" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="5482" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="5508" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="5532" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" points="298" reactiontime="+71" swimtime="00:02:17.40" resultid="5544" heatid="7818" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:45.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5532" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5497" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="5508" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5482" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1679" points="154" reactiontime="+83" swimtime="00:02:51.01" resultid="5551" heatid="7815" lane="6" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:22.86" />
                    <SPLIT distance="150" swimtime="00:02:09.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5526" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="5463" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5490" number="3" reactiontime="+98" />
                    <RELAYPOSITION athleteid="5456" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MKS AQUATI" name="Mks Aquatic Gubin" nation="POL">
          <CONTACT city="Gubin" email="mks@gubin.com.pl" name="Patek Ziemowit" phone="693323270" state="LUBUS" street="Świerczewskiego 20/4" zip="66-620" />
          <ATHLETES>
            <ATHLETE birthdate="1953-05-24" firstname="Anna" gender="F" lastname="Krupińska" nation="POL" athleteid="4036">
              <RESULTS>
                <RESULT eventid="1217" points="186" reactiontime="+118" swimtime="00:03:55.60" resultid="4037" heatid="7465" lane="6" entrytime="00:03:57.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.35" />
                    <SPLIT distance="100" swimtime="00:01:53.63" />
                    <SPLIT distance="150" swimtime="00:02:54.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="191" reactiontime="+112" swimtime="00:01:48.78" resultid="4038" heatid="7585" lane="1" entrytime="00:01:50.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="203" reactiontime="+109" swimtime="00:00:48.96" resultid="4039" heatid="7779" lane="4" entrytime="00:00:50.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-29" firstname="Sylwia" gender="F" lastname="Gorockiewicz" nation="POL" athleteid="4040">
              <RESULTS>
                <RESULT eventid="1385" points="92" reactiontime="+119" swimtime="00:02:18.48" resultid="4041" heatid="7582" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="92" reactiontime="+111" swimtime="00:01:03.69" resultid="4042" heatid="7777" lane="6" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="UKS G-8 Warszawa" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Krzysztof " gender="M" lastname="Wiater" nation="POL" athleteid="4053" />
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Victory Masters Elbląg" nation="POL">
          <CONTACT city="Elbląg" name="Latecki Grzegorz" street="Łokietka 45" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1966-06-06" firstname="Andrzej" gender="M" lastname="Pasieczny" nation="POL" athleteid="4074">
              <RESULTS>
                <RESULT eventid="1075" points="381" reactiontime="+86" swimtime="00:00:28.00" resultid="4075" heatid="7369" lane="1" entrytime="00:00:28.22" />
                <RESULT eventid="1336" points="434" reactiontime="+90" swimtime="00:02:24.05" resultid="4076" heatid="7571" lane="2" entrytime="00:02:23.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:07.37" />
                    <SPLIT distance="150" swimtime="00:01:44.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="455" reactiontime="+87" swimtime="00:02:09.17" resultid="4077" heatid="7704" lane="2" entrytime="00:02:09.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="100" swimtime="00:01:02.46" />
                    <SPLIT distance="150" swimtime="00:01:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="419" reactiontime="+89" swimtime="00:01:04.78" resultid="4078" heatid="7751" lane="6" entrytime="00:01:03.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1710" points="453" reactiontime="+88" swimtime="00:04:37.02" resultid="4079" heatid="8055" lane="3" entrytime="00:04:45.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:05.90" />
                    <SPLIT distance="150" swimtime="00:01:40.39" />
                    <SPLIT distance="200" swimtime="00:02:15.39" />
                    <SPLIT distance="250" swimtime="00:02:50.53" />
                    <SPLIT distance="300" swimtime="00:03:26.24" />
                    <SPLIT distance="350" swimtime="00:04:01.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-05" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="4080">
              <RESULTS>
                <RESULT comment="Przekroczony limit czasu. (14:00.00)" eventid="1148" reactiontime="+110" status="DSQ" swimtime="00:14:38.50" resultid="4081" heatid="7903" lane="4" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.06" />
                    <SPLIT distance="100" swimtime="00:01:47.26" />
                    <SPLIT distance="150" swimtime="00:02:43.66" />
                    <SPLIT distance="200" swimtime="00:03:39.61" />
                    <SPLIT distance="250" swimtime="00:04:35.94" />
                    <SPLIT distance="300" swimtime="00:05:31.96" />
                    <SPLIT distance="350" swimtime="00:06:27.71" />
                    <SPLIT distance="400" swimtime="00:07:23.11" />
                    <SPLIT distance="450" swimtime="00:08:18.79" />
                    <SPLIT distance="500" swimtime="00:09:14.56" />
                    <SPLIT distance="550" swimtime="00:10:09.21" />
                    <SPLIT distance="600" swimtime="00:11:03.53" />
                    <SPLIT distance="650" swimtime="00:11:58.06" />
                    <SPLIT distance="700" swimtime="00:12:52.58" />
                    <SPLIT distance="750" swimtime="00:13:47.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="151" reactiontime="+101" swimtime="00:01:35.72" resultid="4082" heatid="7489" lane="1" entrytime="00:01:36.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="145" reactiontime="+105" swimtime="00:03:31.22" resultid="4083" heatid="7676" lane="3" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.60" />
                    <SPLIT distance="100" swimtime="00:01:44.96" />
                    <SPLIT distance="150" swimtime="00:02:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="155" swimtime="00:07:16.68" resultid="4084" heatid="8020" lane="5" entrytime="00:07:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.54" />
                    <SPLIT distance="100" swimtime="00:01:45.00" />
                    <SPLIT distance="150" swimtime="00:02:40.15" />
                    <SPLIT distance="200" swimtime="00:03:35.85" />
                    <SPLIT distance="250" swimtime="00:04:32.62" />
                    <SPLIT distance="300" swimtime="00:05:29.51" />
                    <SPLIT distance="350" swimtime="00:06:24.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karaś" nation="POL" athleteid="4085">
              <RESULTS>
                <RESULT eventid="1148" points="172" swimtime="00:14:30.47" resultid="4086" heatid="7903" lane="5" entrytime="00:14:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                    <SPLIT distance="100" swimtime="00:01:43.83" />
                    <SPLIT distance="150" swimtime="00:02:37.65" />
                    <SPLIT distance="200" swimtime="00:03:31.69" />
                    <SPLIT distance="250" swimtime="00:04:26.35" />
                    <SPLIT distance="300" swimtime="00:05:21.18" />
                    <SPLIT distance="350" swimtime="00:06:16.78" />
                    <SPLIT distance="400" swimtime="00:07:12.31" />
                    <SPLIT distance="450" swimtime="00:08:08.54" />
                    <SPLIT distance="500" swimtime="00:09:04.44" />
                    <SPLIT distance="550" swimtime="00:09:59.69" />
                    <SPLIT distance="600" swimtime="00:10:55.78" />
                    <SPLIT distance="650" swimtime="00:11:50.44" />
                    <SPLIT distance="700" swimtime="00:12:45.77" />
                    <SPLIT distance="750" swimtime="00:13:39.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="121" reactiontime="+118" swimtime="00:04:03.84" resultid="4087" heatid="7562" lane="6" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.93" />
                    <SPLIT distance="100" swimtime="00:01:56.11" />
                    <SPLIT distance="150" swimtime="00:03:00.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="142" reactiontime="+115" swimtime="00:08:19.76" resultid="4088" heatid="7717" lane="6" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.46" />
                    <SPLIT distance="100" swimtime="00:01:56.43" />
                    <SPLIT distance="150" swimtime="00:03:02.47" />
                    <SPLIT distance="200" swimtime="00:04:05.92" />
                    <SPLIT distance="250" swimtime="00:05:19.84" />
                    <SPLIT distance="300" swimtime="00:06:36.89" />
                    <SPLIT distance="350" swimtime="00:07:28.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="115" reactiontime="+106" swimtime="00:01:53.18" resultid="4089" heatid="7732" lane="1" entrytime="00:01:47.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="156" reactiontime="+114" swimtime="00:07:16.15" resultid="4090" heatid="8020" lane="2" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.23" />
                    <SPLIT distance="100" swimtime="00:01:45.53" />
                    <SPLIT distance="150" swimtime="00:02:41.41" />
                    <SPLIT distance="200" swimtime="00:03:37.70" />
                    <SPLIT distance="250" swimtime="00:04:33.36" />
                    <SPLIT distance="300" swimtime="00:05:28.15" />
                    <SPLIT distance="350" swimtime="00:06:24.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-12-08" firstname="Pawł" gender="M" lastname="Stawiarz" nation="POL" athleteid="4091">
              <RESULTS>
                <RESULT eventid="1075" points="374" reactiontime="+92" swimtime="00:00:28.17" resultid="4092" heatid="7368" lane="1" entrytime="00:00:28.50" />
                <RESULT eventid="1268" points="342" reactiontime="+76" swimtime="00:01:04.22" resultid="4093" heatid="7514" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="4094" heatid="7695" lane="3" entrytime="00:02:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-12" firstname="Grzegorz" gender="M" lastname="Latecki" nation="POL" athleteid="4095">
              <RESULTS>
                <RESULT eventid="1200" points="295" reactiontime="+69" swimtime="00:00:33.94" resultid="4096" heatid="7453" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1436" points="351" reactiontime="+84" swimtime="00:00:30.90" resultid="4097" heatid="7638" lane="2" entrytime="00:00:30.50" />
                <RESULT eventid="1470" points="277" reactiontime="+68" swimtime="00:01:15.01" resultid="4098" heatid="7668" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="4100" heatid="7769" lane="2" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-06-10" firstname="Tomasz" gender="M" lastname="Gleb" nation="POL" athleteid="4101">
              <RESULTS>
                <RESULT eventid="1075" points="313" reactiontime="+88" swimtime="00:00:29.89" resultid="4102" heatid="7366" lane="2" entrytime="00:00:29.20" />
                <RESULT eventid="1165" points="297" reactiontime="+93" swimtime="00:21:13.84" resultid="4103" heatid="7914" lane="1" entrytime="00:21:49.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:01:56.66" />
                    <SPLIT distance="200" swimtime="00:02:37.84" />
                    <SPLIT distance="250" swimtime="00:03:19.75" />
                    <SPLIT distance="300" swimtime="00:04:01.43" />
                    <SPLIT distance="350" swimtime="00:04:43.56" />
                    <SPLIT distance="400" swimtime="00:05:25.67" />
                    <SPLIT distance="450" swimtime="00:06:08.21" />
                    <SPLIT distance="500" swimtime="00:06:51.42" />
                    <SPLIT distance="550" swimtime="00:07:34.36" />
                    <SPLIT distance="600" swimtime="00:08:17.28" />
                    <SPLIT distance="650" swimtime="00:09:00.41" />
                    <SPLIT distance="700" swimtime="00:09:43.22" />
                    <SPLIT distance="750" swimtime="00:10:26.70" />
                    <SPLIT distance="800" swimtime="00:11:09.59" />
                    <SPLIT distance="850" swimtime="00:11:52.61" />
                    <SPLIT distance="900" swimtime="00:12:36.47" />
                    <SPLIT distance="950" swimtime="00:13:20.78" />
                    <SPLIT distance="1000" swimtime="00:14:04.63" />
                    <SPLIT distance="1050" swimtime="00:14:48.52" />
                    <SPLIT distance="1100" swimtime="00:15:32.96" />
                    <SPLIT distance="1150" swimtime="00:16:16.86" />
                    <SPLIT distance="1200" swimtime="00:16:59.96" />
                    <SPLIT distance="1250" swimtime="00:17:43.69" />
                    <SPLIT distance="1300" swimtime="00:18:27.24" />
                    <SPLIT distance="1350" swimtime="00:19:09.66" />
                    <SPLIT distance="1400" swimtime="00:19:53.01" />
                    <SPLIT distance="1450" swimtime="00:20:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="273" reactiontime="+98" swimtime="00:03:06.00" resultid="4104" heatid="7478" lane="1" entrytime="00:03:09.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                    <SPLIT distance="100" swimtime="00:01:27.16" />
                    <SPLIT distance="150" swimtime="00:02:16.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="321" swimtime="00:01:05.58" resultid="4105" heatid="7514" lane="5" entrytime="00:01:05.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="4106" heatid="7602" lane="2" entrytime="00:01:25.45" />
                <RESULT eventid="1559" points="214" reactiontime="+96" swimtime="00:06:33.48" resultid="4107" heatid="7979" lane="6" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:26.18" />
                    <SPLIT distance="150" swimtime="00:02:19.30" />
                    <SPLIT distance="200" swimtime="00:03:12.51" />
                    <SPLIT distance="250" swimtime="00:04:09.53" />
                    <SPLIT distance="300" swimtime="00:05:06.81" />
                    <SPLIT distance="350" swimtime="00:05:51.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="308" swimtime="00:05:14.84" resultid="4108" heatid="8053" lane="5" entrytime="00:05:15.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:01:57.45" />
                    <SPLIT distance="200" swimtime="00:02:37.96" />
                    <SPLIT distance="250" swimtime="00:03:18.64" />
                    <SPLIT distance="300" swimtime="00:03:58.33" />
                    <SPLIT distance="350" swimtime="00:04:37.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03801" name="UKS DELFINEK Legnica" nation="POL">
          <CONTACT name="Malchar" phone="506034671" />
          <ATHLETES>
            <ATHLETE birthdate="1982-12-28" firstname="Jowita" gender="F" lastname="Malchar" nation="POL" athleteid="4110">
              <RESULTS>
                <RESULT eventid="1058" points="425" reactiontime="+80" swimtime="00:00:30.90" resultid="4111" heatid="7342" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1092" points="387" reactiontime="+84" swimtime="00:02:50.91" resultid="4112" heatid="7388" lane="1" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:18.93" />
                    <SPLIT distance="150" swimtime="00:02:08.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="352" reactiontime="+83" swimtime="00:03:10.51" resultid="4113" heatid="7468" lane="1" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                    <SPLIT distance="100" swimtime="00:01:31.76" />
                    <SPLIT distance="150" swimtime="00:02:21.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="292" reactiontime="+91" swimtime="00:03:01.95" resultid="4114" heatid="7563" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:25.52" />
                    <SPLIT distance="150" swimtime="00:02:13.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="367" reactiontime="+84" swimtime="00:01:27.57" resultid="4115" heatid="7590" lane="1" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1542" points="373" reactiontime="+97" swimtime="00:06:02.57" resultid="4116" heatid="7718" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:22.18" />
                    <SPLIT distance="150" swimtime="00:02:08.32" />
                    <SPLIT distance="200" swimtime="00:02:54.24" />
                    <SPLIT distance="250" swimtime="00:03:46.05" />
                    <SPLIT distance="300" swimtime="00:04:36.98" />
                    <SPLIT distance="350" swimtime="00:05:20.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="338" swimtime="00:01:18.96" resultid="4117" heatid="7734" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="383" swimtime="00:00:39.65" resultid="4118" heatid="7785" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00308" name="MKP Bobry Dębica" nation="POL" region="PDK">
          <CONTACT name="GOGACZ" phone="506694816" />
          <ATHLETES>
            <ATHLETE birthdate="1981-04-11" firstname="Przemysław" gender="M" lastname="Jurek" nation="POL" athleteid="4120">
              <RESULTS>
                <RESULT eventid="1075" points="540" reactiontime="+80" swimtime="00:00:24.92" resultid="4121" heatid="7378" lane="2" entrytime="00:00:25.89" />
                <RESULT eventid="1165" points="444" reactiontime="+88" swimtime="00:18:33.50" resultid="4122" heatid="7916" lane="2" entrytime="00:18:35.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:42.32" />
                    <SPLIT distance="200" swimtime="00:02:18.34" />
                    <SPLIT distance="250" swimtime="00:02:54.92" />
                    <SPLIT distance="300" swimtime="00:03:31.92" />
                    <SPLIT distance="350" swimtime="00:04:08.91" />
                    <SPLIT distance="400" swimtime="00:04:45.95" />
                    <SPLIT distance="450" swimtime="00:05:23.04" />
                    <SPLIT distance="500" swimtime="00:06:00.22" />
                    <SPLIT distance="550" swimtime="00:06:37.49" />
                    <SPLIT distance="600" swimtime="00:07:14.80" />
                    <SPLIT distance="650" swimtime="00:07:51.96" />
                    <SPLIT distance="700" swimtime="00:08:29.05" />
                    <SPLIT distance="750" swimtime="00:09:06.09" />
                    <SPLIT distance="800" swimtime="00:09:43.15" />
                    <SPLIT distance="850" swimtime="00:10:20.30" />
                    <SPLIT distance="900" swimtime="00:10:57.47" />
                    <SPLIT distance="950" swimtime="00:11:35.30" />
                    <SPLIT distance="1000" swimtime="00:12:13.05" />
                    <SPLIT distance="1050" swimtime="00:12:50.38" />
                    <SPLIT distance="1100" swimtime="00:13:28.02" />
                    <SPLIT distance="1150" swimtime="00:14:05.86" />
                    <SPLIT distance="1200" swimtime="00:14:43.75" />
                    <SPLIT distance="1250" swimtime="00:15:22.39" />
                    <SPLIT distance="1300" swimtime="00:16:00.57" />
                    <SPLIT distance="1350" swimtime="00:16:38.84" />
                    <SPLIT distance="1400" swimtime="00:17:17.45" />
                    <SPLIT distance="1450" swimtime="00:17:56.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="508" swimtime="00:01:03.58" resultid="4123" heatid="7557" lane="5" entrytime="00:01:06.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="509" reactiontime="+85" swimtime="00:00:27.30" resultid="4124" heatid="7645" lane="3" entrytime="00:00:27.03" />
                <RESULT eventid="1594" points="473" reactiontime="+90" swimtime="00:01:02.21" resultid="4125" heatid="7751" lane="2" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="484" reactiontime="+92" swimtime="00:04:30.95" resultid="4126" heatid="8057" lane="6" entrytime="00:04:42.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                    <SPLIT distance="100" swimtime="00:01:03.08" />
                    <SPLIT distance="150" swimtime="00:01:37.44" />
                    <SPLIT distance="200" swimtime="00:02:12.19" />
                    <SPLIT distance="250" swimtime="00:02:46.65" />
                    <SPLIT distance="300" swimtime="00:03:21.51" />
                    <SPLIT distance="350" swimtime="00:03:56.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-23" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" athleteid="4127">
              <RESULTS>
                <RESULT eventid="1148" points="372" reactiontime="+92" swimtime="00:11:13.30" resultid="4128" heatid="7906" lane="6" entrytime="00:10:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:15.18" />
                    <SPLIT distance="150" swimtime="00:01:55.68" />
                    <SPLIT distance="200" swimtime="00:02:36.73" />
                    <SPLIT distance="250" swimtime="00:03:18.63" />
                    <SPLIT distance="300" swimtime="00:04:01.18" />
                    <SPLIT distance="350" swimtime="00:04:43.90" />
                    <SPLIT distance="400" swimtime="00:05:26.68" />
                    <SPLIT distance="450" swimtime="00:06:09.43" />
                    <SPLIT distance="500" swimtime="00:06:52.24" />
                    <SPLIT distance="550" swimtime="00:07:35.32" />
                    <SPLIT distance="600" swimtime="00:08:18.71" />
                    <SPLIT distance="650" swimtime="00:09:02.62" />
                    <SPLIT distance="700" swimtime="00:09:46.81" />
                    <SPLIT distance="750" swimtime="00:10:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="431" reactiontime="+66" swimtime="00:00:34.01" resultid="4129" heatid="7440" lane="5" entrytime="00:00:34.90" />
                <RESULT eventid="1285" points="417" reactiontime="+93" swimtime="00:01:17.27" resultid="4130" heatid="7535" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="429" reactiontime="+68" swimtime="00:01:13.22" resultid="4131" heatid="7657" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="433" reactiontime="+72" swimtime="00:02:38.55" resultid="4132" heatid="7761" lane="6" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:16.77" />
                    <SPLIT distance="150" swimtime="00:01:57.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-27" firstname="Miłosz" gender="M" lastname="Pagacz" nation="POL" athleteid="4133">
              <RESULTS>
                <RESULT eventid="1075" points="213" reactiontime="+93" swimtime="00:00:33.96" resultid="4134" heatid="7351" lane="3" entrytime="00:00:36.20" />
                <RESULT eventid="1268" points="192" swimtime="00:01:17.82" resultid="4136" heatid="7503" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="182" reactiontime="+95" swimtime="00:02:55.15" resultid="4137" heatid="7691" lane="1" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:19.12" />
                    <SPLIT distance="150" swimtime="00:02:04.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="167" reactiontime="+89" swimtime="00:06:26.11" resultid="4138" heatid="8046" lane="2" entrytime="00:06:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:01:25.62" />
                    <SPLIT distance="150" swimtime="00:02:11.55" />
                    <SPLIT distance="200" swimtime="00:03:01.56" />
                    <SPLIT distance="250" swimtime="00:03:54.48" />
                    <SPLIT distance="300" swimtime="00:04:43.48" />
                    <SPLIT distance="350" swimtime="00:05:34.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-24" firstname="Radosław" gender="M" lastname="Jurek" nation="POL" athleteid="4139">
              <RESULTS>
                <RESULT eventid="1075" points="366" swimtime="00:00:28.36" resultid="4140" heatid="7371" lane="5" entrytime="00:00:27.90" />
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="4141" heatid="7639" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="4142" heatid="7695" lane="2" entrytime="00:02:35.00" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="4143" heatid="7744" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="4144" heatid="8049" lane="4" entrytime="00:05:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-14" firstname="Agnieszka" gender="F" lastname="Opitz" nation="POL" athleteid="4145">
              <RESULTS>
                <RESULT eventid="1217" points="394" swimtime="00:03:03.55" resultid="4146" heatid="7468" lane="5" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:29.88" />
                    <SPLIT distance="150" swimtime="00:02:17.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="424" swimtime="00:01:23.43" resultid="4147" heatid="7589" lane="5" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="427" reactiontime="+77" swimtime="00:00:38.23" resultid="4148" heatid="7787" lane="6" entrytime="00:00:38.21" />
                <RESULT eventid="1693" points="364" reactiontime="+82" swimtime="00:05:28.91" resultid="4149" heatid="8025" lane="6" entrytime="00:05:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:17.07" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                    <SPLIT distance="200" swimtime="00:02:42.19" />
                    <SPLIT distance="250" swimtime="00:03:24.86" />
                    <SPLIT distance="300" swimtime="00:04:07.58" />
                    <SPLIT distance="350" swimtime="00:04:49.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-07-08" firstname="Andrzej" gender="M" lastname="Maciejczak" nation="POL" athleteid="4150">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4151" heatid="7356" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1165" points="153" reactiontime="+108" swimtime="00:26:28.89" resultid="4152" heatid="7910" lane="6" entrytime="00:26:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                    <SPLIT distance="100" swimtime="00:01:29.51" />
                    <SPLIT distance="150" swimtime="00:02:20.39" />
                    <SPLIT distance="200" swimtime="00:03:11.45" />
                    <SPLIT distance="250" swimtime="00:04:03.40" />
                    <SPLIT distance="300" swimtime="00:04:55.45" />
                    <SPLIT distance="350" swimtime="00:05:49.89" />
                    <SPLIT distance="400" swimtime="00:06:42.22" />
                    <SPLIT distance="450" swimtime="00:07:34.74" />
                    <SPLIT distance="500" swimtime="00:08:27.62" />
                    <SPLIT distance="550" swimtime="00:09:20.25" />
                    <SPLIT distance="600" swimtime="00:10:13.35" />
                    <SPLIT distance="650" swimtime="00:11:06.56" />
                    <SPLIT distance="700" swimtime="00:12:00.83" />
                    <SPLIT distance="750" swimtime="00:12:53.96" />
                    <SPLIT distance="800" swimtime="00:13:47.16" />
                    <SPLIT distance="850" swimtime="00:14:40.55" />
                    <SPLIT distance="900" swimtime="00:15:33.66" />
                    <SPLIT distance="950" swimtime="00:16:27.93" />
                    <SPLIT distance="1000" swimtime="00:17:21.15" />
                    <SPLIT distance="1050" swimtime="00:18:15.60" />
                    <SPLIT distance="1100" swimtime="00:19:10.28" />
                    <SPLIT distance="1150" swimtime="00:20:05.17" />
                    <SPLIT distance="1200" swimtime="00:20:59.69" />
                    <SPLIT distance="1250" swimtime="00:21:54.84" />
                    <SPLIT distance="1300" swimtime="00:22:50.12" />
                    <SPLIT distance="1350" swimtime="00:23:44.30" />
                    <SPLIT distance="1400" swimtime="00:24:39.89" />
                    <SPLIT distance="1450" swimtime="00:25:36.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="176" reactiontime="+109" swimtime="00:01:20.07" resultid="4153" heatid="7505" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="172" reactiontime="+109" swimtime="00:06:22.04" resultid="4154" heatid="8047" lane="4" entrytime="00:06:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:02:14.48" />
                    <SPLIT distance="200" swimtime="00:03:04.47" />
                    <SPLIT distance="250" swimtime="00:03:54.52" />
                    <SPLIT distance="300" swimtime="00:04:44.60" />
                    <SPLIT distance="350" swimtime="00:05:34.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4155" heatid="7710" lane="2" />
                <RESULT eventid="1377" status="DNS" swimtime="00:00:00.00" resultid="4156" heatid="7929" lane="1" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1679" points="377" reactiontime="+66" swimtime="00:02:06.98" resultid="5260" heatid="7814" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:12.03" />
                    <SPLIT distance="150" swimtime="00:01:39.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4127" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4145" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="4120" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="4139" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1126" points="360" reactiontime="+94" swimtime="00:01:53.48" resultid="5261" heatid="7408" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:00:59.17" />
                    <SPLIT distance="150" swimtime="00:01:29.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4127" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="4139" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="4145" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4120" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="UKS Energetyk Zgorzelec" nation="POL" region="DOL">
          <CONTACT name="Daszyński" phone="607151541" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="4206">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4207" heatid="7350" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4208" heatid="7393" lane="2" entrytime="00:03:58.65" />
                <RESULT eventid="1234" points="92" swimtime="00:04:26.83" resultid="4209" heatid="7472" lane="5" entrytime="00:04:25.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.34" />
                    <SPLIT distance="100" swimtime="00:02:11.27" />
                    <SPLIT distance="150" swimtime="00:03:21.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="57" reactiontime="+97" swimtime="00:04:43.19" resultid="4210" heatid="7565" lane="1" entrytime="00:04:31.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.45" />
                    <SPLIT distance="100" swimtime="00:02:11.35" />
                    <SPLIT distance="150" swimtime="00:03:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="90" reactiontime="+81" swimtime="00:01:49.02" resultid="4211" heatid="7662" lane="2" entrytime="00:01:47.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="91" reactiontime="+95" swimtime="00:08:41.88" resultid="4212" heatid="7975" lane="3" entrytime="00:08:29.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.43" />
                    <SPLIT distance="100" swimtime="00:02:08.81" />
                    <SPLIT distance="150" swimtime="00:03:13.17" />
                    <SPLIT distance="200" swimtime="00:04:16.63" />
                    <SPLIT distance="250" swimtime="00:05:31.02" />
                    <SPLIT distance="300" swimtime="00:06:41.28" />
                    <SPLIT distance="350" swimtime="00:07:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="54" reactiontime="+108" swimtime="00:02:07.96" resultid="4213" heatid="7738" lane="2" entrytime="00:02:02.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="91" reactiontime="+83" swimtime="00:03:55.84" resultid="4214" heatid="7764" lane="2" entrytime="00:03:52.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.91" />
                    <SPLIT distance="100" swimtime="00:01:56.07" />
                    <SPLIT distance="150" swimtime="00:02:58.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Aquasfera Masters Olsztyn" nation="POL">
          <CONTACT email="gozdzik@uwm.edu.pl" name="Gożdziejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="Piekut" nation="POL" athleteid="4255">
              <RESULTS>
                <RESULT eventid="1092" points="388" reactiontime="+85" swimtime="00:02:50.72" resultid="4256" heatid="7388" lane="4" entrytime="00:02:48.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:18.58" />
                    <SPLIT distance="150" swimtime="00:02:08.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="354" reactiontime="+70" swimtime="00:00:36.31" resultid="4257" heatid="7439" lane="5" entrytime="00:00:36.49" />
                <RESULT eventid="1319" points="419" reactiontime="+88" swimtime="00:02:41.33" resultid="4258" heatid="7563" lane="3" entrytime="00:02:42.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:18.44" />
                    <SPLIT distance="150" swimtime="00:02:00.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="380" reactiontime="+81" swimtime="00:00:33.63" resultid="4259" heatid="7620" lane="1" entrytime="00:00:33.78" />
                <RESULT eventid="1542" points="375" reactiontime="+92" swimtime="00:06:01.86" resultid="4260" heatid="7718" lane="3" entrytime="00:05:27.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="100" swimtime="00:01:20.33" />
                    <SPLIT distance="150" swimtime="00:02:08.54" />
                    <SPLIT distance="200" swimtime="00:02:56.20" />
                    <SPLIT distance="250" swimtime="00:03:48.56" />
                    <SPLIT distance="300" swimtime="00:04:40.18" />
                    <SPLIT distance="350" swimtime="00:05:21.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="362" reactiontime="+88" swimtime="00:01:17.21" resultid="4261" heatid="7735" lane="2" entrytime="00:01:14.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="4262" heatid="7784" lane="2" entrytime="00:00:42.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-12-05" firstname="Aleksandra" gender="F" lastname="Góralska" nation="POL" athleteid="4263">
              <RESULTS>
                <RESULT eventid="1058" points="246" reactiontime="+93" swimtime="00:00:37.10" resultid="4264" heatid="7335" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1148" points="251" reactiontime="+105" swimtime="00:12:47.76" resultid="4265" heatid="7903" lane="2" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:31.11" />
                    <SPLIT distance="150" swimtime="00:02:19.06" />
                    <SPLIT distance="200" swimtime="00:03:07.60" />
                    <SPLIT distance="250" swimtime="00:03:56.81" />
                    <SPLIT distance="300" swimtime="00:04:45.99" />
                    <SPLIT distance="350" swimtime="00:05:34.73" />
                    <SPLIT distance="400" swimtime="00:06:23.17" />
                    <SPLIT distance="450" swimtime="00:07:11.51" />
                    <SPLIT distance="500" swimtime="00:07:59.79" />
                    <SPLIT distance="550" swimtime="00:08:48.46" />
                    <SPLIT distance="600" swimtime="00:09:36.68" />
                    <SPLIT distance="650" swimtime="00:10:26.05" />
                    <SPLIT distance="700" swimtime="00:11:14.60" />
                    <SPLIT distance="750" swimtime="00:12:02.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="253" swimtime="00:06:11.40" resultid="4266" heatid="8021" lane="5" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:01:26.62" />
                    <SPLIT distance="150" swimtime="00:02:13.68" />
                    <SPLIT distance="200" swimtime="00:03:01.28" />
                    <SPLIT distance="250" swimtime="00:03:49.35" />
                    <SPLIT distance="300" swimtime="00:04:37.05" />
                    <SPLIT distance="350" swimtime="00:05:24.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-02" firstname="Piotr" gender="M" lastname="Suchecki" nation="POL" athleteid="4267">
              <RESULTS>
                <RESULT eventid="1200" points="360" reactiontime="+76" swimtime="00:00:31.76" resultid="4268" heatid="7456" lane="2" entrytime="00:00:30.90" />
                <RESULT eventid="1302" points="361" reactiontime="+87" swimtime="00:01:11.23" resultid="4269" heatid="7554" lane="3" entrytime="00:01:08.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="400" reactiontime="+82" swimtime="00:00:29.58" resultid="4270" heatid="7642" lane="3" entrytime="00:00:28.92" />
                <RESULT eventid="1470" points="313" reactiontime="+77" swimtime="00:01:12.05" resultid="4271" heatid="7671" lane="6" entrytime="00:01:09.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="4272" heatid="7748" lane="2" entrytime="00:01:09.37" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="4273" heatid="7802" lane="1" entrytime="00:00:37.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="4274">
              <RESULTS>
                <RESULT eventid="1092" points="289" reactiontime="+90" swimtime="00:03:08.33" resultid="4275" heatid="7386" lane="2" entrytime="00:03:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="100" swimtime="00:01:29.76" />
                    <SPLIT distance="150" swimtime="00:02:24.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="337" reactiontime="+89" swimtime="00:11:36.23" resultid="4276" heatid="7905" lane="6" entrytime="00:11:36.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:21.30" />
                    <SPLIT distance="150" swimtime="00:02:04.68" />
                    <SPLIT distance="200" swimtime="00:02:48.53" />
                    <SPLIT distance="250" swimtime="00:03:32.12" />
                    <SPLIT distance="300" swimtime="00:04:15.83" />
                    <SPLIT distance="350" swimtime="00:04:59.36" />
                    <SPLIT distance="400" swimtime="00:05:43.39" />
                    <SPLIT distance="450" swimtime="00:06:26.76" />
                    <SPLIT distance="500" swimtime="00:07:10.84" />
                    <SPLIT distance="550" swimtime="00:07:55.70" />
                    <SPLIT distance="600" swimtime="00:08:40.67" />
                    <SPLIT distance="650" swimtime="00:09:25.14" />
                    <SPLIT distance="700" swimtime="00:10:09.35" />
                    <SPLIT distance="750" swimtime="00:10:53.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="268" reactiontime="+89" swimtime="00:03:28.47" resultid="4277" heatid="7467" lane="1" entrytime="00:03:25.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                    <SPLIT distance="100" swimtime="00:01:41.32" />
                    <SPLIT distance="150" swimtime="00:02:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="342" swimtime="00:01:12.90" resultid="4278" heatid="7495" lane="5" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="339" swimtime="00:02:39.40" resultid="4279" heatid="7682" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:18.12" />
                    <SPLIT distance="150" swimtime="00:01:58.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K-14 (275m)" eventid="1542" reactiontime="+94" status="DSQ" swimtime="00:06:41.74" resultid="4280" heatid="7717" lane="3" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                    <SPLIT distance="100" swimtime="00:01:44.06" />
                    <SPLIT distance="150" swimtime="00:02:34.35" />
                    <SPLIT distance="200" swimtime="00:03:25.02" />
                    <SPLIT distance="250" swimtime="00:04:18.91" />
                    <SPLIT distance="300" swimtime="00:05:13.70" />
                    <SPLIT distance="350" swimtime="00:05:58.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="324" reactiontime="+88" swimtime="00:05:41.71" resultid="4281" heatid="8023" lane="2" entrytime="00:05:36.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                    <SPLIT distance="150" swimtime="00:02:07.26" />
                    <SPLIT distance="200" swimtime="00:02:51.46" />
                    <SPLIT distance="250" swimtime="00:03:35.13" />
                    <SPLIT distance="300" swimtime="00:04:18.66" />
                    <SPLIT distance="350" swimtime="00:05:01.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-26" firstname="Aleksandra" gender="F" lastname="Przybysz" nation="POL" athleteid="4282">
              <RESULTS>
                <RESULT eventid="1577" points="229" reactiontime="+102" swimtime="00:01:29.89" resultid="4283" heatid="7733" lane="1" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="300" reactiontime="+109" swimtime="00:05:50.89" resultid="4284" heatid="8023" lane="1" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:10.30" />
                    <SPLIT distance="200" swimtime="00:02:55.11" />
                    <SPLIT distance="250" swimtime="00:03:39.65" />
                    <SPLIT distance="300" swimtime="00:04:24.14" />
                    <SPLIT distance="350" swimtime="00:05:08.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="4285">
              <RESULTS>
                <RESULT eventid="1183" points="319" reactiontime="+73" swimtime="00:00:37.61" resultid="4286" heatid="7438" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1285" points="387" swimtime="00:01:19.19" resultid="4287" heatid="7534" lane="5" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="358" reactiontime="+84" swimtime="00:00:34.31" resultid="4288" heatid="7619" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1453" points="312" reactiontime="+70" swimtime="00:01:21.37" resultid="4289" heatid="7655" lane="2" entrytime="00:01:21.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="311" reactiontime="+89" swimtime="00:01:21.21" resultid="4290" heatid="7734" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="309" reactiontime="+79" swimtime="00:02:57.42" resultid="4291" heatid="7759" lane="4" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                    <SPLIT distance="100" swimtime="00:01:27.44" />
                    <SPLIT distance="150" swimtime="00:02:14.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="4292">
              <RESULTS>
                <RESULT eventid="1075" points="471" swimtime="00:00:26.08" resultid="4293" heatid="7373" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1109" points="437" swimtime="00:02:25.03" resultid="4294" heatid="7404" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="505" reactiontime="+79" swimtime="00:00:56.43" resultid="4295" heatid="7504" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="456" reactiontime="+77" swimtime="00:01:05.92" resultid="4296" heatid="7556" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="448" reactiontime="+79" swimtime="00:00:28.49" resultid="4297" heatid="7631" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1504" points="484" reactiontime="+77" swimtime="00:02:06.54" resultid="4298" heatid="7704" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                    <SPLIT distance="100" swimtime="00:01:01.45" />
                    <SPLIT distance="150" swimtime="00:01:34.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="441" swimtime="00:01:03.65" resultid="4299" heatid="7739" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="482" reactiontime="+86" swimtime="00:04:31.36" resultid="4300" heatid="8057" lane="2" entrytime="00:04:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:05.70" />
                    <SPLIT distance="150" swimtime="00:01:40.46" />
                    <SPLIT distance="200" swimtime="00:02:15.21" />
                    <SPLIT distance="250" swimtime="00:02:49.26" />
                    <SPLIT distance="300" swimtime="00:03:23.91" />
                    <SPLIT distance="350" swimtime="00:03:58.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="4301">
              <RESULTS>
                <RESULT eventid="1075" points="367" reactiontime="+88" swimtime="00:00:28.34" resultid="4302" heatid="7367" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1109" points="360" reactiontime="+90" swimtime="00:02:34.62" resultid="4303" heatid="7402" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="150" swimtime="00:01:57.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="330" reactiontime="+79" swimtime="00:00:32.70" resultid="4304" heatid="7450" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="364" reactiontime="+92" swimtime="00:01:11.03" resultid="4305" heatid="7552" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="370" reactiontime="+89" swimtime="00:00:30.35" resultid="4306" heatid="7625" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1504" points="371" reactiontime="+93" swimtime="00:02:18.20" resultid="4307" heatid="7698" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:08.37" />
                    <SPLIT distance="150" swimtime="00:01:43.84" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1594" points="364" reactiontime="+91" swimtime="00:01:07.88" resultid="4308" heatid="7744" lane="4" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="361" reactiontime="+100" swimtime="00:04:58.61" resultid="4309" heatid="8055" lane="6" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="150" swimtime="00:01:50.35" />
                    <SPLIT distance="200" swimtime="00:02:28.25" />
                    <SPLIT distance="250" swimtime="00:03:06.78" />
                    <SPLIT distance="300" swimtime="00:03:45.11" />
                    <SPLIT distance="350" swimtime="00:04:22.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-24" firstname="Przemysław" gender="M" lastname="Bielski" nation="POL" athleteid="4310">
              <RESULTS>
                <RESULT eventid="1075" points="317" swimtime="00:00:29.77" resultid="4311" heatid="7365" lane="5" entrytime="00:00:29.71" />
                <RESULT eventid="1268" points="334" reactiontime="+96" swimtime="00:01:04.77" resultid="4312" heatid="7516" lane="1" entrytime="00:01:04.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="285" reactiontime="+99" swimtime="00:00:33.10" resultid="4313" heatid="7625" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1504" points="298" reactiontime="+99" swimtime="00:02:28.65" resultid="4314" heatid="7697" lane="3" entrytime="00:02:25.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                    <SPLIT distance="150" swimtime="00:01:52.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="4315" heatid="8053" lane="6" entrytime="00:05:22.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-29" firstname="Jakub" gender="M" lastname="Stępień" nation="POL" athleteid="4316">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4317" heatid="7365" lane="6" entrytime="00:00:29.95" />
                <RESULT eventid="1268" points="297" swimtime="00:01:07.30" resultid="4318" heatid="7510" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="265" reactiontime="+91" swimtime="00:02:34.61" resultid="4319" heatid="7686" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:01:54.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="230" reactiontime="+97" swimtime="00:05:47.09" resultid="4320" heatid="8043" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                    <SPLIT distance="100" swimtime="00:01:17.35" />
                    <SPLIT distance="150" swimtime="00:02:01.35" />
                    <SPLIT distance="200" swimtime="00:02:47.48" />
                    <SPLIT distance="250" swimtime="00:03:34.31" />
                    <SPLIT distance="300" swimtime="00:04:20.36" />
                    <SPLIT distance="350" swimtime="00:05:05.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-08" firstname="Paweł" gender="M" lastname="Suchecki" nation="POL" athleteid="4321">
              <RESULTS>
                <RESULT eventid="1268" points="308" reactiontime="+87" swimtime="00:01:06.53" resultid="4322" heatid="7513" lane="4" entrytime="00:01:06.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="318" swimtime="00:00:31.92" resultid="4323" heatid="7634" lane="5" entrytime="00:00:32.04" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-13" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="4324">
              <RESULTS>
                <RESULT eventid="1109" points="433" reactiontime="+84" swimtime="00:02:25.48" resultid="4325" heatid="7403" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                    <SPLIT distance="150" swimtime="00:01:48.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="453" reactiontime="+80" swimtime="00:02:37.05" resultid="4326" heatid="7483" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:13.47" />
                    <SPLIT distance="150" swimtime="00:01:54.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="443" reactiontime="+81" swimtime="00:01:06.54" resultid="4327" heatid="7553" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="488" swimtime="00:01:10.61" resultid="4328" heatid="7609" lane="5" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="369" reactiontime="+78" swimtime="00:05:28.28" resultid="4329" heatid="7978" lane="6" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:18.99" />
                    <SPLIT distance="150" swimtime="00:02:01.65" />
                    <SPLIT distance="200" swimtime="00:02:44.18" />
                    <SPLIT distance="250" swimtime="00:03:27.00" />
                    <SPLIT distance="300" swimtime="00:04:10.27" />
                    <SPLIT distance="350" swimtime="00:04:49.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="482" reactiontime="+76" swimtime="00:00:32.20" resultid="4330" heatid="7808" lane="6" entrytime="00:00:34.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-01" firstname="Małgorzata" gender="F" lastname="Polito" nation="POL" athleteid="4331">
              <RESULTS>
                <RESULT eventid="1148" points="317" swimtime="00:11:50.48" resultid="4332" heatid="7904" lane="3" entrytime="00:11:47.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="100" swimtime="00:01:27.54" />
                    <SPLIT distance="150" swimtime="00:02:13.45" />
                    <SPLIT distance="200" swimtime="00:02:59.95" />
                    <SPLIT distance="250" swimtime="00:03:45.43" />
                    <SPLIT distance="300" swimtime="00:04:31.31" />
                    <SPLIT distance="350" swimtime="00:05:16.64" />
                    <SPLIT distance="400" swimtime="00:06:01.73" />
                    <SPLIT distance="450" swimtime="00:06:46.11" />
                    <SPLIT distance="500" swimtime="00:07:30.81" />
                    <SPLIT distance="550" swimtime="00:08:14.93" />
                    <SPLIT distance="600" swimtime="00:08:59.20" />
                    <SPLIT distance="650" swimtime="00:09:42.59" />
                    <SPLIT distance="700" swimtime="00:10:26.62" />
                    <SPLIT distance="750" swimtime="00:11:09.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="337" reactiontime="+83" swimtime="00:03:13.29" resultid="4333" heatid="7468" lane="3" entrytime="00:03:08.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                    <SPLIT distance="100" swimtime="00:01:33.49" />
                    <SPLIT distance="150" swimtime="00:02:23.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="347" swimtime="00:01:29.19" resultid="4334" heatid="7590" lane="5" entrytime="00:01:26.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="326" reactiontime="+83" swimtime="00:02:41.37" resultid="4335" heatid="7682" lane="4" entrytime="00:02:37.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:18.17" />
                    <SPLIT distance="150" swimtime="00:02:00.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="325" reactiontime="+85" swimtime="00:05:41.63" resultid="4336" heatid="8023" lane="4" entrytime="00:05:31.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:22.31" />
                    <SPLIT distance="150" swimtime="00:02:07.01" />
                    <SPLIT distance="200" swimtime="00:02:51.53" />
                    <SPLIT distance="250" swimtime="00:03:35.73" />
                    <SPLIT distance="300" swimtime="00:04:19.28" />
                    <SPLIT distance="350" swimtime="00:05:02.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-30" firstname="Karol" gender="M" lastname="Dziemian" nation="POL" athleteid="4337">
              <RESULTS>
                <RESULT eventid="1075" points="202" reactiontime="+96" swimtime="00:00:34.56" resultid="4338" heatid="7353" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1268" points="189" swimtime="00:01:18.30" resultid="4339" heatid="7505" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="155" reactiontime="+90" swimtime="00:00:40.55" resultid="4340" heatid="7626" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1504" points="164" swimtime="00:03:01.49" resultid="4341" heatid="7690" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                    <SPLIT distance="100" swimtime="00:01:27.89" />
                    <SPLIT distance="150" swimtime="00:02:15.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="210" reactiontime="+85" swimtime="00:00:42.46" resultid="4342" heatid="7793" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-01" firstname="Grzegorz" gender="M" lastname="Mówiński" nation="POL" athleteid="4343">
              <RESULTS>
                <RESULT eventid="1075" points="247" reactiontime="+86" swimtime="00:00:32.33" resultid="4344" heatid="7355" lane="6" entrytime="00:00:33.75" />
                <RESULT eventid="1336" points="194" reactiontime="+85" swimtime="00:03:08.29" resultid="4345" heatid="7568" lane="4" entrytime="00:03:08.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                    <SPLIT distance="100" swimtime="00:01:27.62" />
                    <SPLIT distance="150" swimtime="00:02:17.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="241" reactiontime="+85" swimtime="00:02:39.57" resultid="4346" heatid="7692" lane="3" entrytime="00:02:45.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:01:59.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="182" reactiontime="+91" swimtime="00:01:25.45" resultid="4347" heatid="7742" lane="2" entrytime="00:01:23.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Aquasfera Masters Olsztyn B" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="237" reactiontime="+73" swimtime="00:02:28.34" resultid="4352" heatid="7930" lane="3" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:01:54.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4321" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4316" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4343" number="3" reactiontime="+20" />
                    <RELAYPOSITION athleteid="4337" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Aquasfera Masters Olsztyn C" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="414" reactiontime="+71" swimtime="00:02:03.16" resultid="4353" heatid="7933" lane="4" entrytime="00:02:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:04.83" />
                    <SPLIT distance="150" swimtime="00:01:36.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4267" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4324" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="4301" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="4292" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Aquasfera Masters Olsztyn C" number="1">
              <RESULTS>
                <RESULT eventid="1528" points="400" reactiontime="+84" swimtime="00:01:49.55" resultid="4354" heatid="7714" lane="4" entrytime="00:01:51.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="100" swimtime="00:00:56.44" />
                    <SPLIT distance="150" swimtime="00:01:23.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4292" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="4324" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="4321" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="4267" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Aquasfera Masters Olsztyn C" number="2">
              <RESULTS>
                <RESULT eventid="1528" points="292" reactiontime="+94" swimtime="00:02:01.71" resultid="4348" heatid="7712" lane="4" entrytime="00:02:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="100" swimtime="00:00:59.72" />
                    <SPLIT distance="150" swimtime="00:01:33.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4310" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="4316" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="4337" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="4301" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Aquasfera Masters Olsztyn B" number="1">
              <RESULTS>
                <RESULT eventid="1370" points="339" reactiontime="+72" swimtime="00:02:27.25" resultid="4350" heatid="7573" lane="1" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:19.66" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4285" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4331" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="4255" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4274" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1521" points="365" reactiontime="+94" swimtime="00:02:10.40" resultid="4351" heatid="7708" lane="1" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:03.55" />
                    <SPLIT distance="150" swimtime="00:01:37.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4285" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="4255" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4331" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="4274" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Aquasfera Masters Olsztyn B" number="1">
              <RESULTS>
                <RESULT eventid="1679" points="334" reactiontime="+75" swimtime="00:02:12.21" resultid="4355" heatid="7818" lane="4" entrytime="00:02:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:09.43" />
                    <SPLIT distance="150" swimtime="00:01:37.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4255" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4324" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="4292" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="4282" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1126" points="326" swimtime="00:01:57.31" resultid="4356" heatid="7411" lane="5" entrytime="00:01:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                    <SPLIT distance="100" swimtime="00:00:53.27" />
                    <SPLIT distance="150" swimtime="00:01:24.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4292" number="1" />
                    <RELAYPOSITION athleteid="4324" number="2" />
                    <RELAYPOSITION athleteid="4255" number="3" />
                    <RELAYPOSITION athleteid="4331" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Aquasfera Masters Olsztyn C" number="1">
              <RESULTS>
                <RESULT eventid="1126" points="245" reactiontime="+104" swimtime="00:02:09.08" resultid="4349" heatid="7409" lane="3" entrytime="00:02:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:00:58.38" />
                    <SPLIT distance="150" swimtime="00:01:32.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4310" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="4301" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="4274" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="4263" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Aquasfera Masters Olsztyn C" number="2">
              <RESULTS>
                <RESULT eventid="1679" points="231" reactiontime="+85" swimtime="00:02:29.55" resultid="4357" heatid="7817" lane="5" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="150" swimtime="00:01:53.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4301" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="4331" number="2" />
                    <RELAYPOSITION athleteid="4343" number="3" />
                    <RELAYPOSITION athleteid="4263" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AWBIA" name="AZS AWF Biała Podlaska" nation="POL" region="LU">
          <CONTACT email="zielakk@gmail.com" name="Kamil Zieliński" phone="781529483" />
          <ATHLETES>
            <ATHLETE birthdate="1989-04-27" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" license="S02203200002" athleteid="4378">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4379" heatid="7377" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4380" heatid="7406" lane="5" entrytime="00:02:20.00" />
                <RESULT eventid="1234" points="570" swimtime="00:02:25.47" resultid="4381" heatid="7485" lane="5" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:10.08" />
                    <SPLIT distance="150" swimtime="00:01:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="506" reactiontime="+70" swimtime="00:01:03.67" resultid="4382" heatid="7559" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="605" reactiontime="+72" swimtime="00:01:05.74" resultid="4383" heatid="7611" lane="4" entrytime="00:01:03.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="471" reactiontime="+73" swimtime="00:00:28.00" resultid="4384" heatid="7640" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1662" points="583" reactiontime="+71" swimtime="00:00:30.21" resultid="4385" heatid="7813" lane="3" entrytime="00:00:29.26" />
                <RESULT eventid="1710" points="402" reactiontime="+76" swimtime="00:04:48.28" resultid="4386" heatid="8054" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:44.36" />
                    <SPLIT distance="200" swimtime="00:02:20.89" />
                    <SPLIT distance="250" swimtime="00:02:57.76" />
                    <SPLIT distance="300" swimtime="00:03:35.30" />
                    <SPLIT distance="350" swimtime="00:04:12.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01910" name="KS Delfin Gdynia" nation="POL" region="POM">
          <ATHLETES>
            <ATHLETE birthdate="1971-11-04" firstname="Jakub" gender="M" lastname="Mańczak" nation="POL" license="101910200065" athleteid="4388">
              <RESULTS>
                <RESULT eventid="1268" points="407" reactiontime="+77" swimtime="00:01:00.61" resultid="4389" heatid="7520" lane="6" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="290" reactiontime="+84" swimtime="00:02:44.71" resultid="4390" heatid="7570" lane="6" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="100" swimtime="00:01:16.92" />
                    <SPLIT distance="150" swimtime="00:02:01.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="397" reactiontime="+76" swimtime="00:00:29.64" resultid="4391" heatid="7641" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1504" points="342" swimtime="00:02:22.06" resultid="4392" heatid="7700" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                    <SPLIT distance="150" swimtime="00:01:46.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KRA" name="Masters Korona Kraków" nation="POL" region="MAL">
          <CONTACT city="Kraków" email="masterskorona@wp.pl" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="4394">
              <RESULTS>
                <RESULT eventid="1058" points="465" reactiontime="+79" swimtime="00:00:30.01" resultid="4395" heatid="7343" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1183" points="393" reactiontime="+62" swimtime="00:00:35.06" resultid="4396" heatid="7434" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1285" points="442" reactiontime="+73" swimtime="00:01:15.76" resultid="4397" heatid="7536" lane="6" entrytime="00:01:15.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1385" points="404" reactiontime="+84" swimtime="00:01:24.80" resultid="4398" heatid="7583" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="413" swimtime="00:00:32.72" resultid="4399" heatid="7620" lane="5" entrytime="00:00:33.50" />
                <RESULT comment="Rekord Polski Masters" eventid="1645" points="454" reactiontime="+82" swimtime="00:00:37.47" resultid="4400" heatid="7786" lane="3" entrytime="00:00:38.36" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1933-04-07" firstname="Tadeusz" gender="M" lastname="Banach" nation="POL" athleteid="4401">
              <RESULTS>
                <RESULT eventid="1075" points="16" reactiontime="+115" swimtime="00:01:20.08" resultid="4402" heatid="7345" lane="2" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="4403" heatid="7442" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-04-24" firstname="Krzysztof" gender="M" lastname="Chołda" nation="POL" athleteid="4404">
              <RESULTS>
                <RESULT eventid="1165" points="238" reactiontime="+111" swimtime="00:22:51.00" resultid="4405" heatid="7913" lane="6" entrytime="00:22:36.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                    <SPLIT distance="100" swimtime="00:01:19.99" />
                    <SPLIT distance="150" swimtime="00:02:03.71" />
                    <SPLIT distance="200" swimtime="00:02:48.00" />
                    <SPLIT distance="250" swimtime="00:04:18.20" />
                    <SPLIT distance="300" swimtime="00:05:03.41" />
                    <SPLIT distance="350" swimtime="00:05:48.74" />
                    <SPLIT distance="400" swimtime="00:06:34.82" />
                    <SPLIT distance="450" swimtime="00:08:07.74" />
                    <SPLIT distance="500" swimtime="00:09:40.98" />
                    <SPLIT distance="550" swimtime="00:10:28.16" />
                    <SPLIT distance="600" swimtime="00:11:14.88" />
                    <SPLIT distance="650" swimtime="00:12:02.28" />
                    <SPLIT distance="700" swimtime="00:12:48.13" />
                    <SPLIT distance="750" swimtime="00:13:35.21" />
                    <SPLIT distance="800" swimtime="00:14:21.60" />
                    <SPLIT distance="850" swimtime="00:15:08.59" />
                    <SPLIT distance="900" swimtime="00:15:55.79" />
                    <SPLIT distance="950" swimtime="00:16:42.65" />
                    <SPLIT distance="1000" swimtime="00:17:29.77" />
                    <SPLIT distance="1050" swimtime="00:18:16.38" />
                    <SPLIT distance="1100" swimtime="00:19:03.46" />
                    <SPLIT distance="1150" swimtime="00:19:49.79" />
                    <SPLIT distance="1200" swimtime="00:20:36.47" />
                    <SPLIT distance="1300" swimtime="00:21:23.24" />
                    <SPLIT distance="1400" swimtime="00:22:08.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="218" reactiontime="+100" swimtime="00:01:24.32" resultid="4406" heatid="7543" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="223" reactiontime="+98" swimtime="00:01:31.64" resultid="4407" heatid="7599" lane="3" entrytime="00:01:30.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="222" reactiontime="+102" swimtime="00:00:41.64" resultid="4408" heatid="7792" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1710" points="252" swimtime="00:05:36.42" resultid="4409" heatid="8051" lane="5" entrytime="00:05:35.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:16.58" />
                    <SPLIT distance="150" swimtime="00:02:39.74" />
                    <SPLIT distance="200" swimtime="00:03:23.36" />
                    <SPLIT distance="250" swimtime="00:04:07.39" />
                    <SPLIT distance="300" swimtime="00:04:52.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="Frączek" nation="POL" athleteid="4410">
              <RESULTS>
                <RESULT eventid="1058" points="470" swimtime="00:00:29.90" resultid="4411" heatid="7343" lane="5" entrytime="00:00:29.50" />
                <RESULT eventid="1251" points="458" reactiontime="+78" swimtime="00:01:06.17" resultid="4412" heatid="7497" lane="1" entrytime="00:01:06.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" status="DNS" swimtime="00:00:00.00" resultid="4413" heatid="7535" lane="4" entrytime="00:01:16.00" />
                <RESULT eventid="1419" points="370" reactiontime="+76" swimtime="00:00:33.95" resultid="4414" heatid="7619" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1453" points="297" reactiontime="+72" swimtime="00:01:22.75" resultid="4415" heatid="7656" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-09-19" firstname="Maciej" gender="M" lastname="Grudzień" nation="POL" athleteid="4416">
              <RESULTS>
                <RESULT eventid="1109" points="216" reactiontime="+93" swimtime="00:03:03.21" resultid="4417" heatid="7396" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                    <SPLIT distance="100" swimtime="00:01:30.69" />
                    <SPLIT distance="150" swimtime="00:02:23.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="191" reactiontime="+101" swimtime="00:03:29.49" resultid="4418" heatid="7477" lane="6" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.60" />
                    <SPLIT distance="100" swimtime="00:01:42.62" />
                    <SPLIT distance="150" swimtime="00:02:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="196" reactiontime="+82" swimtime="00:03:02.41" resultid="4419" heatid="7766" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:01:27.62" />
                    <SPLIT distance="150" swimtime="00:02:15.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-12" firstname="Wojciech" gender="M" lastname="Hoffman" nation="POL" athleteid="4420">
              <RESULTS>
                <RESULT eventid="1165" points="333" reactiontime="+86" swimtime="00:20:26.16" resultid="4421" heatid="7914" lane="3" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                    <SPLIT distance="100" swimtime="00:01:14.80" />
                    <SPLIT distance="150" swimtime="00:01:55.46" />
                    <SPLIT distance="200" swimtime="00:02:35.94" />
                    <SPLIT distance="250" swimtime="00:03:16.44" />
                    <SPLIT distance="300" swimtime="00:03:57.82" />
                    <SPLIT distance="350" swimtime="00:04:38.53" />
                    <SPLIT distance="400" swimtime="00:05:18.90" />
                    <SPLIT distance="450" swimtime="00:05:59.85" />
                    <SPLIT distance="500" swimtime="00:06:42.10" />
                    <SPLIT distance="550" swimtime="00:07:23.03" />
                    <SPLIT distance="600" swimtime="00:08:05.04" />
                    <SPLIT distance="650" swimtime="00:08:46.47" />
                    <SPLIT distance="700" swimtime="00:09:27.82" />
                    <SPLIT distance="750" swimtime="00:10:09.09" />
                    <SPLIT distance="800" swimtime="00:10:49.27" />
                    <SPLIT distance="850" swimtime="00:11:30.19" />
                    <SPLIT distance="900" swimtime="00:12:11.79" />
                    <SPLIT distance="950" swimtime="00:12:53.41" />
                    <SPLIT distance="1000" swimtime="00:13:36.05" />
                    <SPLIT distance="1050" swimtime="00:14:18.03" />
                    <SPLIT distance="1100" swimtime="00:14:59.40" />
                    <SPLIT distance="1150" swimtime="00:15:41.76" />
                    <SPLIT distance="1200" swimtime="00:16:21.70" />
                    <SPLIT distance="1250" swimtime="00:17:03.93" />
                    <SPLIT distance="1300" swimtime="00:17:45.65" />
                    <SPLIT distance="1350" swimtime="00:18:27.49" />
                    <SPLIT distance="1400" swimtime="00:19:07.65" />
                    <SPLIT distance="1450" swimtime="00:19:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="338" reactiontime="+77" swimtime="00:01:04.50" resultid="4422" heatid="7516" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="339" swimtime="00:02:22.48" resultid="4423" heatid="7698" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:09.27" />
                    <SPLIT distance="150" swimtime="00:01:46.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="347" reactiontime="+84" swimtime="00:05:02.65" resultid="4424" heatid="8054" lane="1" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                    <SPLIT distance="150" swimtime="00:01:50.47" />
                    <SPLIT distance="200" swimtime="00:02:28.82" />
                    <SPLIT distance="250" swimtime="00:03:07.28" />
                    <SPLIT distance="300" swimtime="00:03:45.56" />
                    <SPLIT distance="350" swimtime="00:04:25.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="4425">
              <RESULTS>
                <RESULT eventid="1058" points="332" reactiontime="+92" swimtime="00:00:33.56" resultid="4426" heatid="7339" lane="2" entrytime="00:00:34.50" />
                <RESULT eventid="1183" points="274" reactiontime="+85" swimtime="00:00:39.54" resultid="4427" heatid="7437" lane="5" entrytime="00:00:39.95" />
                <RESULT eventid="1285" status="DNS" swimtime="00:00:00.00" resultid="4428" heatid="7529" lane="1" entrytime="00:01:35.00" />
                <RESULT eventid="1419" points="299" swimtime="00:00:36.44" resultid="4429" heatid="7618" lane="5" entrytime="00:00:36.80" />
                <RESULT eventid="1453" points="225" reactiontime="+86" swimtime="00:01:30.78" resultid="4430" heatid="7651" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="142" reactiontime="+99" swimtime="00:01:45.47" resultid="4431" heatid="7732" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="218" reactiontime="+87" swimtime="00:03:19.38" resultid="4432" heatid="7757" lane="6" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                    <SPLIT distance="100" swimtime="00:01:38.37" />
                    <SPLIT distance="150" swimtime="00:02:31.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-26" firstname="Anna" gender="F" lastname="Kasprzykowska" nation="POL" athleteid="4433">
              <RESULTS>
                <RESULT eventid="1251" points="130" reactiontime="+98" swimtime="00:01:40.62" resultid="4434" heatid="7487" lane="3" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="104" swimtime="00:00:51.79" resultid="4435" heatid="7613" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1487" points="111" reactiontime="+104" swimtime="00:03:50.84" resultid="4436" heatid="7676" lane="1" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.98" />
                    <SPLIT distance="100" swimtime="00:01:50.88" />
                    <SPLIT distance="150" swimtime="00:02:50.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-07-26" firstname="Anna" gender="F" lastname="Koźmin" nation="POL" athleteid="4437">
              <RESULTS>
                <RESULT eventid="1092" points="102" reactiontime="+110" swimtime="00:04:25.84" resultid="4438" heatid="7383" lane="4" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.53" />
                    <SPLIT distance="100" swimtime="00:02:09.40" />
                    <SPLIT distance="150" swimtime="00:03:20.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="112" reactiontime="+120" swimtime="00:04:39.08" resultid="4439" heatid="7464" lane="6" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.77" />
                    <SPLIT distance="100" swimtime="00:02:13.19" />
                    <SPLIT distance="150" swimtime="00:03:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="108" reactiontime="+122" swimtime="00:02:01.00" resultid="4440" heatid="7527" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="101" reactiontime="+119" swimtime="00:00:52.27" resultid="4441" heatid="7613" lane="3" entrytime="00:00:52.00" />
                <RESULT eventid="1645" points="170" reactiontime="+113" swimtime="00:00:51.89" resultid="4442" heatid="7779" lane="1" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-06-03" firstname="Antoni" gender="M" lastname="Kubis" nation="POL" athleteid="4443">
              <RESULTS>
                <RESULT eventid="1075" points="125" swimtime="00:00:40.54" resultid="4444" heatid="7348" lane="5" entrytime="00:00:47.00" />
                <RESULT eventid="1302" points="120" reactiontime="+123" swimtime="00:01:42.66" resultid="4445" heatid="7540" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="100" swimtime="00:01:59.79" resultid="4446" heatid="7595" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="4447" heatid="7790" lane="4" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-24" firstname="Bogusław" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="4448">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4449" heatid="7348" lane="6" entrytime="00:00:58.00" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="4450" heatid="7442" lane="3" entrytime="00:01:15.00" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="4451" heatid="7501" lane="1" entrytime="00:02:24.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="4452" heatid="7594" lane="6" entrytime="00:02:57.00" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="4453" heatid="7660" lane="3" entrytime="00:02:40.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="4454" heatid="7790" lane="6" entrytime="00:01:17.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-16" firstname="Kamil" gender="M" lastname="Latuszek" nation="POL" athleteid="4455">
              <RESULTS>
                <RESULT eventid="1075" points="474" reactiontime="+79" swimtime="00:00:26.02" resultid="4456" heatid="7373" lane="2" entrytime="00:00:27.00" />
                <RESULT eventid="1268" points="473" reactiontime="+78" swimtime="00:00:57.65" resultid="4457" heatid="7522" lane="6" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="411" reactiontime="+79" swimtime="00:00:29.32" resultid="4458" heatid="7639" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1504" points="375" reactiontime="+82" swimtime="00:02:17.79" resultid="4459" heatid="7700" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:08.36" />
                    <SPLIT distance="150" swimtime="00:01:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="344" swimtime="00:01:09.16" resultid="4460" heatid="7746" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="4461">
              <RESULTS>
                <RESULT eventid="1058" points="241" reactiontime="+99" swimtime="00:00:37.32" resultid="4462" heatid="7332" lane="1" />
                <RESULT eventid="1092" points="180" reactiontime="+110" swimtime="00:03:40.64" resultid="4463" heatid="7385" lane="6" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.55" />
                    <SPLIT distance="100" swimtime="00:01:45.04" />
                    <SPLIT distance="150" swimtime="00:02:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" status="DNS" swimtime="00:00:00.00" resultid="4464" heatid="7434" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1319" points="133" reactiontime="+114" swimtime="00:03:56.59" resultid="4465" heatid="7561" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.85" />
                    <SPLIT distance="100" swimtime="00:01:53.62" />
                    <SPLIT distance="150" swimtime="00:02:55.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="175" reactiontime="+108" swimtime="00:00:43.54" resultid="4466" heatid="7612" lane="2" />
                <RESULT eventid="1487" points="179" reactiontime="+113" swimtime="00:03:17.11" resultid="4467" heatid="7678" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:33.21" />
                    <SPLIT distance="150" swimtime="00:02:24.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="133" reactiontime="+120" swimtime="00:01:47.84" resultid="4468" heatid="7730" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="181" reactiontime="+118" swimtime="00:06:55.26" resultid="4469" heatid="8018" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                    <SPLIT distance="100" swimtime="00:01:37.26" />
                    <SPLIT distance="150" swimtime="00:02:30.25" />
                    <SPLIT distance="200" swimtime="00:03:24.17" />
                    <SPLIT distance="250" swimtime="00:04:16.48" />
                    <SPLIT distance="300" swimtime="00:05:10.39" />
                    <SPLIT distance="350" swimtime="00:06:05.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="4470">
              <RESULTS>
                <RESULT eventid="1092" points="244" reactiontime="+104" swimtime="00:03:19.36" resultid="4471" heatid="7382" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:01:34.02" />
                    <SPLIT distance="150" swimtime="00:02:34.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="257" reactiontime="+104" swimtime="00:12:41.28" resultid="4472" heatid="7904" lane="6" entrytime="00:13:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:24.48" />
                    <SPLIT distance="150" swimtime="00:02:11.69" />
                    <SPLIT distance="200" swimtime="00:02:59.11" />
                    <SPLIT distance="250" swimtime="00:03:46.65" />
                    <SPLIT distance="300" swimtime="00:04:34.64" />
                    <SPLIT distance="350" swimtime="00:05:23.35" />
                    <SPLIT distance="400" swimtime="00:06:12.17" />
                    <SPLIT distance="450" swimtime="00:07:01.29" />
                    <SPLIT distance="500" swimtime="00:07:50.52" />
                    <SPLIT distance="550" swimtime="00:08:40.12" />
                    <SPLIT distance="600" swimtime="00:09:29.12" />
                    <SPLIT distance="650" swimtime="00:10:17.83" />
                    <SPLIT distance="700" swimtime="00:11:07.06" />
                    <SPLIT distance="750" swimtime="00:11:55.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="260" reactiontime="+104" swimtime="00:01:30.43" resultid="4473" heatid="7526" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="200" swimtime="00:03:26.51" resultid="4474" heatid="7561" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                    <SPLIT distance="100" swimtime="00:01:35.12" />
                    <SPLIT distance="150" swimtime="00:02:31.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="202" swimtime="00:00:41.50" resultid="4475" heatid="7612" lane="5" />
                <RESULT eventid="1487" points="271" reactiontime="+99" swimtime="00:02:51.72" resultid="4476" heatid="7680" lane="1" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                    <SPLIT distance="150" swimtime="00:02:09.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="209" reactiontime="+91" swimtime="00:01:32.74" resultid="4477" heatid="7730" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="241" reactiontime="+113" swimtime="00:06:17.41" resultid="4478" heatid="8021" lane="4" entrytime="00:06:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:25.59" />
                    <SPLIT distance="150" swimtime="00:02:14.24" />
                    <SPLIT distance="200" swimtime="00:03:02.87" />
                    <SPLIT distance="250" swimtime="00:03:51.47" />
                    <SPLIT distance="300" swimtime="00:04:40.49" />
                    <SPLIT distance="350" swimtime="00:05:29.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="4479">
              <RESULTS>
                <RESULT eventid="1075" points="217" reactiontime="+120" swimtime="00:00:33.78" resultid="4480" heatid="7357" lane="4" entrytime="00:00:32.50" />
                <RESULT eventid="1165" reactiontime="+146" status="DNF" swimtime="00:00:00.00" resultid="4481" heatid="7909" lane="2" entrytime="00:26:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="100" swimtime="00:02:46.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="221" reactiontime="+114" swimtime="00:01:14.25" resultid="4482" heatid="7508" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="74" swimtime="00:04:19.86" resultid="4483" heatid="7566" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.34" />
                    <SPLIT distance="100" swimtime="00:02:07.85" />
                    <SPLIT distance="150" swimtime="00:03:12.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="168" reactiontime="+124" swimtime="00:02:59.89" resultid="4484" heatid="7692" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:25.54" />
                    <SPLIT distance="150" swimtime="00:02:13.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="97" reactiontime="+141" swimtime="00:08:31.03" resultid="4485" heatid="7976" lane="6" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.58" />
                    <SPLIT distance="100" swimtime="00:02:07.38" />
                    <SPLIT distance="150" swimtime="00:03:11.23" />
                    <SPLIT distance="200" swimtime="00:04:17.61" />
                    <SPLIT distance="250" swimtime="00:05:25.33" />
                    <SPLIT distance="300" swimtime="00:06:36.94" />
                    <SPLIT distance="350" swimtime="00:07:35.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="80" reactiontime="+124" swimtime="00:01:52.36" resultid="4486" heatid="7740" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="135" reactiontime="+130" swimtime="00:06:54.23" resultid="4487" heatid="8048" lane="6" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                    <SPLIT distance="100" swimtime="00:01:36.81" />
                    <SPLIT distance="150" swimtime="00:02:30.08" />
                    <SPLIT distance="200" swimtime="00:03:24.87" />
                    <SPLIT distance="250" swimtime="00:04:19.31" />
                    <SPLIT distance="300" swimtime="00:05:12.99" />
                    <SPLIT distance="350" swimtime="00:06:06.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="4488">
              <RESULTS>
                <RESULT eventid="1058" points="54" reactiontime="+108" swimtime="00:01:01.25" resultid="4489" heatid="7333" lane="1" entrytime="00:00:59.00" />
                <RESULT eventid="1092" points="58" reactiontime="+113" swimtime="00:05:21.75" resultid="4490" heatid="7382" lane="3" entrytime="00:05:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.77" />
                    <SPLIT distance="100" swimtime="00:02:43.66" />
                    <SPLIT distance="150" swimtime="00:04:09.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="71" reactiontime="+106" swimtime="00:05:24.23" resultid="4491" heatid="7462" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.81" />
                    <SPLIT distance="100" swimtime="00:02:32.69" />
                    <SPLIT distance="150" swimtime="00:04:00.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="60" reactiontime="+115" swimtime="00:02:09.85" resultid="4492" heatid="7487" lane="6" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="39" reactiontime="+108" swimtime="00:01:11.43" resultid="4493" heatid="7613" lane="6" entrytime="00:01:15.00" />
                <RESULT eventid="1487" points="56" reactiontime="+106" swimtime="00:04:49.88" resultid="4494" heatid="7675" lane="4" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.33" />
                    <SPLIT distance="100" swimtime="00:02:17.07" />
                    <SPLIT distance="150" swimtime="00:03:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="90" reactiontime="+109" swimtime="00:01:04.09" resultid="4495" heatid="7776" lane="4" entrytime="00:01:01.00" />
                <RESULT eventid="1693" points="59" reactiontime="+113" swimtime="00:10:03.07" resultid="4496" heatid="8019" lane="1" entrytime="00:09:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.37" />
                    <SPLIT distance="100" swimtime="00:02:15.77" />
                    <SPLIT distance="150" swimtime="00:04:47.34" />
                    <SPLIT distance="200" swimtime="00:06:07.27" />
                    <SPLIT distance="250" swimtime="00:07:24.62" />
                    <SPLIT distance="300" swimtime="00:08:48.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="Palmowska" nation="POL" athleteid="4497">
              <RESULTS>
                <RESULT eventid="1092" points="470" reactiontime="+66" swimtime="00:02:40.21" resultid="4498" heatid="7388" lane="3" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="150" swimtime="00:02:02.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="449" reactiontime="+72" swimtime="00:00:33.54" resultid="4499" heatid="7440" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1285" points="482" reactiontime="+73" swimtime="00:01:13.60" resultid="4500" heatid="7535" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="464" reactiontime="+62" swimtime="00:01:11.34" resultid="4501" heatid="7658" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="442" reactiontime="+63" swimtime="00:02:37.54" resultid="4502" heatid="7761" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:15.02" />
                    <SPLIT distance="150" swimtime="00:01:56.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="412" reactiontime="+70" swimtime="00:05:15.49" resultid="4503" heatid="8024" lane="6" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:01:50.94" />
                    <SPLIT distance="200" swimtime="00:02:31.10" />
                    <SPLIT distance="250" swimtime="00:03:12.38" />
                    <SPLIT distance="300" swimtime="00:03:53.99" />
                    <SPLIT distance="350" swimtime="00:04:35.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="4504">
              <RESULTS>
                <RESULT eventid="1075" points="316" swimtime="00:00:29.80" resultid="4505" heatid="7366" lane="5" entrytime="00:00:29.21" />
                <RESULT eventid="1200" points="246" reactiontime="+81" swimtime="00:00:36.04" resultid="4506" heatid="7450" lane="6" entrytime="00:00:35.63" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="4507" heatid="7548" lane="3" entrytime="00:01:15.28" />
                <RESULT eventid="1436" points="335" swimtime="00:00:31.36" resultid="4508" heatid="7636" lane="5" entrytime="00:00:31.60" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="4509" heatid="7666" lane="5" entrytime="00:01:19.21" />
                <RESULT eventid="1662" points="301" reactiontime="+91" swimtime="00:00:37.66" resultid="4511" heatid="7803" lane="1" entrytime="00:00:37.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-18" firstname="Bartosz" gender="M" lastname="Próchniewicz" nation="POL" athleteid="4512">
              <RESULTS>
                <RESULT eventid="1200" points="117" reactiontime="+68" swimtime="00:00:46.10" resultid="4513" heatid="7444" lane="5" entrytime="00:00:52.00" />
                <RESULT eventid="1470" points="113" reactiontime="+74" swimtime="00:01:41.20" resultid="4514" heatid="7662" lane="1" entrytime="00:01:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-02-21" firstname="Adam" gender="M" lastname="Pycia" nation="POL" athleteid="4515">
              <RESULTS>
                <RESULT eventid="1268" points="258" reactiontime="+108" swimtime="00:01:10.52" resultid="4516" heatid="7509" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="208" reactiontime="+118" swimtime="00:01:33.72" resultid="4517" heatid="7596" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="216" reactiontime="+116" swimtime="00:02:45.37" resultid="4518" heatid="7693" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="150" swimtime="00:02:02.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-22" firstname="Alicja" gender="F" lastname="Romańska" nation="POL" athleteid="4519">
              <RESULTS>
                <RESULT eventid="1251" points="148" reactiontime="+99" swimtime="00:01:36.23" resultid="4520" heatid="7488" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="81" reactiontime="+103" swimtime="00:00:56.26" resultid="4521" heatid="7613" lane="1" entrytime="00:00:58.00" />
                <RESULT eventid="1487" points="151" reactiontime="+106" swimtime="00:03:28.74" resultid="4522" heatid="7677" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.67" />
                    <SPLIT distance="100" swimtime="00:01:43.60" />
                    <SPLIT distance="150" swimtime="00:02:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="136" reactiontime="+101" swimtime="00:00:55.92" resultid="4523" heatid="7779" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1693" points="150" reactiontime="+103" swimtime="00:07:21.24" resultid="4524" heatid="8020" lane="6" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.96" />
                    <SPLIT distance="100" swimtime="00:01:48.38" />
                    <SPLIT distance="150" swimtime="00:02:44.26" />
                    <SPLIT distance="200" swimtime="00:03:40.37" />
                    <SPLIT distance="250" swimtime="00:04:35.31" />
                    <SPLIT distance="300" swimtime="00:05:30.49" />
                    <SPLIT distance="350" swimtime="00:06:25.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="4525">
              <RESULTS>
                <RESULT eventid="1075" points="98" reactiontime="+107" swimtime="00:00:44.03" resultid="4526" heatid="7348" lane="3" entrytime="00:00:42.00" />
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1165" reactiontime="+92" status="DSQ" swimtime="00:31:21.34" resultid="4527" heatid="7907" lane="3" entrytime="00:41:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.17" />
                    <SPLIT distance="100" swimtime="00:01:55.48" />
                    <SPLIT distance="150" swimtime="00:02:58.29" />
                    <SPLIT distance="200" swimtime="00:04:02.03" />
                    <SPLIT distance="250" swimtime="00:05:05.05" />
                    <SPLIT distance="300" swimtime="00:06:09.99" />
                    <SPLIT distance="350" swimtime="00:07:12.63" />
                    <SPLIT distance="400" swimtime="00:08:16.97" />
                    <SPLIT distance="450" swimtime="00:09:21.20" />
                    <SPLIT distance="500" swimtime="00:10:24.84" />
                    <SPLIT distance="550" swimtime="00:11:27.72" />
                    <SPLIT distance="600" swimtime="00:12:31.27" />
                    <SPLIT distance="650" swimtime="00:13:35.35" />
                    <SPLIT distance="700" swimtime="00:14:39.17" />
                    <SPLIT distance="750" swimtime="00:15:42.62" />
                    <SPLIT distance="800" swimtime="00:16:46.25" />
                    <SPLIT distance="850" swimtime="00:17:49.70" />
                    <SPLIT distance="900" swimtime="00:18:53.32" />
                    <SPLIT distance="950" swimtime="00:19:56.48" />
                    <SPLIT distance="1000" swimtime="00:21:00.58" />
                    <SPLIT distance="1050" swimtime="00:22:03.81" />
                    <SPLIT distance="1100" swimtime="00:23:06.67" />
                    <SPLIT distance="1150" swimtime="00:24:09.12" />
                    <SPLIT distance="1200" swimtime="00:25:12.38" />
                    <SPLIT distance="1250" swimtime="00:26:14.19" />
                    <SPLIT distance="1300" swimtime="00:27:16.23" />
                    <SPLIT distance="1350" swimtime="00:28:19.17" />
                    <SPLIT distance="1400" swimtime="00:29:21.21" />
                    <SPLIT distance="1450" swimtime="00:30:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="22" reactiontime="+89" swimtime="00:01:20.40" resultid="4528" heatid="7443" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1268" points="88" reactiontime="+98" swimtime="00:01:40.76" resultid="4529" heatid="7501" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="4530" heatid="7661" lane="3" entrytime="00:02:00.00" />
                <RESULT eventid="1504" points="84" reactiontime="+111" swimtime="00:03:46.15" resultid="4531" heatid="7688" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.42" />
                    <SPLIT distance="100" swimtime="00:01:48.34" />
                    <SPLIT distance="150" swimtime="00:02:47.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="88" reactiontime="+134" swimtime="00:07:57.05" resultid="4532" heatid="8045" lane="6" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                    <SPLIT distance="100" swimtime="00:01:51.55" />
                    <SPLIT distance="150" swimtime="00:02:53.26" />
                    <SPLIT distance="200" swimtime="00:03:55.24" />
                    <SPLIT distance="250" swimtime="00:04:56.42" />
                    <SPLIT distance="300" swimtime="00:05:57.73" />
                    <SPLIT distance="350" swimtime="00:06:59.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="4533">
              <RESULTS>
                <RESULT eventid="1092" points="325" reactiontime="+83" swimtime="00:03:01.07" resultid="4534" heatid="7386" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:24.74" />
                    <SPLIT distance="150" swimtime="00:02:18.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="321" swimtime="00:01:24.28" resultid="4535" heatid="7530" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="304" reactiontime="+80" swimtime="00:00:36.24" resultid="4536" heatid="7618" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1487" points="283" swimtime="00:02:49.29" resultid="4537" heatid="7679" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:20.92" />
                    <SPLIT distance="150" swimtime="00:02:04.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="286" swimtime="00:01:23.51" resultid="4538" heatid="7733" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="Wysocka" nation="POL" athleteid="4539">
              <RESULTS>
                <RESULT eventid="1058" points="283" reactiontime="+94" swimtime="00:00:35.40" resultid="4540" heatid="7339" lane="4" entrytime="00:00:34.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1217" points="329" reactiontime="+90" swimtime="00:03:14.80" resultid="4541" heatid="7467" lane="4" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                    <SPLIT distance="100" swimtime="00:01:32.45" />
                    <SPLIT distance="150" swimtime="00:02:23.60" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1385" points="342" reactiontime="+93" swimtime="00:01:29.61" resultid="4542" heatid="7588" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="4543" heatid="7652" lane="6" entrytime="00:01:35.00" />
                <RESULT eventid="1645" points="324" reactiontime="+93" swimtime="00:00:41.91" resultid="4544" heatid="7785" lane="6" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-12-07" firstname="Jarosław" gender="M" lastname="Zadożny" nation="POL" athleteid="4545">
              <RESULTS>
                <RESULT eventid="1075" points="197" reactiontime="+88" swimtime="00:00:34.86" resultid="4546" heatid="7356" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1165" points="207" swimtime="00:23:55.23" resultid="4547" heatid="7910" lane="5" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="150" swimtime="00:02:10.28" />
                    <SPLIT distance="200" swimtime="00:02:56.43" />
                    <SPLIT distance="250" swimtime="00:03:42.97" />
                    <SPLIT distance="300" swimtime="00:04:29.95" />
                    <SPLIT distance="350" swimtime="00:05:17.13" />
                    <SPLIT distance="400" swimtime="00:06:04.99" />
                    <SPLIT distance="450" swimtime="00:06:52.84" />
                    <SPLIT distance="500" swimtime="00:07:40.80" />
                    <SPLIT distance="550" swimtime="00:08:29.11" />
                    <SPLIT distance="600" swimtime="00:09:17.91" />
                    <SPLIT distance="650" swimtime="00:10:06.76" />
                    <SPLIT distance="700" swimtime="00:10:56.06" />
                    <SPLIT distance="750" swimtime="00:11:45.42" />
                    <SPLIT distance="800" swimtime="00:12:34.85" />
                    <SPLIT distance="850" swimtime="00:13:24.21" />
                    <SPLIT distance="900" swimtime="00:14:13.46" />
                    <SPLIT distance="950" swimtime="00:15:02.72" />
                    <SPLIT distance="1000" swimtime="00:15:52.12" />
                    <SPLIT distance="1050" swimtime="00:16:40.82" />
                    <SPLIT distance="1100" swimtime="00:17:30.77" />
                    <SPLIT distance="1150" swimtime="00:18:19.30" />
                    <SPLIT distance="1200" swimtime="00:19:10.06" />
                    <SPLIT distance="1250" swimtime="00:19:58.90" />
                    <SPLIT distance="1300" swimtime="00:20:47.25" />
                    <SPLIT distance="1350" swimtime="00:21:36.12" />
                    <SPLIT distance="1400" swimtime="00:22:25.04" />
                    <SPLIT distance="1450" swimtime="00:23:13.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="219" reactiontime="+94" swimtime="00:05:52.95" resultid="4548" heatid="8050" lane="2" entrytime="00:05:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:19.47" />
                    <SPLIT distance="150" swimtime="00:02:03.53" />
                    <SPLIT distance="200" swimtime="00:02:50.16" />
                    <SPLIT distance="250" swimtime="00:03:37.01" />
                    <SPLIT distance="300" swimtime="00:04:23.93" />
                    <SPLIT distance="350" swimtime="00:05:10.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-05-14" firstname="Piotr" gender="M" lastname="Kowalski" nation="POL" athleteid="4549">
              <RESULTS>
                <RESULT eventid="1268" points="220" swimtime="00:01:14.41" resultid="4550" heatid="7507" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="168" reactiontime="+81" swimtime="00:00:39.48" resultid="4551" heatid="7627" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1504" points="202" reactiontime="+84" swimtime="00:02:49.32" resultid="4552" heatid="7690" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:19.16" />
                    <SPLIT distance="150" swimtime="00:02:05.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-02" firstname="Wojciech" gender="M" lastname="Kaczmarczyk" nation="POL" athleteid="4553">
              <RESULTS>
                <RESULT eventid="1075" points="71" swimtime="00:00:48.82" resultid="4554" heatid="7346" lane="5" />
                <RESULT eventid="1234" points="107" reactiontime="+128" swimtime="00:04:13.94" resultid="4555" heatid="7470" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.46" />
                    <SPLIT distance="100" swimtime="00:01:59.88" />
                    <SPLIT distance="150" swimtime="00:03:09.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="114" reactiontime="+114" swimtime="00:01:54.50" resultid="4556" heatid="7593" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-04" firstname="Andrzej" gender="M" lastname="Data" nation="POL" athleteid="4557">
              <RESULTS>
                <RESULT eventid="1165" points="175" reactiontime="+120" swimtime="00:25:18.74" resultid="4558" heatid="7912" lane="3" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:23.06" />
                    <SPLIT distance="150" swimtime="00:02:10.30" />
                    <SPLIT distance="200" swimtime="00:02:59.58" />
                    <SPLIT distance="250" swimtime="00:03:49.29" />
                    <SPLIT distance="300" swimtime="00:04:39.53" />
                    <SPLIT distance="350" swimtime="00:05:30.05" />
                    <SPLIT distance="400" swimtime="00:06:20.90" />
                    <SPLIT distance="450" swimtime="00:07:11.61" />
                    <SPLIT distance="500" swimtime="00:08:02.71" />
                    <SPLIT distance="550" swimtime="00:08:54.54" />
                    <SPLIT distance="600" swimtime="00:09:45.74" />
                    <SPLIT distance="650" swimtime="00:10:36.87" />
                    <SPLIT distance="700" swimtime="00:11:28.28" />
                    <SPLIT distance="750" swimtime="00:12:20.18" />
                    <SPLIT distance="800" swimtime="00:13:11.67" />
                    <SPLIT distance="850" swimtime="00:14:02.59" />
                    <SPLIT distance="900" swimtime="00:14:54.33" />
                    <SPLIT distance="950" swimtime="00:15:47.59" />
                    <SPLIT distance="1000" swimtime="00:16:39.18" />
                    <SPLIT distance="1050" swimtime="00:17:31.21" />
                    <SPLIT distance="1100" swimtime="00:18:24.08" />
                    <SPLIT distance="1150" swimtime="00:19:16.18" />
                    <SPLIT distance="1200" swimtime="00:20:09.28" />
                    <SPLIT distance="1250" swimtime="00:21:02.19" />
                    <SPLIT distance="1300" swimtime="00:21:54.55" />
                    <SPLIT distance="1350" swimtime="00:22:47.80" />
                    <SPLIT distance="1400" swimtime="00:23:38.91" />
                    <SPLIT distance="1450" swimtime="00:24:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="162" reactiontime="+108" swimtime="00:03:41.08" resultid="4559" heatid="7475" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="100" swimtime="00:01:41.48" />
                    <SPLIT distance="150" swimtime="00:02:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="167" reactiontime="+113" swimtime="00:01:32.07" resultid="4560" heatid="7541" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="4561" heatid="7598" lane="1" entrytime="00:01:35.00" />
                <RESULT eventid="1504" points="173" swimtime="00:02:58.27" resultid="4562" heatid="7692" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:23.96" />
                    <SPLIT distance="150" swimtime="00:02:11.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="4563" heatid="7793" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1710" points="170" swimtime="00:06:23.41" resultid="4564" heatid="8048" lane="5" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:24.11" />
                    <SPLIT distance="150" swimtime="00:02:12.39" />
                    <SPLIT distance="200" swimtime="00:03:01.96" />
                    <SPLIT distance="250" swimtime="00:03:52.59" />
                    <SPLIT distance="300" swimtime="00:04:44.32" />
                    <SPLIT distance="350" swimtime="00:05:34.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-16" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="4565">
              <RESULTS>
                <RESULT eventid="1075" points="88" reactiontime="+91" swimtime="00:00:45.62" resultid="4566" heatid="7348" lane="2" entrytime="00:00:46.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4567" heatid="7391" lane="4" entrytime="00:04:45.00" />
                <RESULT eventid="1268" points="81" reactiontime="+127" swimtime="00:01:43.76" resultid="4568" heatid="7501" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="38" reactiontime="+123" swimtime="00:02:29.73" resultid="4569" heatid="7539" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="21" reactiontime="+112" swimtime="00:01:18.78" resultid="4570" heatid="7623" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="4571" heatid="7687" lane="3" entrytime="00:04:03.00" />
                <RESULT eventid="1628" points="37" reactiontime="+76" swimtime="00:05:16.72" resultid="4572" heatid="7763" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.88" />
                    <SPLIT distance="100" swimtime="00:02:35.49" />
                    <SPLIT distance="150" swimtime="00:03:57.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="58" reactiontime="+134" swimtime="00:09:06.69" resultid="4573" heatid="8044" lane="4" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.90" />
                    <SPLIT distance="100" swimtime="00:01:59.67" />
                    <SPLIT distance="150" swimtime="00:03:08.48" />
                    <SPLIT distance="200" swimtime="00:04:19.13" />
                    <SPLIT distance="250" swimtime="00:05:29.49" />
                    <SPLIT distance="300" swimtime="00:06:42.19" />
                    <SPLIT distance="350" swimtime="00:07:54.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Masters Korona E" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="147" reactiontime="+71" swimtime="00:02:53.79" resultid="4582" heatid="7930" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.37" />
                    <SPLIT distance="100" swimtime="00:01:48.61" />
                    <SPLIT distance="150" swimtime="00:02:19.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4565" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4404" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4504" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4479" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="199" reactiontime="+97" swimtime="00:02:18.18" resultid="4583" heatid="7711" lane="1" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:48.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4525" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="4404" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="4479" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4504" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="Masters Korona C" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1521" points="438" reactiontime="+70" swimtime="00:02:02.72" resultid="4578" heatid="7708" lane="4" entrytime="00:02:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:00:59.82" />
                    <SPLIT distance="150" swimtime="00:01:33.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4497" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4394" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4425" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="4410" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Masters Korona E" number="2">
              <RESULTS>
                <RESULT eventid="1521" points="273" swimtime="00:02:23.58" resultid="4579" heatid="7707" lane="5" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                    <SPLIT distance="150" swimtime="00:01:48.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4533" number="1" />
                    <RELAYPOSITION athleteid="4470" number="2" />
                    <RELAYPOSITION athleteid="4461" number="3" />
                    <RELAYPOSITION athleteid="4539" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Masters Korona C" number="3">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1370" points="343" reactiontime="+61" swimtime="00:02:26.61" resultid="4580" heatid="7573" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:01:52.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4394" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4539" number="2" />
                    <RELAYPOSITION athleteid="4410" number="3" />
                    <RELAYPOSITION athleteid="4470" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Masters Korona D" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1126" points="294" swimtime="00:02:01.44" resultid="4574" heatid="7410" lane="5" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="100" swimtime="00:00:59.03" />
                    <SPLIT distance="150" swimtime="00:01:32.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4504" number="1" />
                    <RELAYPOSITION athleteid="4394" number="2" />
                    <RELAYPOSITION athleteid="4479" number="3" />
                    <RELAYPOSITION athleteid="4410" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" points="291" reactiontime="+62" swimtime="00:02:18.42" resultid="4575" heatid="7818" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:45.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4394" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4504" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="4410" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4479" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Masters Korona E" number="2">
              <RESULTS>
                <RESULT eventid="1126" points="141" reactiontime="+100" swimtime="00:02:35.14" resultid="4576" heatid="7409" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.13" />
                    <SPLIT distance="100" swimtime="00:02:00.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4470" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="4525" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="4443" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4539" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" points="106" reactiontime="+77" swimtime="00:03:13.45" resultid="4577" heatid="7815" lane="4" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.50" />
                    <SPLIT distance="100" swimtime="00:01:50.37" />
                    <SPLIT distance="150" swimtime="00:02:27.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4565" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4539" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4533" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4525" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SMMK" name="Straż Miejska Miasta Kraków" nation="POL" region="MAL">
          <CONTACT city="Kraków" name="Jawień Krzysztof" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1971-06-11" firstname="Krzysztof" gender="M" lastname="Jawień" nation="POL" athleteid="4604">
              <RESULTS>
                <RESULT eventid="1109" points="342" reactiontime="+80" swimtime="00:02:37.33" resultid="4605" heatid="7400" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:01:57.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="342" reactiontime="+81" swimtime="00:02:52.45" resultid="4606" heatid="7472" lane="6" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                    <SPLIT distance="100" swimtime="00:01:21.56" />
                    <SPLIT distance="150" swimtime="00:02:06.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="260" reactiontime="+83" swimtime="00:02:50.91" resultid="4607" heatid="7569" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                    <SPLIT distance="150" swimtime="00:02:03.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="374" reactiontime="+82" swimtime="00:01:17.12" resultid="4608" heatid="7608" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="262" reactiontime="+73" swimtime="00:02:45.70" resultid="4610" heatid="7763" lane="3" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:18.46" />
                    <SPLIT distance="150" swimtime="00:02:02.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="365" reactiontime="+69" swimtime="00:00:35.32" resultid="4611" heatid="7806" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1559" points="296" reactiontime="+80" swimtime="00:05:53.36" resultid="8002" heatid="7979" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:02:04.19" />
                    <SPLIT distance="200" swimtime="00:02:52.63" />
                    <SPLIT distance="250" swimtime="00:03:41.16" />
                    <SPLIT distance="300" swimtime="00:04:30.28" />
                    <SPLIT distance="350" swimtime="00:05:11.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00315" name="Akwawit Astromal Leszno" nation="POL" region="PO">
          <CONTACT email="krzychutomczyk@o2.pl" name="Tomczyk Krzysztof" phone="723524682" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-14" firstname="Krzysztof" gender="M" lastname="Tomczyk" nation="POL" athleteid="4613">
              <RESULTS>
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="4614" heatid="7482" lane="4" entrytime="00:02:50.00" />
                <RESULT eventid="1402" points="439" reactiontime="+85" swimtime="00:01:13.12" resultid="4615" heatid="7608" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="445" swimtime="00:00:28.54" resultid="4616" heatid="7642" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1662" points="457" reactiontime="+80" swimtime="00:00:32.78" resultid="4617" heatid="7811" lane="6" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Tp Masters Opole" nation="POL">
          <CONTACT city="OPOLE" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="4619">
              <RESULTS>
                <RESULT eventid="1075" points="397" reactiontime="+78" swimtime="00:00:27.61" resultid="4620" heatid="7368" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="1200" points="358" reactiontime="+62" swimtime="00:00:31.82" resultid="4621" heatid="7453" lane="6" entrytime="00:00:33.50" />
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1268" status="DSQ" swimtime="00:01:00.02" resultid="4622" heatid="7521" lane="5" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="393" reactiontime="+77" swimtime="00:00:29.75" resultid="4623" heatid="7637" lane="3" entrytime="00:00:30.90" />
                <RESULT eventid="1470" points="371" reactiontime="+63" swimtime="00:01:08.08" resultid="4624" heatid="7671" lane="5" entrytime="00:01:08.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Grzegorz" gender="M" lastname="Radomski" nation="POL" athleteid="4625">
              <RESULTS>
                <RESULT eventid="1109" points="557" reactiontime="+76" swimtime="00:02:13.73" resultid="4626" heatid="7406" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                    <SPLIT distance="100" swimtime="00:01:01.74" />
                    <SPLIT distance="150" swimtime="00:01:40.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="467" reactiontime="+78" swimtime="00:18:15.10" resultid="4627" heatid="7916" lane="3" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                    <SPLIT distance="150" swimtime="00:01:40.59" />
                    <SPLIT distance="200" swimtime="00:02:16.15" />
                    <SPLIT distance="250" swimtime="00:02:51.80" />
                    <SPLIT distance="300" swimtime="00:03:27.82" />
                    <SPLIT distance="350" swimtime="00:04:03.93" />
                    <SPLIT distance="400" swimtime="00:04:40.07" />
                    <SPLIT distance="450" swimtime="00:05:16.10" />
                    <SPLIT distance="500" swimtime="00:05:52.71" />
                    <SPLIT distance="550" swimtime="00:06:29.11" />
                    <SPLIT distance="600" swimtime="00:07:05.60" />
                    <SPLIT distance="650" swimtime="00:07:41.49" />
                    <SPLIT distance="700" swimtime="00:08:17.98" />
                    <SPLIT distance="750" swimtime="00:08:54.44" />
                    <SPLIT distance="800" swimtime="00:09:31.23" />
                    <SPLIT distance="850" swimtime="00:10:07.81" />
                    <SPLIT distance="900" swimtime="00:10:45.23" />
                    <SPLIT distance="950" swimtime="00:11:22.29" />
                    <SPLIT distance="1000" swimtime="00:11:59.39" />
                    <SPLIT distance="1050" swimtime="00:12:36.38" />
                    <SPLIT distance="1100" swimtime="00:13:14.09" />
                    <SPLIT distance="1150" swimtime="00:13:51.49" />
                    <SPLIT distance="1200" swimtime="00:14:29.06" />
                    <SPLIT distance="1250" swimtime="00:15:06.75" />
                    <SPLIT distance="1300" swimtime="00:15:44.58" />
                    <SPLIT distance="1350" swimtime="00:16:22.24" />
                    <SPLIT distance="1400" swimtime="00:17:00.31" />
                    <SPLIT distance="1450" swimtime="00:17:38.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="534" reactiontime="+77" swimtime="00:04:50.19" resultid="4628" heatid="7977" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:43.84" />
                    <SPLIT distance="200" swimtime="00:02:20.45" />
                    <SPLIT distance="250" swimtime="00:03:00.26" />
                    <SPLIT distance="300" swimtime="00:03:41.35" />
                    <SPLIT distance="350" swimtime="00:04:16.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Jan" gender="M" lastname="Bryniak" nation="POL" athleteid="4629">
              <RESULTS>
                <RESULT eventid="1234" points="201" reactiontime="+114" swimtime="00:03:25.88" resultid="4630" heatid="7474" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                    <SPLIT distance="100" swimtime="00:01:37.68" />
                    <SPLIT distance="150" swimtime="00:02:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="139" reactiontime="+107" swimtime="00:03:30.20" resultid="4631" heatid="7567" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                    <SPLIT distance="100" swimtime="00:01:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="214" reactiontime="+122" swimtime="00:01:32.95" resultid="4632" heatid="7595" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="166" swimtime="00:07:07.70" resultid="4633" heatid="7976" lane="5" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                    <SPLIT distance="100" swimtime="00:01:38.98" />
                    <SPLIT distance="150" swimtime="00:02:35.59" />
                    <SPLIT distance="200" swimtime="00:03:34.38" />
                    <SPLIT distance="250" swimtime="00:04:30.11" />
                    <SPLIT distance="300" swimtime="00:05:27.25" />
                    <SPLIT distance="350" swimtime="00:06:18.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Oskar" gender="M" lastname="Orski" nation="POL" athleteid="4634">
              <RESULTS>
                <RESULT eventid="1075" points="329" reactiontime="+99" swimtime="00:00:29.39" resultid="4635" heatid="7367" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1268" points="302" reactiontime="+91" swimtime="00:01:06.97" resultid="4636" heatid="7512" lane="6" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Witkowski" nation="POL" athleteid="4637">
              <RESULTS>
                <RESULT eventid="1075" points="170" reactiontime="+119" swimtime="00:00:36.64" resultid="4638" heatid="7351" lane="4" entrytime="00:00:36.50" />
                <RESULT eventid="1109" points="62" reactiontime="+116" swimtime="00:04:37.19" resultid="4639" heatid="7391" lane="3" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.46" />
                    <SPLIT distance="100" swimtime="00:02:13.94" />
                    <SPLIT distance="150" swimtime="00:03:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="89" reactiontime="+85" swimtime="00:00:50.46" resultid="4640" heatid="7445" lane="5" entrytime="00:00:49.00" />
                <RESULT eventid="1268" points="122" reactiontime="+119" swimtime="00:01:30.47" resultid="4641" heatid="7503" lane="4" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="50" reactiontime="+116" swimtime="00:00:59.08" resultid="4642" heatid="7624" lane="2" entrytime="00:00:58.00" />
                <RESULT eventid="1470" points="77" reactiontime="+91" swimtime="00:01:54.86" resultid="4643" heatid="7662" lane="5" entrytime="00:01:51.00" />
                <RESULT eventid="1628" points="68" reactiontime="+86" swimtime="00:04:19.22" resultid="4644" heatid="7764" lane="1" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.17" />
                    <SPLIT distance="100" swimtime="00:02:05.01" />
                    <SPLIT distance="150" swimtime="00:03:14.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="4645" heatid="7791" lane="4" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Jerzy" gender="M" lastname="Minkiewicz" nation="POL" athleteid="4646">
              <RESULTS>
                <RESULT eventid="1075" points="280" reactiontime="+88" swimtime="00:00:31.00" resultid="4647" heatid="7361" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1268" points="262" reactiontime="+84" swimtime="00:01:10.17" resultid="4648" heatid="7511" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="227" reactiontime="+90" swimtime="00:01:23.12" resultid="4649" heatid="7544" lane="3" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="229" reactiontime="+85" swimtime="00:00:35.60" resultid="4650" heatid="7631" lane="2" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Zbigniew" gender="M" lastname="Krasnodębski" nation="POL" athleteid="4651">
              <RESULTS>
                <RESULT eventid="1402" points="207" reactiontime="+93" swimtime="00:01:33.92" resultid="4652" heatid="7598" lane="6" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="237" reactiontime="+59" swimtime="00:02:28.27" resultid="4653" heatid="7930" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:15.08" />
                    <SPLIT distance="150" swimtime="00:01:51.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4619" number="1" reactiontime="+59" />
                    <RELAYPOSITION athleteid="4651" number="2" />
                    <RELAYPOSITION athleteid="4646" number="3" />
                    <RELAYPOSITION athleteid="4637" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1528" points="362" reactiontime="+78" swimtime="00:01:53.28" resultid="4654" heatid="7713" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                    <SPLIT distance="100" swimtime="00:00:58.69" />
                    <SPLIT distance="150" swimtime="00:01:27.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4619" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4646" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4634" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="4625" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SOPMAST" name="Sopot Masters" nation="POL" region="POM">
          <CONTACT city="SOPOT" email="sopotmasters@o2.pl" internet="www.sopotmasters.pl" name="Gorbaczow Mirosław" phone="696 258 185" state="POMOR" street="ul. Haffnera 57" zip="81-715" />
          <ATHLETES>
            <ATHLETE birthdate="1958-12-28" firstname="Dariusz" gender="M" lastname="Gorbaczow" nation="POL" athleteid="4663">
              <RESULTS>
                <RESULT eventid="1200" points="314" reactiontime="+89" swimtime="00:00:33.25" resultid="4664" heatid="7451" lane="1" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1268" points="339" reactiontime="+85" swimtime="00:01:04.41" resultid="4665" heatid="7514" lane="2" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="344" swimtime="00:00:31.11" resultid="4666" heatid="7630" lane="5" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1470" points="260" reactiontime="+83" swimtime="00:01:16.59" resultid="4667" heatid="7667" lane="5" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="237" reactiontime="+82" swimtime="00:02:51.45" resultid="4668" heatid="7767" lane="6" entrytime="00:02:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.92" />
                    <SPLIT distance="100" swimtime="00:01:26.41" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STEEF" name="Steef Wrocław" nation="POL" region="DOL">
          <CONTACT city="Wrocław" email="ste1@wp.pl" name="Skrzypek Stefan" phone="500 388 374" street="Szewska 18" zip="50-139" />
          <ATHLETES>
            <ATHLETE birthdate="1978-02-26" firstname="Kuba" gender="M" lastname="Zwiernik" nation="POL" athleteid="4670">
              <RESULTS>
                <RESULT eventid="1075" points="273" reactiontime="+100" swimtime="00:00:31.26" resultid="4671" heatid="7369" lane="3" entrytime="00:00:28.05" />
                <RESULT eventid="1268" points="239" swimtime="00:01:12.33" resultid="4672" heatid="7512" lane="5" entrytime="00:01:07.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="208" swimtime="00:02:47.55" resultid="4673" heatid="7699" lane="5" entrytime="00:02:23.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:16.61" />
                    <SPLIT distance="150" swimtime="00:02:01.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-05-27" firstname="Krzysztof" gender="M" lastname="Nowak" nation="POL" athleteid="4674">
              <RESULTS>
                <RESULT eventid="1109" points="100" reactiontime="+112" swimtime="00:03:56.57" resultid="4675" heatid="7393" lane="1" entrytime="00:04:05.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.90" />
                    <SPLIT distance="100" swimtime="00:01:56.47" />
                    <SPLIT distance="150" swimtime="00:03:00.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="119" swimtime="00:04:04.70" resultid="4676" heatid="7473" lane="5" entrytime="00:03:58.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                    <SPLIT distance="100" swimtime="00:01:53.86" />
                    <SPLIT distance="150" swimtime="00:02:58.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="130" reactiontime="+115" swimtime="00:01:49.73" resultid="4677" heatid="7595" lane="1" entrytime="00:01:50.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="146" swimtime="00:00:47.90" resultid="4678" heatid="7792" lane="5" entrytime="00:00:49.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="4679">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski 50 motylkowym." eventid="1092" points="343" reactiontime="+94" swimtime="00:02:57.90" resultid="4680" heatid="7388" lane="6" entrytime="00:02:55.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:23.60" />
                    <SPLIT distance="150" swimtime="00:02:15.74" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1148" points="317" swimtime="00:11:49.91" resultid="4681" heatid="7904" lane="5" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:26.40" />
                    <SPLIT distance="150" swimtime="00:02:12.17" />
                    <SPLIT distance="200" swimtime="00:02:58.77" />
                    <SPLIT distance="250" swimtime="00:03:44.58" />
                    <SPLIT distance="300" swimtime="00:04:30.41" />
                    <SPLIT distance="350" swimtime="00:05:15.84" />
                    <SPLIT distance="400" swimtime="00:06:01.21" />
                    <SPLIT distance="450" swimtime="00:06:44.91" />
                    <SPLIT distance="500" swimtime="00:07:30.05" />
                    <SPLIT distance="550" swimtime="00:08:14.29" />
                    <SPLIT distance="600" swimtime="00:08:58.70" />
                    <SPLIT distance="650" swimtime="00:09:42.09" />
                    <SPLIT distance="700" swimtime="00:10:26.03" />
                    <SPLIT distance="750" swimtime="00:11:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="252" reactiontime="+95" swimtime="00:00:40.64" resultid="4682" heatid="7437" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1251" points="296" reactiontime="+91" swimtime="00:01:16.50" resultid="4683" heatid="7494" lane="4" entrytime="00:01:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="285" reactiontime="+89" swimtime="00:01:23.84" resultid="4684" heatid="7655" lane="5" entrytime="00:01:21.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="296" reactiontime="+102" swimtime="00:06:31.68" resultid="4685" heatid="7718" lane="6" entrytime="00:06:24.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                    <SPLIT distance="100" swimtime="00:01:34.18" />
                    <SPLIT distance="150" swimtime="00:02:23.31" />
                    <SPLIT distance="200" swimtime="00:03:11.58" />
                    <SPLIT distance="250" swimtime="00:04:07.42" />
                    <SPLIT distance="300" swimtime="00:05:03.64" />
                    <SPLIT distance="350" swimtime="00:05:48.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="300" reactiontime="+88" swimtime="00:02:59.28" resultid="4686" heatid="7759" lane="3" entrytime="00:02:55.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                    <SPLIT distance="100" swimtime="00:01:28.03" />
                    <SPLIT distance="150" swimtime="00:02:13.85" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1693" points="318" swimtime="00:05:43.84" resultid="4687" heatid="8022" lane="5" entrytime="00:05:56.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                    <SPLIT distance="150" swimtime="00:02:05.36" />
                    <SPLIT distance="200" swimtime="00:02:49.10" />
                    <SPLIT distance="250" swimtime="00:03:32.97" />
                    <SPLIT distance="300" swimtime="00:04:17.39" />
                    <SPLIT distance="350" swimtime="00:05:01.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="4688">
              <RESULTS>
                <RESULT eventid="1075" points="209" reactiontime="+96" swimtime="00:00:34.17" resultid="4689" heatid="7355" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1165" points="208" reactiontime="+106" swimtime="00:23:54.66" resultid="4690" heatid="7910" lane="4" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:24.19" />
                    <SPLIT distance="150" swimtime="00:02:09.40" />
                    <SPLIT distance="200" swimtime="00:02:55.51" />
                    <SPLIT distance="250" swimtime="00:03:42.01" />
                    <SPLIT distance="300" swimtime="00:04:28.82" />
                    <SPLIT distance="350" swimtime="00:05:16.29" />
                    <SPLIT distance="400" swimtime="00:06:03.86" />
                    <SPLIT distance="450" swimtime="00:06:51.42" />
                    <SPLIT distance="500" swimtime="00:07:38.64" />
                    <SPLIT distance="550" swimtime="00:08:25.67" />
                    <SPLIT distance="600" swimtime="00:09:13.42" />
                    <SPLIT distance="650" swimtime="00:10:01.57" />
                    <SPLIT distance="700" swimtime="00:10:50.70" />
                    <SPLIT distance="750" swimtime="00:11:40.30" />
                    <SPLIT distance="800" swimtime="00:12:29.48" />
                    <SPLIT distance="850" swimtime="00:13:18.37" />
                    <SPLIT distance="900" swimtime="00:14:07.31" />
                    <SPLIT distance="950" swimtime="00:14:56.80" />
                    <SPLIT distance="1000" swimtime="00:15:46.41" />
                    <SPLIT distance="1050" swimtime="00:16:35.42" />
                    <SPLIT distance="1100" swimtime="00:17:24.52" />
                    <SPLIT distance="1150" swimtime="00:18:14.40" />
                    <SPLIT distance="1200" swimtime="00:19:03.22" />
                    <SPLIT distance="1250" swimtime="00:19:51.76" />
                    <SPLIT distance="1300" swimtime="00:20:41.19" />
                    <SPLIT distance="1350" swimtime="00:21:29.41" />
                    <SPLIT distance="1400" swimtime="00:22:18.02" />
                    <SPLIT distance="1450" swimtime="00:23:07.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="4691" heatid="7448" lane="4" entrytime="00:00:37.50" />
                <RESULT eventid="1336" points="148" reactiontime="+104" swimtime="00:03:26.19" resultid="4692" heatid="7567" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                    <SPLIT distance="100" swimtime="00:01:38.14" />
                    <SPLIT distance="150" swimtime="00:02:34.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="4693" heatid="7629" lane="6" entrytime="00:00:37.65" />
                <RESULT eventid="1504" points="225" reactiontime="+96" swimtime="00:02:43.22" resultid="4694" heatid="7692" lane="2" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:19.22" />
                    <SPLIT distance="150" swimtime="00:02:00.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="4695" heatid="7797" lane="4" entrytime="00:00:40.50" />
                <RESULT eventid="1710" points="228" swimtime="00:05:48.10" resultid="4696" heatid="8050" lane="5" entrytime="00:05:54.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:23.37" />
                    <SPLIT distance="150" swimtime="00:02:06.87" />
                    <SPLIT distance="200" swimtime="00:02:50.94" />
                    <SPLIT distance="250" swimtime="00:03:35.03" />
                    <SPLIT distance="300" swimtime="00:04:19.20" />
                    <SPLIT distance="350" swimtime="00:05:03.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Weteran  Zabrze" nation="POL">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW.JANA  4A/4" zip="41803" />
          <ATHLETES>
            <ATHLETE birthdate="1951-02-18" firstname="Genowefa" gender="F" lastname="Drużyńska" nation="POL" athleteid="4698">
              <RESULTS>
                <RESULT eventid="1385" points="122" swimtime="00:02:06.24" resultid="4699" heatid="7583" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="131" reactiontime="+94" swimtime="00:00:56.68" resultid="4700" heatid="7777" lane="4" entrytime="00:00:57.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-23" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" license="502611100004" athleteid="4701">
              <RESULTS>
                <RESULT eventid="1058" points="121" reactiontime="+94" swimtime="00:00:46.95" resultid="4702" heatid="7334" lane="6" entrytime="00:00:47.00" />
                <RESULT eventid="1183" points="99" reactiontime="+75" swimtime="00:00:55.43" resultid="4703" heatid="7431" lane="3" />
                <RESULT eventid="1453" points="75" reactiontime="+79" swimtime="00:02:10.55" resultid="4704" heatid="7648" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="4705" heatid="7753" lane="2" />
                <RESULT eventid="1645" points="173" swimtime="00:00:51.67" resultid="4706" heatid="7778" lane="5" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" license="502611200004" athleteid="4707">
              <RESULTS>
                <RESULT eventid="1200" points="150" reactiontime="+66" swimtime="00:00:42.52" resultid="4708" heatid="7446" lane="5" entrytime="00:00:42.54" />
                <RESULT eventid="1470" points="127" reactiontime="+67" swimtime="00:01:37.25" resultid="4709" heatid="7663" lane="6" entrytime="00:01:37.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="113" reactiontime="+63" swimtime="00:03:39.30" resultid="4710" heatid="7764" lane="4" entrytime="00:03:41.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.47" />
                    <SPLIT distance="100" swimtime="00:01:44.27" />
                    <SPLIT distance="150" swimtime="00:02:41.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="502611100009" athleteid="4711">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="4712" heatid="7389" lane="6" entrytime="00:02:45.00" />
                <RESULT eventid="1148" points="482" swimtime="00:10:17.72" resultid="4713" heatid="7906" lane="5" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:12.13" />
                    <SPLIT distance="150" swimtime="00:01:50.38" />
                    <SPLIT distance="200" swimtime="00:02:28.87" />
                    <SPLIT distance="250" swimtime="00:03:07.94" />
                    <SPLIT distance="300" swimtime="00:03:47.19" />
                    <SPLIT distance="350" swimtime="00:04:26.37" />
                    <SPLIT distance="400" swimtime="00:05:05.68" />
                    <SPLIT distance="450" swimtime="00:05:44.85" />
                    <SPLIT distance="500" swimtime="00:06:23.91" />
                    <SPLIT distance="550" swimtime="00:07:03.18" />
                    <SPLIT distance="600" swimtime="00:07:42.53" />
                    <SPLIT distance="650" swimtime="00:08:22.02" />
                    <SPLIT distance="700" swimtime="00:09:01.02" />
                    <SPLIT distance="750" swimtime="00:09:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1217" points="428" reactiontime="+92" swimtime="00:02:58.56" resultid="4714" heatid="7469" lane="1" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:24.94" />
                    <SPLIT distance="150" swimtime="00:02:11.11" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1385" points="440" reactiontime="+89" swimtime="00:01:22.40" resultid="4715" heatid="7591" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1542" points="457" reactiontime="+90" swimtime="00:05:38.73" resultid="4716" heatid="7718" lane="4" entrytime="00:05:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:15.30" />
                    <SPLIT distance="150" swimtime="00:02:01.97" />
                    <SPLIT distance="200" swimtime="00:02:47.45" />
                    <SPLIT distance="250" swimtime="00:03:34.08" />
                    <SPLIT distance="300" swimtime="00:04:21.31" />
                    <SPLIT distance="350" swimtime="00:05:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1693" points="472" reactiontime="+94" swimtime="00:05:01.56" resultid="4717" heatid="8025" lane="1" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                    <SPLIT distance="150" swimtime="00:01:49.65" />
                    <SPLIT distance="200" swimtime="00:02:27.99" />
                    <SPLIT distance="250" swimtime="00:03:06.66" />
                    <SPLIT distance="300" swimtime="00:03:45.57" />
                    <SPLIT distance="350" swimtime="00:04:24.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-09" firstname="Anna" gender="F" lastname="Karlsson" nation="POL" license="502611100011" athleteid="4718">
              <RESULTS>
                <RESULT eventid="1058" points="352" reactiontime="+86" swimtime="00:00:32.92" resultid="4719" heatid="7340" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1251" points="295" reactiontime="+91" swimtime="00:01:16.61" resultid="4720" heatid="7492" lane="1" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-05-27" firstname="Dawid" gender="M" lastname="Muszala" nation="POL" athleteid="4721">
              <RESULTS>
                <RESULT eventid="1504" points="194" reactiontime="+74" swimtime="00:02:51.52" resultid="4723" heatid="7692" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:21.99" />
                    <SPLIT distance="150" swimtime="00:02:05.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="199" swimtime="00:06:03.90" resultid="4724" heatid="8049" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:01:22.18" />
                    <SPLIT distance="150" swimtime="00:02:08.96" />
                    <SPLIT distance="200" swimtime="00:02:56.59" />
                    <SPLIT distance="250" swimtime="00:03:44.63" />
                    <SPLIT distance="300" swimtime="00:04:33.39" />
                    <SPLIT distance="350" swimtime="00:05:21.48" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Przekroczony limit czasu." eventid="1165" reactiontime="+76" status="DSQ" swimtime="00:25:03.36" resultid="7927" heatid="7907" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:21.29" />
                    <SPLIT distance="150" swimtime="00:02:06.14" />
                    <SPLIT distance="200" swimtime="00:02:58.13" />
                    <SPLIT distance="250" swimtime="00:03:46.56" />
                    <SPLIT distance="300" swimtime="00:04:36.06" />
                    <SPLIT distance="350" swimtime="00:05:27.40" />
                    <SPLIT distance="400" swimtime="00:06:19.46" />
                    <SPLIT distance="450" swimtime="00:07:11.26" />
                    <SPLIT distance="500" swimtime="00:08:03.50" />
                    <SPLIT distance="550" swimtime="00:08:54.47" />
                    <SPLIT distance="600" swimtime="00:09:44.53" />
                    <SPLIT distance="650" swimtime="00:10:34.58" />
                    <SPLIT distance="700" swimtime="00:11:25.38" />
                    <SPLIT distance="750" swimtime="00:12:17.37" />
                    <SPLIT distance="800" swimtime="00:13:09.23" />
                    <SPLIT distance="850" swimtime="00:14:02.42" />
                    <SPLIT distance="900" swimtime="00:14:53.86" />
                    <SPLIT distance="950" swimtime="00:15:44.66" />
                    <SPLIT distance="1000" swimtime="00:16:36.15" />
                    <SPLIT distance="1050" swimtime="00:17:27.25" />
                    <SPLIT distance="1100" swimtime="00:18:19.02" />
                    <SPLIT distance="1150" swimtime="00:19:10.03" />
                    <SPLIT distance="1200" swimtime="00:19:59.90" />
                    <SPLIT distance="1250" swimtime="00:20:52.65" />
                    <SPLIT distance="1300" swimtime="00:21:45.31" />
                    <SPLIT distance="1350" swimtime="00:22:37.46" />
                    <SPLIT distance="1400" swimtime="00:23:28.21" />
                    <SPLIT distance="1450" swimtime="00:24:19.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="502611100001" athleteid="4725">
              <RESULTS>
                <RESULT eventid="1058" points="272" reactiontime="+85" swimtime="00:00:35.85" resultid="4726" heatid="7337" lane="4" entrytime="00:00:36.78" />
                <RESULT eventid="1183" points="191" reactiontime="+69" swimtime="00:00:44.62" resultid="4727" heatid="7434" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1251" points="226" reactiontime="+81" swimtime="00:01:23.72" resultid="4728" heatid="7491" lane="6" entrytime="00:01:24.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="164" reactiontime="+65" swimtime="00:01:40.71" resultid="4729" heatid="7651" lane="2" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="502611200002" athleteid="4730">
              <RESULTS>
                <RESULT eventid="1234" points="179" swimtime="00:03:33.93" resultid="4731" heatid="7474" lane="5" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.77" />
                    <SPLIT distance="100" swimtime="00:01:43.57" />
                    <SPLIT distance="150" swimtime="00:02:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="182" reactiontime="+100" swimtime="00:01:38.09" resultid="4732" heatid="7597" lane="2" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="168" reactiontime="+96" swimtime="00:00:45.76" resultid="4733" heatid="7794" lane="4" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="502611100002" athleteid="4734">
              <RESULTS>
                <RESULT eventid="1148" points="114" reactiontime="+110" swimtime="00:16:38.66" resultid="4735" heatid="7902" lane="4" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.62" />
                    <SPLIT distance="100" swimtime="00:01:54.20" />
                    <SPLIT distance="150" swimtime="00:02:56.47" />
                    <SPLIT distance="200" swimtime="00:03:58.79" />
                    <SPLIT distance="250" swimtime="00:05:01.84" />
                    <SPLIT distance="300" swimtime="00:06:05.45" />
                    <SPLIT distance="350" swimtime="00:07:08.49" />
                    <SPLIT distance="400" swimtime="00:08:11.22" />
                    <SPLIT distance="450" swimtime="00:09:14.26" />
                    <SPLIT distance="500" swimtime="00:10:18.56" />
                    <SPLIT distance="550" swimtime="00:11:21.33" />
                    <SPLIT distance="600" swimtime="00:12:23.64" />
                    <SPLIT distance="650" swimtime="00:13:28.20" />
                    <SPLIT distance="700" swimtime="00:14:30.87" />
                    <SPLIT distance="750" swimtime="00:15:36.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="163" swimtime="00:04:05.91" resultid="4736" heatid="7464" lane="5" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.93" />
                    <SPLIT distance="100" swimtime="00:02:00.39" />
                    <SPLIT distance="150" swimtime="00:03:03.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="163" reactiontime="+106" swimtime="00:01:54.57" resultid="4737" heatid="7584" lane="4" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="168" reactiontime="+108" swimtime="00:00:52.19" resultid="4738" heatid="7778" lane="2" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-28" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="502611200007" athleteid="4739">
              <RESULTS>
                <RESULT eventid="1075" points="261" reactiontime="+83" swimtime="00:00:31.74" resultid="4740" heatid="7358" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1302" points="169" reactiontime="+90" swimtime="00:01:31.79" resultid="4741" heatid="7542" lane="2" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="241" reactiontime="+84" swimtime="00:00:35.03" resultid="4742" heatid="7631" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-05" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" license="502611100005" athleteid="4743">
              <RESULTS>
                <RESULT eventid="1058" points="186" reactiontime="+95" swimtime="00:00:40.66" resultid="4744" heatid="7335" lane="6" entrytime="00:00:40.30" />
                <RESULT eventid="1251" points="172" reactiontime="+91" swimtime="00:01:31.70" resultid="4745" heatid="7489" lane="3" entrytime="00:01:33.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="126" reactiontime="+98" swimtime="00:03:41.73" resultid="4746" heatid="7676" lane="4" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.24" />
                    <SPLIT distance="100" swimtime="00:01:43.26" />
                    <SPLIT distance="150" swimtime="00:02:42.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="502611200008" athleteid="4747">
              <RESULTS>
                <RESULT eventid="1075" points="269" reactiontime="+85" swimtime="00:00:31.41" resultid="4748" heatid="7360" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1200" points="194" reactiontime="+67" swimtime="00:00:39.01" resultid="4749" heatid="7447" lane="3" entrytime="00:00:39.30" />
                <RESULT eventid="1470" points="156" reactiontime="+72" swimtime="00:01:30.89" resultid="4750" heatid="7664" lane="6" entrytime="00:01:28.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" reactiontime="+58" status="DNF" swimtime="00:00:00.00" resultid="4751" heatid="7766" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:31.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-04" firstname="Ulasz" gender="M" lastname="Szanli" nation="POL" license="502611200015" athleteid="4752">
              <RESULTS>
                <RESULT eventid="1075" points="207" reactiontime="+92" swimtime="00:00:34.27" resultid="4753" heatid="7352" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1268" points="131" reactiontime="+104" swimtime="00:01:28.45" resultid="4754" heatid="7502" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-14" firstname="Maciej" gender="M" lastname="Kunicki" nation="POL" license="502611200011" athleteid="4755">
              <RESULTS>
                <RESULT eventid="1336" points="240" reactiontime="+89" swimtime="00:02:55.41" resultid="4756" heatid="7569" lane="1" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:21.89" />
                    <SPLIT distance="150" swimtime="00:02:08.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="324" reactiontime="+89" swimtime="00:00:31.72" resultid="4757" heatid="7634" lane="1" entrytime="00:00:32.50" />
                <RESULT eventid="1594" points="288" reactiontime="+83" swimtime="00:01:13.40" resultid="4758" heatid="7746" lane="2" entrytime="00:01:12.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="502611200005" athleteid="4759">
              <RESULTS>
                <RESULT eventid="1075" points="131" reactiontime="+108" swimtime="00:00:39.90" resultid="4760" heatid="7351" lane="1" entrytime="00:00:37.50" />
                <RESULT eventid="1200" points="82" reactiontime="+91" swimtime="00:00:51.84" resultid="4761" heatid="7444" lane="6" entrytime="00:00:55.45" />
                <RESULT eventid="1302" points="88" reactiontime="+104" swimtime="00:01:53.96" resultid="4762" heatid="7540" lane="4" entrytime="00:01:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="92" reactiontime="+101" swimtime="00:00:48.14" resultid="4763" heatid="7626" lane="2" entrytime="00:00:42.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1377" points="189" reactiontime="+73" swimtime="00:02:39.77" resultid="4767" heatid="7930" lane="1" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:24.40" />
                    <SPLIT distance="150" swimtime="00:02:01.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4747" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4730" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4739" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="4759" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1528" points="202" reactiontime="+91" swimtime="00:02:17.58" resultid="4769" heatid="7711" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:15.74" />
                    <SPLIT distance="150" swimtime="00:01:47.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4707" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="4759" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="4739" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4755" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1370" points="218" reactiontime="+66" swimtime="00:02:50.59" resultid="4766" heatid="7572" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                    <SPLIT distance="100" swimtime="00:01:36.76" />
                    <SPLIT distance="150" swimtime="00:02:11.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4725" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4734" number="2" />
                    <RELAYPOSITION athleteid="4711" number="3" />
                    <RELAYPOSITION athleteid="4743" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="1521" points="201" reactiontime="+79" swimtime="00:02:39.04" resultid="4768" heatid="7707" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:25.47" />
                    <SPLIT distance="150" swimtime="00:02:07.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4725" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4701" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="4743" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4711" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="319" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1126" points="128" reactiontime="+80" swimtime="00:02:40.08" resultid="6439" heatid="7409" lane="6" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:25.63" />
                    <SPLIT distance="150" swimtime="00:02:05.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4725" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4734" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4730" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4739" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="1679" points="211" reactiontime="+68" swimtime="00:02:34.08" resultid="4765" heatid="7815" lane="1" entrytime="00:02:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:01:21.90" />
                    <SPLIT distance="150" swimtime="00:01:57.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4707" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4711" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4739" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="4725" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" name="MOTYL -SENIOR MOSiR Stalowa Wola" nation="POL" region="PDK" shortname="MOTYL -SENIOR MOSiR Stalowa Wo">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" state="PDK" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="4784">
              <RESULTS>
                <RESULT eventid="1075" points="451" swimtime="00:00:26.47" resultid="4785" heatid="7377" lane="5" entrytime="00:00:26.07" />
                <RESULT eventid="1109" points="394" reactiontime="+96" swimtime="00:02:30.03" resultid="4786" heatid="7405" lane="1" entrytime="00:02:27.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:09.38" />
                    <SPLIT distance="150" swimtime="00:01:54.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="425" reactiontime="+73" swimtime="00:00:30.06" resultid="4787" heatid="7458" lane="6" entrytime="00:00:29.96" />
                <RESULT eventid="1268" points="443" reactiontime="+85" swimtime="00:00:58.94" resultid="4788" heatid="7523" lane="4" entrytime="00:00:57.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="404" reactiontime="+84" swimtime="00:00:29.48" resultid="4789" heatid="7638" lane="1" entrytime="00:00:30.66" />
                <RESULT eventid="1470" points="408" reactiontime="+79" swimtime="00:01:05.98" resultid="4790" heatid="7672" lane="4" entrytime="00:01:05.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="388" reactiontime="+73" swimtime="00:02:25.47" resultid="4791" heatid="7773" lane="1" entrytime="00:02:26.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:11.15" />
                    <SPLIT distance="150" swimtime="00:01:48.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="346" reactiontime="+89" swimtime="00:00:35.96" resultid="4792" heatid="7804" lane="2" entrytime="00:00:36.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="4793">
              <RESULTS>
                <RESULT eventid="1075" points="479" swimtime="00:00:25.93" resultid="4794" heatid="7349" lane="5" entrytime="00:00:41.99" />
                <RESULT eventid="1109" points="526" reactiontime="+71" swimtime="00:02:16.30" resultid="4795" heatid="7407" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                    <SPLIT distance="100" swimtime="00:01:04.55" />
                    <SPLIT distance="150" swimtime="00:01:44.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="520" reactiontime="+66" swimtime="00:00:55.87" resultid="4796" heatid="7524" lane="6" entrytime="00:00:56.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="520" reactiontime="+74" swimtime="00:01:03.12" resultid="4797" heatid="7559" lane="2" entrytime="00:01:03.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="512" reactiontime="+76" swimtime="00:00:27.24" resultid="4798" heatid="7645" lane="4" entrytime="00:00:27.29" />
                <RESULT eventid="1504" points="512" reactiontime="+75" swimtime="00:02:04.19" resultid="4799" heatid="7705" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                    <SPLIT distance="100" swimtime="00:01:00.90" />
                    <SPLIT distance="150" swimtime="00:01:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="530" reactiontime="+74" swimtime="00:00:59.89" resultid="4800" heatid="7752" lane="1" entrytime="00:00:59.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="408" reactiontime="+71" swimtime="00:02:23.01" resultid="4801" heatid="7773" lane="2" entrytime="00:02:22.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:09.69" />
                    <SPLIT distance="150" swimtime="00:01:46.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-06-01" firstname="Arkadiusz" gender="M" lastname="Janik" nation="POL" athleteid="4802">
              <RESULTS>
                <RESULT eventid="1075" points="315" reactiontime="+85" swimtime="00:00:29.81" resultid="4803" heatid="7365" lane="4" entrytime="00:00:29.51" />
                <RESULT eventid="1165" points="241" reactiontime="+90" swimtime="00:22:44.87" resultid="4804" heatid="7911" lane="2" entrytime="00:24:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:23.97" />
                    <SPLIT distance="150" swimtime="00:02:08.71" />
                    <SPLIT distance="200" swimtime="00:02:54.39" />
                    <SPLIT distance="250" swimtime="00:03:39.50" />
                    <SPLIT distance="300" swimtime="00:04:25.47" />
                    <SPLIT distance="350" swimtime="00:07:28.98" />
                    <SPLIT distance="400" swimtime="00:08:16.07" />
                    <SPLIT distance="450" swimtime="00:09:02.16" />
                    <SPLIT distance="500" swimtime="00:09:48.04" />
                    <SPLIT distance="550" swimtime="00:10:33.78" />
                    <SPLIT distance="600" swimtime="00:11:19.81" />
                    <SPLIT distance="650" swimtime="00:12:06.27" />
                    <SPLIT distance="700" swimtime="00:12:53.03" />
                    <SPLIT distance="750" swimtime="00:13:38.79" />
                    <SPLIT distance="800" swimtime="00:14:25.12" />
                    <SPLIT distance="850" swimtime="00:15:11.03" />
                    <SPLIT distance="900" swimtime="00:16:42.87" />
                    <SPLIT distance="950" swimtime="00:18:14.82" />
                    <SPLIT distance="1000" swimtime="00:20:32.93" />
                    <SPLIT distance="1050" swimtime="00:22:02.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="296" reactiontime="+86" swimtime="00:01:07.38" resultid="4805" heatid="7512" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="271" swimtime="00:01:18.42" resultid="4806" heatid="7546" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="282" reactiontime="+89" swimtime="00:00:33.23" resultid="4807" heatid="7633" lane="6" entrytime="00:00:33.50" />
                <RESULT eventid="1504" points="249" reactiontime="+88" swimtime="00:02:37.84" resultid="4808" heatid="7697" lane="1" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="150" swimtime="00:01:57.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="162" reactiontime="+89" swimtime="00:01:28.88" resultid="4809" heatid="7743" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="4810" heatid="8052" lane="4" entrytime="00:05:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzinierz" gender="M" lastname="Jarzyna" nation="POL" athleteid="4811">
              <RESULTS>
                <RESULT eventid="1075" points="236" reactiontime="+87" swimtime="00:00:32.81" resultid="4812" heatid="7355" lane="4" entrytime="00:00:33.49" />
                <RESULT eventid="1109" points="153" reactiontime="+92" swimtime="00:03:25.41" resultid="4813" heatid="7395" lane="2" entrytime="00:03:22.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.48" />
                    <SPLIT distance="100" swimtime="00:01:38.04" />
                    <SPLIT distance="150" swimtime="00:02:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="146" reactiontime="+67" swimtime="00:00:42.88" resultid="4814" heatid="7446" lane="6" entrytime="00:00:43.41" />
                <RESULT eventid="1302" points="171" swimtime="00:01:31.31" resultid="4815" heatid="7542" lane="5" entrytime="00:01:34.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="144" reactiontime="+82" swimtime="00:01:33.26" resultid="4816" heatid="7663" lane="5" entrytime="00:01:33.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="149" reactiontime="+101" swimtime="00:07:23.37" resultid="4817" heatid="7977" lane="1" entrytime="00:07:24.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.44" />
                    <SPLIT distance="100" swimtime="00:01:53.07" />
                    <SPLIT distance="150" swimtime="00:03:42.85" />
                    <SPLIT distance="200" swimtime="00:04:45.67" />
                    <SPLIT distance="250" swimtime="00:05:47.61" />
                    <SPLIT distance="300" swimtime="00:06:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="141" reactiontime="+73" swimtime="00:03:23.51" resultid="4818" heatid="7765" lane="2" entrytime="00:03:28.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.71" />
                    <SPLIT distance="100" swimtime="00:01:40.22" />
                    <SPLIT distance="150" swimtime="00:02:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="168" reactiontime="+102" swimtime="00:06:24.87" resultid="4819" heatid="8047" lane="2" entrytime="00:06:27.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:30.60" />
                    <SPLIT distance="150" swimtime="00:02:20.81" />
                    <SPLIT distance="200" swimtime="00:03:11.54" />
                    <SPLIT distance="250" swimtime="00:04:02.13" />
                    <SPLIT distance="300" swimtime="00:04:52.68" />
                    <SPLIT distance="350" swimtime="00:05:40.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-18" firstname="Waldemar" gender="M" lastname="Kalbarczyk" nation="POL" athleteid="4820">
              <RESULTS>
                <RESULT eventid="1075" points="301" reactiontime="+90" swimtime="00:00:30.29" resultid="4821" heatid="7362" lane="6" entrytime="00:00:30.32" />
                <RESULT eventid="1109" points="269" reactiontime="+93" swimtime="00:02:50.41" resultid="4822" heatid="7397" lane="3" entrytime="00:02:55.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:02:10.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="290" reactiontime="+91" swimtime="00:01:07.84" resultid="4823" heatid="7510" lane="4" entrytime="00:01:09.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="271" swimtime="00:01:18.40" resultid="4824" heatid="7547" lane="5" entrytime="00:01:18.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="276" reactiontime="+91" swimtime="00:00:33.45" resultid="4825" heatid="7632" lane="1" entrytime="00:00:34.50" />
                <RESULT eventid="1470" points="223" reactiontime="+83" swimtime="00:01:20.64" resultid="4826" heatid="7665" lane="6" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="212" reactiontime="+99" swimtime="00:01:21.22" resultid="4827" heatid="7743" lane="1" entrytime="00:01:21.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="235" swimtime="00:02:51.93" resultid="4828" heatid="7767" lane="2" entrytime="00:02:56.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:02:08.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="4829">
              <RESULTS>
                <RESULT eventid="1075" points="303" reactiontime="+94" swimtime="00:00:30.22" resultid="4830" heatid="7361" lane="3" entrytime="00:00:30.41" />
                <RESULT eventid="1109" points="282" reactiontime="+90" swimtime="00:02:47.72" resultid="4831" heatid="7398" lane="4" entrytime="00:02:51.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                    <SPLIT distance="150" swimtime="00:02:09.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="307" reactiontime="+86" swimtime="00:01:06.61" resultid="4832" heatid="7512" lane="2" entrytime="00:01:07.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="196" reactiontime="+93" swimtime="00:03:07.67" resultid="4833" heatid="7568" lane="3" entrytime="00:03:07.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:24.21" />
                    <SPLIT distance="150" swimtime="00:02:13.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="4834" heatid="7665" lane="5" entrytime="00:01:21.30" />
                <RESULT eventid="1559" points="269" reactiontime="+98" swimtime="00:06:04.57" resultid="4835" heatid="7979" lane="4" entrytime="00:06:05.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:24.21" />
                    <SPLIT distance="150" swimtime="00:02:09.80" />
                    <SPLIT distance="200" swimtime="00:02:54.93" />
                    <SPLIT distance="250" swimtime="00:03:49.36" />
                    <SPLIT distance="300" swimtime="00:04:42.98" />
                    <SPLIT distance="350" swimtime="00:05:24.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="234" reactiontime="+91" swimtime="00:01:18.64" resultid="4836" heatid="7742" lane="4" entrytime="00:01:22.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="236" reactiontime="+91" swimtime="00:02:51.50" resultid="4837" heatid="7768" lane="1" entrytime="00:02:51.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:01:22.33" />
                    <SPLIT distance="150" swimtime="00:02:07.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="4838">
              <RESULTS>
                <RESULT eventid="1109" points="308" reactiontime="+82" swimtime="00:02:42.83" resultid="4839" heatid="7400" lane="4" entrytime="00:02:44.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:17.46" />
                    <SPLIT distance="150" swimtime="00:02:04.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="311" reactiontime="+86" swimtime="00:02:57.93" resultid="4841" heatid="7479" lane="6" entrytime="00:03:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:24.53" />
                    <SPLIT distance="150" swimtime="00:02:11.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="196" reactiontime="+90" swimtime="00:03:07.56" resultid="4842" heatid="7567" lane="2" entrytime="00:03:27.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                    <SPLIT distance="100" swimtime="00:01:27.54" />
                    <SPLIT distance="150" swimtime="00:02:17.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="333" swimtime="00:01:20.17" resultid="4843" heatid="7605" lane="5" entrytime="00:01:21.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="271" reactiontime="+88" swimtime="00:06:03.57" resultid="4844" heatid="7979" lane="2" entrytime="00:06:05.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                    <SPLIT distance="100" swimtime="00:01:28.66" />
                    <SPLIT distance="150" swimtime="00:02:16.13" />
                    <SPLIT distance="200" swimtime="00:03:02.05" />
                    <SPLIT distance="250" swimtime="00:03:52.51" />
                    <SPLIT distance="300" swimtime="00:04:42.61" />
                    <SPLIT distance="350" swimtime="00:05:24.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="257" reactiontime="+82" swimtime="00:02:46.89" resultid="4845" heatid="7769" lane="4" entrytime="00:02:44.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:20.89" />
                    <SPLIT distance="150" swimtime="00:02:04.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="351" reactiontime="+79" swimtime="00:00:35.77" resultid="4846" heatid="7804" lane="3" entrytime="00:00:36.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="4847">
              <RESULTS>
                <RESULT eventid="1058" points="292" reactiontime="+74" swimtime="00:00:35.01" resultid="4848" heatid="7338" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1092" points="277" reactiontime="+84" swimtime="00:03:11.02" resultid="4849" heatid="7385" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                    <SPLIT distance="100" swimtime="00:01:33.30" />
                    <SPLIT distance="150" swimtime="00:02:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="272" swimtime="00:03:27.53" resultid="4850" heatid="7466" lane="5" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                    <SPLIT distance="100" swimtime="00:01:41.01" />
                    <SPLIT distance="150" swimtime="00:02:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="190" reactiontime="+94" swimtime="00:03:29.74" resultid="4851" heatid="7562" lane="2" entrytime="00:03:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.60" />
                    <SPLIT distance="100" swimtime="00:01:39.37" />
                    <SPLIT distance="150" swimtime="00:02:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="246" reactiontime="+94" swimtime="00:01:40.00" resultid="4852" heatid="7587" lane="6" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="264" swimtime="00:00:37.99" resultid="4853" heatid="7616" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1577" points="210" reactiontime="+91" swimtime="00:01:32.51" resultid="4854" heatid="7732" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="259" reactiontime="+85" swimtime="00:00:45.17" resultid="4855" heatid="7782" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-12" firstname="Adam" gender="M" lastname="Przybylski" nation="POL" athleteid="4856">
              <RESULTS>
                <RESULT eventid="1075" points="395" reactiontime="+79" swimtime="00:00:27.65" resultid="4857" heatid="7372" lane="3" entrytime="00:00:27.44" />
                <RESULT eventid="1109" points="285" reactiontime="+73" swimtime="00:02:47.21" resultid="4858" heatid="7398" lane="3" entrytime="00:02:50.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:02:09.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="281" reactiontime="+66" swimtime="00:00:34.51" resultid="4859" heatid="7451" lane="5" entrytime="00:00:34.95" />
                <RESULT eventid="1268" points="376" swimtime="00:01:02.24" resultid="4860" heatid="7518" lane="5" entrytime="00:01:02.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="324" reactiontime="+84" swimtime="00:00:31.73" resultid="4861" heatid="7636" lane="3" entrytime="00:00:31.19" />
                <RESULT eventid="1470" points="252" reactiontime="+72" swimtime="00:01:17.39" resultid="4862" heatid="7667" lane="6" entrytime="00:01:17.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="260" reactiontime="+89" swimtime="00:01:15.90" resultid="4863" heatid="7745" lane="6" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="240" reactiontime="+72" swimtime="00:02:50.57" resultid="4864" heatid="7768" lane="2" entrytime="00:02:49.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:22.07" />
                    <SPLIT distance="150" swimtime="00:02:06.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-07" firstname="Marcin" gender="M" lastname="Musialik" nation="POL" athleteid="4865">
              <RESULTS>
                <RESULT eventid="1200" points="321" reactiontime="+66" swimtime="00:00:33.02" resultid="4866" heatid="7452" lane="1" entrytime="00:00:34.21" />
                <RESULT eventid="1336" points="371" reactiontime="+88" swimtime="00:02:31.78" resultid="4867" heatid="7570" lane="1" entrytime="00:02:40.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:10.99" />
                    <SPLIT distance="150" swimtime="00:01:51.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="441" reactiontime="+88" swimtime="00:02:10.46" resultid="4868" heatid="7702" lane="2" entrytime="00:02:14.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="100" swimtime="00:01:01.76" />
                    <SPLIT distance="150" swimtime="00:01:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="425" reactiontime="+95" swimtime="00:05:13.20" resultid="4869" heatid="7982" lane="1" entrytime="00:05:28.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:12.47" />
                    <SPLIT distance="150" swimtime="00:01:52.74" />
                    <SPLIT distance="200" swimtime="00:02:32.19" />
                    <SPLIT distance="250" swimtime="00:03:17.50" />
                    <SPLIT distance="300" swimtime="00:04:02.87" />
                    <SPLIT distance="350" swimtime="00:04:39.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="364" reactiontime="+71" swimtime="00:02:28.51" resultid="4870" heatid="7772" lane="1" entrytime="00:02:32.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="150" swimtime="00:01:51.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="454" reactiontime="+92" swimtime="00:04:36.68" resultid="4871" heatid="8048" lane="4" entrytime="00:04:45.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:07.05" />
                    <SPLIT distance="150" swimtime="00:01:42.37" />
                    <SPLIT distance="200" swimtime="00:02:17.63" />
                    <SPLIT distance="250" swimtime="00:02:52.85" />
                    <SPLIT distance="300" swimtime="00:03:27.84" />
                    <SPLIT distance="350" swimtime="00:04:02.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="433" reactiontime="+76" swimtime="00:02:01.31" resultid="4872" heatid="7934" lane="1" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:05.80" />
                    <SPLIT distance="150" swimtime="00:01:33.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4784" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4838" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="4793" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4856" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1377" points="285" reactiontime="+80" swimtime="00:02:19.41" resultid="4873" heatid="7931" lane="6" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:46.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4829" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4802" number="2" reactiontime="+15" />
                    <RELAYPOSITION athleteid="4820" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="4811" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1528" points="421" swimtime="00:01:47.76" resultid="4874" heatid="7715" lane="5" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.68" />
                    <SPLIT distance="100" swimtime="00:00:52.97" />
                    <SPLIT distance="150" swimtime="00:01:21.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4793" number="1" />
                    <RELAYPOSITION athleteid="4856" number="2" />
                    <RELAYPOSITION athleteid="4838" number="3" />
                    <RELAYPOSITION athleteid="4784" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1528" points="285" reactiontime="+81" swimtime="00:02:02.68" resultid="4875" heatid="7713" lane="6" entrytime="00:02:01.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="100" swimtime="00:00:59.34" />
                    <SPLIT distance="150" swimtime="00:01:32.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4829" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4802" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4811" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="4820" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" name="TS Olimpia Poznań" nation="POL" region="WIE">
          <CONTACT name="Pietraszewski" phone="501648415" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Grażyna" gender="F" lastname="Cabaj-Drela" nation="POL" athleteid="4892">
              <RESULTS>
                <RESULT eventid="1058" points="312" reactiontime="+80" swimtime="00:00:34.27" resultid="4893" heatid="7338" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1092" points="306" swimtime="00:03:04.71" resultid="4894" heatid="7386" lane="5" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                    <SPLIT distance="150" swimtime="00:02:20.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="315" swimtime="00:03:17.67" resultid="4895" heatid="7467" lane="5" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.08" />
                    <SPLIT distance="100" swimtime="00:01:35.10" />
                    <SPLIT distance="150" swimtime="00:02:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="315" reactiontime="+90" swimtime="00:01:24.78" resultid="4896" heatid="7532" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="341" swimtime="00:01:29.67" resultid="4897" heatid="7588" lane="5" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1419" points="255" reactiontime="+91" swimtime="00:00:38.43" resultid="4898" heatid="7615" lane="1" entrytime="00:00:42.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1645" points="339" reactiontime="+89" swimtime="00:00:41.27" resultid="4899" heatid="7784" lane="1" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="4900">
              <RESULTS>
                <RESULT eventid="1058" points="217" reactiontime="+92" swimtime="00:00:38.67" resultid="4901" heatid="7336" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1183" points="151" reactiontime="+81" swimtime="00:00:48.16" resultid="4902" heatid="7433" lane="4" entrytime="00:00:52.00" />
                <RESULT eventid="1251" points="176" swimtime="00:01:30.93" resultid="4903" heatid="7489" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="131" reactiontime="+99" swimtime="00:00:47.95" resultid="4904" heatid="7614" lane="6" entrytime="00:00:52.00" />
                <RESULT eventid="1487" points="181" swimtime="00:03:16.46" resultid="4905" heatid="7677" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                    <SPLIT distance="100" swimtime="00:01:36.21" />
                    <SPLIT distance="150" swimtime="00:02:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="184" reactiontime="+103" swimtime="00:00:50.60" resultid="4906" heatid="7777" lane="3" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Joanna" gender="F" lastname="Puchalska" nation="POL" athleteid="4907">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1092" points="437" swimtime="00:02:44.10" resultid="4908" heatid="7388" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:20.62" />
                    <SPLIT distance="150" swimtime="00:02:05.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="405" reactiontime="+92" swimtime="00:03:01.84" resultid="4909" heatid="7469" lane="6" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:01:27.48" />
                    <SPLIT distance="150" swimtime="00:02:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1385" points="400" reactiontime="+89" swimtime="00:01:25.06" resultid="4910" heatid="7590" lane="4" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1542" points="392" reactiontime="+95" swimtime="00:05:56.61" resultid="4911" heatid="7718" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                    <SPLIT distance="150" swimtime="00:02:56.11" />
                    <SPLIT distance="200" swimtime="00:03:45.62" />
                    <SPLIT distance="250" swimtime="00:04:35.53" />
                    <SPLIT distance="300" swimtime="00:05:16.46" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1577" points="400" swimtime="00:01:14.66" resultid="4912" heatid="7735" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="4913">
              <RESULTS>
                <RESULT eventid="1075" points="146" reactiontime="+101" swimtime="00:00:38.52" resultid="4914" heatid="7346" lane="1" />
                <RESULT eventid="1109" points="120" reactiontime="+109" swimtime="00:03:43.12" resultid="4915" heatid="7394" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.15" />
                    <SPLIT distance="100" swimtime="00:01:48.42" />
                    <SPLIT distance="150" swimtime="00:02:53.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="134" reactiontime="+78" swimtime="00:00:44.14" resultid="4916" heatid="7445" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1302" points="132" swimtime="00:01:39.69" resultid="4917" heatid="7541" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="80" swimtime="00:00:50.49" resultid="4918" heatid="7623" lane="5" />
                <RESULT eventid="1470" points="110" reactiontime="+89" swimtime="00:01:42.11" resultid="4919" heatid="7662" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="101" reactiontime="+82" swimtime="00:03:47.42" resultid="4920" heatid="7764" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.43" />
                    <SPLIT distance="100" swimtime="00:01:48.98" />
                    <SPLIT distance="150" swimtime="00:02:47.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="133" reactiontime="+106" swimtime="00:00:49.45" resultid="4921" heatid="7792" lane="1" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="4922">
              <RESULTS>
                <RESULT eventid="1109" points="202" reactiontime="+99" swimtime="00:03:07.46" resultid="4923" heatid="7396" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                    <SPLIT distance="100" swimtime="00:01:33.15" />
                    <SPLIT distance="150" swimtime="00:02:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="166" reactiontime="+76" swimtime="00:00:41.12" resultid="4924" heatid="7446" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1302" points="211" reactiontime="+94" swimtime="00:01:25.22" resultid="4925" heatid="7544" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="183" reactiontime="+76" swimtime="00:01:26.05" resultid="4926" heatid="7664" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="211" reactiontime="+93" swimtime="00:06:35.27" resultid="4927" heatid="7977" lane="4" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.22" />
                    <SPLIT distance="100" swimtime="00:01:42.10" />
                    <SPLIT distance="150" swimtime="00:02:30.57" />
                    <SPLIT distance="200" swimtime="00:03:19.12" />
                    <SPLIT distance="250" swimtime="00:04:12.40" />
                    <SPLIT distance="300" swimtime="00:05:07.04" />
                    <SPLIT distance="350" swimtime="00:05:52.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="184" reactiontime="+81" swimtime="00:03:06.25" resultid="4928" heatid="7766" lane="5" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                    <SPLIT distance="100" swimtime="00:01:31.17" />
                    <SPLIT distance="150" swimtime="00:02:19.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="4929">
              <RESULTS>
                <RESULT eventid="1109" points="294" reactiontime="+79" swimtime="00:02:45.51" resultid="4930" heatid="7399" lane="4" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:22.09" />
                    <SPLIT distance="150" swimtime="00:02:08.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="318" reactiontime="+81" swimtime="00:02:56.74" resultid="4931" heatid="7481" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:25.12" />
                    <SPLIT distance="150" swimtime="00:02:11.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="328" reactiontime="+82" swimtime="00:01:13.55" resultid="4932" heatid="7548" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="365" reactiontime="+79" swimtime="00:01:17.77" resultid="4933" heatid="7607" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="314" reactiontime="+80" swimtime="00:02:26.10" resultid="4934" heatid="7699" lane="3" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                    <SPLIT distance="150" swimtime="00:01:48.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="274" swimtime="00:01:14.61" resultid="4935" heatid="7744" lane="5" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="359" reactiontime="+82" swimtime="00:00:35.52" resultid="4936" heatid="7805" lane="1" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Bartłomiej" gender="M" lastname="Zadorożny" nation="POL" athleteid="4937">
              <RESULTS>
                <RESULT eventid="1075" points="393" reactiontime="+81" swimtime="00:00:27.71" resultid="4938" heatid="7371" lane="3" entrytime="00:00:27.66" />
                <RESULT eventid="1268" points="381" reactiontime="+84" swimtime="00:01:01.98" resultid="4939" heatid="7519" lane="6" entrytime="00:01:01.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="351" reactiontime="+91" swimtime="00:01:11.94" resultid="4940" heatid="7551" lane="4" entrytime="00:01:11.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="363" reactiontime="+87" swimtime="00:01:17.89" resultid="4941" heatid="7606" lane="1" entrytime="00:01:20.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="346" reactiontime="+83" swimtime="00:00:31.03" resultid="4942" heatid="7637" lane="6" entrytime="00:00:31.02" />
                <RESULT eventid="1662" points="379" reactiontime="+83" swimtime="00:00:34.87" resultid="4943" heatid="7808" lane="2" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1126" points="274" reactiontime="+84" swimtime="00:02:04.32" resultid="4944" heatid="7410" lane="2" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                    <SPLIT distance="100" swimtime="00:01:02.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4937" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="4892" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4907" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4929" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" points="285" reactiontime="+72" swimtime="00:02:19.42" resultid="4945" heatid="7818" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:14.81" />
                    <SPLIT distance="150" swimtime="00:01:50.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4892" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4937" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4907" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4929" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WMT" name="Warsaw Masters Team" nation="POL" region="MAZ">
          <CONTACT email="wojciech.kaluzynski@gmail.com" name="Kałużyński Wojciech" phone="607 45 4444" />
          <ATHLETES>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" athleteid="4947">
              <RESULTS>
                <RESULT eventid="1251" points="613" reactiontime="+77" swimtime="00:01:00.04" resultid="4948" heatid="7498" lane="4" entrytime="00:00:59.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="588" reactiontime="+76" swimtime="00:01:08.90" resultid="4949" heatid="7537" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="535" reactiontime="+74" swimtime="00:00:30.02" resultid="4950" heatid="7621" lane="2" entrytime="00:00:29.60" />
                <RESULT eventid="1487" points="550" reactiontime="+78" swimtime="00:02:15.61" resultid="4951" heatid="7685" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="150" swimtime="00:01:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="580" reactiontime="+74" swimtime="00:01:05.99" resultid="4952" heatid="7735" lane="3" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="4953">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1109" points="327" reactiontime="+90" swimtime="00:02:39.67" resultid="4954" heatid="7399" lane="2" entrytime="00:02:49.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                    <SPLIT distance="150" swimtime="00:02:03.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="265" reactiontime="+68" swimtime="00:00:35.18" resultid="4955" heatid="7449" lane="5" entrytime="00:00:36.89" />
                <RESULT comment="Rekord Polski Masters" eventid="1302" points="345" reactiontime="+86" swimtime="00:01:12.33" resultid="4956" heatid="7549" lane="4" entrytime="00:01:14.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="296" reactiontime="+72" swimtime="00:01:13.42" resultid="4957" heatid="7667" lane="3" entrytime="00:01:14.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="297" reactiontime="+72" swimtime="00:02:38.92" resultid="4958" heatid="7771" lane="6" entrytime="00:02:39.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="100" swimtime="00:01:17.55" />
                    <SPLIT distance="150" swimtime="00:01:58.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-14" firstname="Sebastian" gender="M" lastname="Wojciechowski" nation="POL" athleteid="4959">
              <RESULTS>
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="4961" heatid="7691" lane="6" entrytime="00:02:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="4963">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4964" heatid="7353" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4965" heatid="7403" lane="2" entrytime="00:02:35.00" />
                <RESULT eventid="1200" points="387" reactiontime="+74" swimtime="00:00:31.00" resultid="4966" heatid="7454" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1302" points="439" reactiontime="+82" swimtime="00:01:06.77" resultid="4967" heatid="7556" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="407" reactiontime="+76" swimtime="00:01:06.03" resultid="4968" heatid="7671" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="373" reactiontime="+84" swimtime="00:02:27.40" resultid="4969" heatid="7772" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:49.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-07" firstname="Michał" gender="M" lastname="Wasielak" nation="POL" athleteid="4970">
              <RESULTS>
                <RESULT eventid="1075" points="221" reactiontime="+100" swimtime="00:00:33.55" resultid="4971" heatid="7358" lane="3" entrytime="00:00:32.00" />
                <RESULT comment="Przekroczony limit czasu." eventid="1165" reactiontime="+102" status="DSQ" swimtime="00:24:18.60" resultid="4972" heatid="7911" lane="4" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:01:28.04" />
                    <SPLIT distance="150" swimtime="00:02:14.87" />
                    <SPLIT distance="200" swimtime="00:03:02.62" />
                    <SPLIT distance="250" swimtime="00:03:50.44" />
                    <SPLIT distance="300" swimtime="00:04:38.49" />
                    <SPLIT distance="350" swimtime="00:05:26.64" />
                    <SPLIT distance="400" swimtime="00:06:15.28" />
                    <SPLIT distance="450" swimtime="00:07:04.80" />
                    <SPLIT distance="500" swimtime="00:07:53.11" />
                    <SPLIT distance="550" swimtime="00:08:42.15" />
                    <SPLIT distance="600" swimtime="00:09:29.99" />
                    <SPLIT distance="650" swimtime="00:10:18.57" />
                    <SPLIT distance="700" swimtime="00:11:07.02" />
                    <SPLIT distance="750" swimtime="00:11:55.63" />
                    <SPLIT distance="800" swimtime="00:12:44.91" />
                    <SPLIT distance="850" swimtime="00:13:34.50" />
                    <SPLIT distance="900" swimtime="00:14:23.11" />
                    <SPLIT distance="950" swimtime="00:15:13.08" />
                    <SPLIT distance="1000" swimtime="00:16:02.71" />
                    <SPLIT distance="1050" swimtime="00:16:52.55" />
                    <SPLIT distance="1100" swimtime="00:17:42.19" />
                    <SPLIT distance="1150" swimtime="00:18:32.66" />
                    <SPLIT distance="1200" swimtime="00:19:22.06" />
                    <SPLIT distance="1250" swimtime="00:20:11.75" />
                    <SPLIT distance="1300" swimtime="00:21:01.65" />
                    <SPLIT distance="1350" swimtime="00:21:51.83" />
                    <SPLIT distance="1400" swimtime="00:22:42.20" />
                    <SPLIT distance="1450" swimtime="00:23:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="217" swimtime="00:01:14.74" resultid="4973" heatid="7506" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="207" reactiontime="+97" swimtime="00:02:47.74" resultid="4974" heatid="7694" lane="1" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:20.89" />
                    <SPLIT distance="150" swimtime="00:02:05.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="4975" heatid="8055" lane="4" entrytime="00:06:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="4976">
              <RESULTS>
                <RESULT eventid="1109" points="57" reactiontime="+119" swimtime="00:04:44.82" resultid="4977" heatid="7391" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.74" />
                    <SPLIT distance="100" swimtime="00:02:24.28" />
                    <SPLIT distance="150" swimtime="00:03:39.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="72" reactiontime="+120" swimtime="00:04:48.79" resultid="4978" heatid="7471" lane="4" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.70" />
                    <SPLIT distance="100" swimtime="00:02:22.59" />
                    <SPLIT distance="150" swimtime="00:03:37.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="56" reactiontime="+121" swimtime="00:02:12.08" resultid="4979" heatid="7539" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="72" reactiontime="+123" swimtime="00:02:13.28" resultid="4980" heatid="7594" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="35" reactiontime="+76" swimtime="00:02:28.36" resultid="4981" heatid="7661" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="40" reactiontime="+71" swimtime="00:05:08.26" resultid="4982" heatid="7763" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.10" />
                    <SPLIT distance="100" swimtime="00:02:29.98" />
                    <SPLIT distance="150" swimtime="00:03:51.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="83" reactiontime="+116" swimtime="00:00:57.84" resultid="4983" heatid="7790" lane="3" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-20" firstname="Anna" gender="F" lastname="Stanisławska" nation="POL" athleteid="4984">
              <RESULTS>
                <RESULT eventid="1058" points="284" reactiontime="+94" swimtime="00:00:35.34" resultid="4985" heatid="7338" lane="4" entrytime="00:00:35.34" />
                <RESULT eventid="1251" points="256" reactiontime="+106" swimtime="00:01:20.32" resultid="4986" heatid="7486" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="197" reactiontime="+109" swimtime="00:03:27.48" resultid="4987" heatid="7562" lane="4" entrytime="00:03:28.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.76" />
                    <SPLIT distance="100" swimtime="00:01:39.79" />
                    <SPLIT distance="150" swimtime="00:02:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="220" reactiontime="+99" swimtime="00:00:40.34" resultid="4988" heatid="7615" lane="4" entrytime="00:00:40.65" />
                <RESULT eventid="1487" points="230" reactiontime="+110" swimtime="00:03:01.25" resultid="4989" heatid="7678" lane="4" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:01:26.61" />
                    <SPLIT distance="150" swimtime="00:02:15.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="173" reactiontime="+109" swimtime="00:01:38.61" resultid="4990" heatid="7732" lane="4" entrytime="00:01:36.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="191" reactiontime="+106" swimtime="00:00:49.97" resultid="4991" heatid="7780" lane="2" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="4992">
              <RESULTS>
                <RESULT eventid="1234" points="213" reactiontime="+106" swimtime="00:03:21.86" resultid="4993" heatid="7475" lane="3" entrytime="00:03:22.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                    <SPLIT distance="100" swimtime="00:01:34.77" />
                    <SPLIT distance="150" swimtime="00:02:28.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="83" reactiontime="+108" swimtime="00:04:09.72" resultid="4994" heatid="7565" lane="2" entrytime="00:04:53.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.93" />
                    <SPLIT distance="100" swimtime="00:01:55.88" />
                    <SPLIT distance="150" swimtime="00:03:03.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="222" reactiontime="+108" swimtime="00:01:31.83" resultid="4995" heatid="7599" lane="6" entrytime="00:01:32.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="137" reactiontime="+108" swimtime="00:07:36.81" resultid="4996" heatid="7976" lane="2" entrytime="00:07:44.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                    <SPLIT distance="100" swimtime="00:01:49.09" />
                    <SPLIT distance="150" swimtime="00:02:55.09" />
                    <SPLIT distance="200" swimtime="00:04:00.71" />
                    <SPLIT distance="250" swimtime="00:04:52.45" />
                    <SPLIT distance="300" swimtime="00:05:47.10" />
                    <SPLIT distance="350" swimtime="00:06:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="113" swimtime="00:01:40.20" resultid="4997" heatid="7740" lane="5" entrytime="00:01:42.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="213" reactiontime="+100" swimtime="00:00:42.24" resultid="4998" heatid="7795" lane="1" entrytime="00:00:42.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-07-13" firstname="Sebastian" gender="M" lastname="Ostapczuk" nation="POL" athleteid="4999">
              <RESULTS>
                <RESULT eventid="1234" points="156" reactiontime="+103" swimtime="00:03:43.76" resultid="5000" heatid="7475" lane="6" entrytime="00:03:35.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.28" />
                    <SPLIT distance="100" swimtime="00:01:45.85" />
                    <SPLIT distance="150" swimtime="00:02:44.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="152" reactiontime="+98" swimtime="00:01:24.16" resultid="5001" heatid="7502" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="119" swimtime="00:00:44.31" resultid="5002" heatid="7625" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="1504" points="143" reactiontime="+101" swimtime="00:03:09.94" resultid="5003" heatid="7686" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="100" swimtime="00:01:29.18" />
                    <SPLIT distance="150" swimtime="00:02:19.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="5004">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5005" heatid="7351" lane="2" entrytime="00:00:37.00" />
                <RESULT comment="G-3 - Wynurzenie głowy spod lustra wody po starcie poza 15m" eventid="1200" reactiontime="+80" status="DSQ" swimtime="00:00:49.45" resultid="5006" heatid="7445" lane="1" entrytime="00:00:49.00" />
                <RESULT eventid="1268" points="160" reactiontime="+107" swimtime="00:01:22.69" resultid="5007" heatid="7504" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="91" reactiontime="+77" swimtime="00:01:48.69" resultid="5008" heatid="7660" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="134" reactiontime="+103" swimtime="00:03:14.15" resultid="5009" heatid="7689" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                    <SPLIT distance="100" swimtime="00:01:32.92" />
                    <SPLIT distance="150" swimtime="00:02:24.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="74" reactiontime="+85" swimtime="00:04:12.29" resultid="5010" heatid="7763" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.99" />
                    <SPLIT distance="100" swimtime="00:02:02.16" />
                    <SPLIT distance="150" swimtime="00:03:07.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="121" reactiontime="+103" swimtime="00:07:09.20" resultid="5011" heatid="8046" lane="6" entrytime="00:07:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:37.93" />
                    <SPLIT distance="150" swimtime="00:02:32.58" />
                    <SPLIT distance="200" swimtime="00:03:27.87" />
                    <SPLIT distance="250" swimtime="00:04:24.24" />
                    <SPLIT distance="300" swimtime="00:05:20.16" />
                    <SPLIT distance="350" swimtime="00:06:17.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-02" firstname="Natalia" gender="F" lastname="Kifert" nation="POL" athleteid="5012">
              <RESULTS>
                <RESULT eventid="1183" points="325" reactiontime="+70" swimtime="00:00:37.36" resultid="5013" heatid="7438" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1453" points="326" reactiontime="+66" swimtime="00:01:20.17" resultid="5014" heatid="7655" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5015" heatid="7781" lane="5" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-28" firstname="Katarzyna" gender="F" lastname="Dobczyńska" nation="POL" athleteid="5016">
              <RESULTS>
                <RESULT eventid="1183" points="224" reactiontime="+91" swimtime="00:00:42.26" resultid="5017" heatid="7435" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1251" points="234" reactiontime="+103" swimtime="00:01:22.75" resultid="5018" heatid="7491" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="218" reactiontime="+93" swimtime="00:01:31.75" resultid="5019" heatid="7652" lane="1" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="229" reactiontime="+105" swimtime="00:03:01.54" resultid="5020" heatid="7679" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:01:27.69" />
                    <SPLIT distance="150" swimtime="00:02:15.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-18" firstname="Łukasz" gender="M" lastname="Kubiszewski - Jakubiak" nation="POL" athleteid="5021">
              <RESULTS>
                <RESULT eventid="1268" points="294" reactiontime="+95" swimtime="00:01:07.54" resultid="5022" heatid="7513" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="173" reactiontime="+101" swimtime="00:00:39.10" resultid="5023" heatid="7628" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="5024" heatid="7796" lane="2" entrytime="00:00:41.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-10" firstname="Tomasz" gender="M" lastname="Porada" nation="POL" athleteid="5025">
              <RESULTS>
                <RESULT eventid="1075" points="381" reactiontime="+78" swimtime="00:00:27.98" resultid="5026" heatid="7372" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="1165" points="341" reactiontime="+94" swimtime="00:20:16.36" resultid="5027" heatid="7915" lane="4" entrytime="00:20:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:10.44" />
                    <SPLIT distance="150" swimtime="00:01:48.89" />
                    <SPLIT distance="200" swimtime="00:02:27.60" />
                    <SPLIT distance="250" swimtime="00:03:07.03" />
                    <SPLIT distance="300" swimtime="00:03:46.90" />
                    <SPLIT distance="350" swimtime="00:04:26.70" />
                    <SPLIT distance="400" swimtime="00:05:06.73" />
                    <SPLIT distance="450" swimtime="00:05:46.91" />
                    <SPLIT distance="500" swimtime="00:06:26.70" />
                    <SPLIT distance="550" swimtime="00:07:06.98" />
                    <SPLIT distance="600" swimtime="00:07:46.96" />
                    <SPLIT distance="650" swimtime="00:08:27.51" />
                    <SPLIT distance="700" swimtime="00:09:08.03" />
                    <SPLIT distance="750" swimtime="00:09:48.83" />
                    <SPLIT distance="800" swimtime="00:10:30.28" />
                    <SPLIT distance="850" swimtime="00:11:11.27" />
                    <SPLIT distance="900" swimtime="00:11:52.33" />
                    <SPLIT distance="950" swimtime="00:12:33.54" />
                    <SPLIT distance="1000" swimtime="00:13:14.79" />
                    <SPLIT distance="1050" swimtime="00:13:56.23" />
                    <SPLIT distance="1100" swimtime="00:14:37.76" />
                    <SPLIT distance="1150" swimtime="00:15:19.65" />
                    <SPLIT distance="1200" swimtime="00:16:01.76" />
                    <SPLIT distance="1250" swimtime="00:16:44.45" />
                    <SPLIT distance="1300" swimtime="00:17:27.49" />
                    <SPLIT distance="1350" swimtime="00:18:10.13" />
                    <SPLIT distance="1400" swimtime="00:18:52.73" />
                    <SPLIT distance="1450" swimtime="00:19:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="381" swimtime="00:02:46.41" resultid="5028" heatid="7483" lane="5" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:20.69" />
                    <SPLIT distance="150" swimtime="00:02:03.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="356" reactiontime="+81" swimtime="00:01:11.58" resultid="5029" heatid="7551" lane="3" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="367" reactiontime="+89" swimtime="00:01:17.63" resultid="5030" heatid="7607" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="364" reactiontime="+79" swimtime="00:01:07.88" resultid="5032" heatid="7747" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="374" reactiontime="+87" swimtime="00:04:55.30" resultid="5033" heatid="8053" lane="3" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:09.11" />
                    <SPLIT distance="150" swimtime="00:01:46.73" />
                    <SPLIT distance="200" swimtime="00:02:24.58" />
                    <SPLIT distance="250" swimtime="00:03:02.20" />
                    <SPLIT distance="300" swimtime="00:03:40.51" />
                    <SPLIT distance="350" swimtime="00:04:18.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-04" firstname="Ewa" gender="F" lastname="Matlak" nation="POL" athleteid="5034">
              <RESULTS>
                <RESULT eventid="1251" points="271" reactiontime="+83" swimtime="00:01:18.82" resultid="5035" heatid="7493" lane="2" entrytime="00:01:17.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="241" reactiontime="+94" swimtime="00:01:32.76" resultid="5036" heatid="7529" lane="2" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5037" heatid="7778" lane="3" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-31" firstname="Radek" gender="M" lastname="Wysocki" nation="POL" athleteid="5038">
              <RESULTS>
                <RESULT eventid="1268" points="378" reactiontime="+75" swimtime="00:01:02.10" resultid="5039" heatid="7516" lane="6" entrytime="00:01:04.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="301" reactiontime="+80" swimtime="00:01:15.67" resultid="5040" heatid="7542" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="313" reactiontime="+76" swimtime="00:00:32.09" resultid="5041" heatid="7633" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1504" points="343" reactiontime="+82" swimtime="00:02:21.92" resultid="5042" heatid="7698" lane="6" entrytime="00:02:25.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:08.76" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="5043">
              <RESULTS>
                <RESULT eventid="1165" points="151" reactiontime="+116" swimtime="00:26:33.80" resultid="5044" heatid="7908" lane="2" entrytime="00:28:50.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                    <SPLIT distance="100" swimtime="00:01:40.03" />
                    <SPLIT distance="150" swimtime="00:02:35.26" />
                    <SPLIT distance="200" swimtime="00:03:29.00" />
                    <SPLIT distance="250" swimtime="00:04:23.98" />
                    <SPLIT distance="300" swimtime="00:05:18.54" />
                    <SPLIT distance="350" swimtime="00:06:13.39" />
                    <SPLIT distance="400" swimtime="00:07:08.15" />
                    <SPLIT distance="450" swimtime="00:08:02.04" />
                    <SPLIT distance="500" swimtime="00:08:54.83" />
                    <SPLIT distance="550" swimtime="00:09:48.05" />
                    <SPLIT distance="600" swimtime="00:10:41.41" />
                    <SPLIT distance="650" swimtime="00:11:34.96" />
                    <SPLIT distance="700" swimtime="00:12:28.29" />
                    <SPLIT distance="750" swimtime="00:13:21.75" />
                    <SPLIT distance="800" swimtime="00:14:15.24" />
                    <SPLIT distance="850" swimtime="00:15:08.18" />
                    <SPLIT distance="900" swimtime="00:16:01.25" />
                    <SPLIT distance="950" swimtime="00:16:54.87" />
                    <SPLIT distance="1000" swimtime="00:17:48.30" />
                    <SPLIT distance="1050" swimtime="00:18:42.22" />
                    <SPLIT distance="1100" swimtime="00:19:34.78" />
                    <SPLIT distance="1150" swimtime="00:20:28.26" />
                    <SPLIT distance="1200" swimtime="00:21:21.12" />
                    <SPLIT distance="1250" swimtime="00:22:13.72" />
                    <SPLIT distance="1300" swimtime="00:23:06.88" />
                    <SPLIT distance="1350" swimtime="00:24:00.60" />
                    <SPLIT distance="1400" swimtime="00:24:54.21" />
                    <SPLIT distance="1450" swimtime="00:25:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="76" reactiontime="+81" swimtime="00:00:53.20" resultid="5045" heatid="7444" lane="1" entrytime="00:00:53.01" />
                <RESULT eventid="1268" points="136" reactiontime="+111" swimtime="00:01:27.29" resultid="5046" heatid="7503" lane="2" entrytime="00:01:27.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="93" reactiontime="+116" swimtime="00:00:48.09" resultid="5047" heatid="7626" lane="6" entrytime="00:00:44.92" />
                <RESULT eventid="1504" points="139" reactiontime="+116" swimtime="00:03:11.45" resultid="5048" heatid="7690" lane="1" entrytime="00:03:02.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:32.87" />
                    <SPLIT distance="150" swimtime="00:02:23.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="144" reactiontime="+108" swimtime="00:06:45.32" resultid="5049" heatid="8047" lane="6" entrytime="00:06:42.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                    <SPLIT distance="100" swimtime="00:01:39.78" />
                    <SPLIT distance="150" swimtime="00:02:32.09" />
                    <SPLIT distance="200" swimtime="00:03:23.68" />
                    <SPLIT distance="250" swimtime="00:04:15.69" />
                    <SPLIT distance="300" swimtime="00:05:07.52" />
                    <SPLIT distance="350" swimtime="00:05:58.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-11" firstname="Sara" gender="F" lastname="Debevec" nation="POL" athleteid="5050">
              <RESULTS>
                <RESULT eventid="1251" points="201" reactiontime="+119" swimtime="00:01:26.94" resultid="5051" heatid="7489" lane="6" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1285" reactiontime="+98" status="DSQ" swimtime="00:01:40.55" resultid="5052" heatid="7528" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="159" reactiontime="+112" swimtime="00:00:45.00" resultid="5053" heatid="7616" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1487" points="213" reactiontime="+118" swimtime="00:03:06.09" resultid="5054" heatid="7678" lane="1" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                    <SPLIT distance="100" swimtime="00:01:30.93" />
                    <SPLIT distance="150" swimtime="00:02:19.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="5055" heatid="7732" lane="5" entrytime="00:01:40.00" />
                <RESULT eventid="1693" points="212" reactiontime="+113" swimtime="00:06:33.94" resultid="8061" heatid="8020" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                    <SPLIT distance="100" swimtime="00:01:32.48" />
                    <SPLIT distance="150" swimtime="00:02:21.88" />
                    <SPLIT distance="200" swimtime="00:03:12.66" />
                    <SPLIT distance="250" swimtime="00:04:03.35" />
                    <SPLIT distance="300" swimtime="00:04:54.41" />
                    <SPLIT distance="350" swimtime="00:05:45.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="5057">
              <RESULTS>
                <RESULT eventid="1058" points="95" reactiontime="+96" swimtime="00:00:50.81" resultid="5058" heatid="7333" lane="2" entrytime="00:00:50.75" />
                <RESULT eventid="1148" points="108" reactiontime="+101" swimtime="00:16:55.34" resultid="5059" heatid="7902" lane="2" entrytime="00:17:25.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.07" />
                    <SPLIT distance="100" swimtime="00:03:05.66" />
                    <SPLIT distance="150" swimtime="00:04:10.55" />
                    <SPLIT distance="200" swimtime="00:06:20.93" />
                    <SPLIT distance="250" swimtime="00:07:25.97" />
                    <SPLIT distance="300" swimtime="00:10:35.67" />
                    <SPLIT distance="350" swimtime="00:15:51.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="81" reactiontime="+72" swimtime="00:01:57.78" resultid="5060" heatid="7487" lane="4" entrytime="00:01:52.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="92" reactiontime="+93" swimtime="00:04:05.68" resultid="5061" heatid="7676" lane="6" entrytime="00:04:06.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:57.29" />
                    <SPLIT distance="100" swimtime="00:03:03.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="100" reactiontime="+91" swimtime="00:08:24.91" resultid="5062" heatid="8019" lane="2" entrytime="00:08:07.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.36" />
                    <SPLIT distance="100" swimtime="00:02:01.29" />
                    <SPLIT distance="150" swimtime="00:03:06.73" />
                    <SPLIT distance="200" swimtime="00:04:10.83" />
                    <SPLIT distance="250" swimtime="00:05:15.29" />
                    <SPLIT distance="300" swimtime="00:06:19.79" />
                    <SPLIT distance="350" swimtime="00:07:23.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-16" firstname="Paweł" gender="M" lastname="Witkowski" nation="POL" athleteid="5063">
              <RESULTS>
                <RESULT eventid="1234" points="385" reactiontime="+96" swimtime="00:02:45.76" resultid="5064" heatid="7483" lane="1" entrytime="00:02:48.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:01:18.79" />
                    <SPLIT distance="150" swimtime="00:02:02.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="442" reactiontime="+92" swimtime="00:01:12.95" resultid="5065" heatid="7608" lane="2" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="153" reactiontime="+88" swimtime="00:00:47.13" resultid="5066" heatid="7810" lane="2" entrytime="00:00:33.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-24" firstname="Marlena" gender="F" lastname="Dobrasiewicz" nation="POL" athleteid="5067">
              <RESULTS>
                <RESULT eventid="1217" points="445" reactiontime="+88" swimtime="00:02:56.19" resultid="5068" heatid="7467" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:26.18" />
                    <SPLIT distance="150" swimtime="00:02:11.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="490" reactiontime="+83" swimtime="00:01:04.67" resultid="5069" heatid="7496" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="432" reactiontime="+87" swimtime="00:01:22.92" resultid="5070" heatid="7589" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="455" reactiontime="+89" swimtime="00:02:24.51" resultid="5071" heatid="7683" lane="3" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:10.55" />
                    <SPLIT distance="150" swimtime="00:01:48.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="439" swimtime="00:05:09.04" resultid="5072" heatid="8025" lane="5" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="150" swimtime="00:01:52.80" />
                    <SPLIT distance="200" swimtime="00:02:32.26" />
                    <SPLIT distance="250" swimtime="00:03:11.98" />
                    <SPLIT distance="300" swimtime="00:03:52.08" />
                    <SPLIT distance="350" swimtime="00:04:31.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Olga" gender="F" lastname="Krysiak" nation="POL" athleteid="5073">
              <RESULTS>
                <RESULT eventid="1058" points="508" reactiontime="+76" swimtime="00:00:29.12" resultid="5074" heatid="7344" lane="6" entrytime="00:00:28.77" />
                <RESULT eventid="1148" points="343" reactiontime="+82" swimtime="00:11:31.77" resultid="5075" heatid="7905" lane="4" entrytime="00:10:45.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                    <SPLIT distance="150" swimtime="00:01:57.64" />
                    <SPLIT distance="200" swimtime="00:02:40.67" />
                    <SPLIT distance="250" swimtime="00:03:23.97" />
                    <SPLIT distance="300" swimtime="00:04:07.32" />
                    <SPLIT distance="350" swimtime="00:04:51.23" />
                    <SPLIT distance="400" swimtime="00:05:35.25" />
                    <SPLIT distance="450" swimtime="00:06:20.35" />
                    <SPLIT distance="500" swimtime="00:07:05.07" />
                    <SPLIT distance="550" swimtime="00:07:50.02" />
                    <SPLIT distance="600" swimtime="00:08:35.22" />
                    <SPLIT distance="650" swimtime="00:09:20.20" />
                    <SPLIT distance="700" swimtime="00:10:05.99" />
                    <SPLIT distance="750" swimtime="00:10:50.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="479" reactiontime="+79" swimtime="00:01:05.16" resultid="5076" heatid="7498" lane="1" entrytime="00:01:02.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="447" reactiontime="+82" swimtime="00:02:25.33" resultid="5077" heatid="7684" lane="4" entrytime="00:02:21.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                    <SPLIT distance="150" swimtime="00:01:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" status="DNS" swimtime="00:00:00.00" resultid="5078" heatid="8024" lane="4" entrytime="00:05:13.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="5079">
              <RESULTS>
                <RESULT eventid="1268" points="392" reactiontime="+81" swimtime="00:01:01.38" resultid="5080" heatid="7519" lane="2" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="360" reactiontime="+88" swimtime="00:01:11.35" resultid="5081" heatid="7550" lane="3" entrytime="00:01:13.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="379" reactiontime="+94" swimtime="00:00:30.12" resultid="5082" heatid="7640" lane="4" entrytime="00:00:29.90" />
                <RESULT eventid="1504" points="379" reactiontime="+87" swimtime="00:02:17.20" resultid="5083" heatid="7701" lane="4" entrytime="00:02:16.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                    <SPLIT distance="150" swimtime="00:01:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="301" reactiontime="+85" swimtime="00:01:12.31" resultid="5084" heatid="7745" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="341" reactiontime="+73" swimtime="00:00:36.11" resultid="5085" heatid="7800" lane="4" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-02" firstname="Tomasz" gender="M" lastname="Jąkalski" nation="POL" athleteid="5086">
              <RESULTS>
                <RESULT eventid="1200" points="427" reactiontime="+62" swimtime="00:00:30.02" resultid="5087" heatid="7458" lane="4" entrytime="00:00:29.50" />
                <RESULT eventid="1302" points="449" reactiontime="+89" swimtime="00:01:06.27" resultid="5088" heatid="7558" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="436" reactiontime="+87" swimtime="00:00:28.74" resultid="5089" heatid="7642" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1470" reactiontime="+70" status="DNS" swimtime="00:00:00.00" resultid="5090" heatid="7672" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="5091" heatid="7773" lane="6" entrytime="00:02:30.00" />
                <RESULT eventid="1662" points="409" reactiontime="+90" swimtime="00:00:34.00" resultid="5092" heatid="7809" lane="4" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="5093">
              <RESULTS>
                <RESULT eventid="1217" points="324" reactiontime="+86" swimtime="00:03:15.73" resultid="5094" heatid="7468" lane="2" entrytime="00:03:10.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                    <SPLIT distance="100" swimtime="00:01:36.82" />
                    <SPLIT distance="150" swimtime="00:02:26.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="322" reactiontime="+83" swimtime="00:01:31.46" resultid="5095" heatid="7589" lane="4" entrytime="00:01:28.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="261" reactiontime="+83" swimtime="00:02:53.76" resultid="5096" heatid="7680" lane="2" entrytime="00:02:51.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                    <SPLIT distance="100" swimtime="00:01:26.33" />
                    <SPLIT distance="150" swimtime="00:02:11.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="309" reactiontime="+84" swimtime="00:00:42.56" resultid="5097" heatid="7785" lane="1" entrytime="00:00:40.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-02-17" firstname="Piotr" gender="M" lastname="Barski" nation="POL" athleteid="5098">
              <RESULTS>
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="5099" heatid="7475" lane="5" entrytime="00:03:35.00" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="5100" heatid="7523" lane="6" entrytime="00:00:58.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="5101" heatid="7608" lane="3" entrytime="00:01:15.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="5102" heatid="7811" lane="5" entrytime="00:00:32.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="5103">
              <RESULTS>
                <RESULT eventid="1075" points="476" swimtime="00:00:25.99" resultid="5104" heatid="7379" lane="5" entrytime="00:00:25.50" />
                <RESULT eventid="1109" points="447" reactiontime="+75" swimtime="00:02:23.89" resultid="5105" heatid="7405" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                    <SPLIT distance="100" swimtime="00:01:06.13" />
                    <SPLIT distance="150" swimtime="00:01:50.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="513" swimtime="00:00:56.12" resultid="5106" heatid="7524" lane="5" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="408" reactiontime="+72" swimtime="00:02:27.10" resultid="5107" heatid="7571" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                    <SPLIT distance="150" swimtime="00:01:45.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="508" reactiontime="+71" swimtime="00:00:27.31" resultid="5108" heatid="7646" lane="2" entrytime="00:00:27.00" />
                <RESULT eventid="1594" reactiontime="+72" status="DNF" swimtime="00:00:00.00" resultid="5110" heatid="7751" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="5111" heatid="7805" lane="6" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="5112">
              <RESULTS>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="5113" heatid="7503" lane="6" entrytime="00:01:31.15" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="5114" heatid="7556" lane="1" entrytime="00:01:07.82" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="5115" heatid="7703" lane="2" entrytime="00:02:11.31" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="5116" heatid="7807" lane="4" entrytime="00:00:34.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-18" firstname="Jacek" gender="M" lastname="Czupryn" nation="POL" athleteid="5117">
              <RESULTS>
                <RESULT eventid="1075" points="323" reactiontime="+92" swimtime="00:00:29.56" resultid="5118" heatid="7364" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1268" points="326" reactiontime="+73" swimtime="00:01:05.26" resultid="5119" heatid="7515" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="252" reactiontime="+90" swimtime="00:00:34.51" resultid="5120" heatid="7630" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1504" points="295" reactiontime="+102" swimtime="00:02:29.15" resultid="5121" heatid="7698" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="150" swimtime="00:01:51.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="248" reactiontime="+96" swimtime="00:00:40.15" resultid="5122" heatid="7798" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1710" points="242" reactiontime="+97" swimtime="00:05:41.19" resultid="5123" heatid="8052" lane="2" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                    <SPLIT distance="200" swimtime="00:02:42.74" />
                    <SPLIT distance="250" swimtime="00:03:27.25" />
                    <SPLIT distance="300" swimtime="00:04:11.82" />
                    <SPLIT distance="350" swimtime="00:04:57.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka - Skorykow" nation="POL" athleteid="5124">
              <RESULTS>
                <RESULT eventid="1058" points="404" reactiontime="+83" swimtime="00:00:31.44" resultid="5125" heatid="7342" lane="1" entrytime="00:00:31.84" />
                <RESULT eventid="1217" points="348" reactiontime="+84" swimtime="00:03:11.30" resultid="5126" heatid="7468" lane="6" entrytime="00:03:14.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:01:30.06" />
                    <SPLIT distance="150" swimtime="00:02:19.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="374" reactiontime="+87" swimtime="00:01:20.10" resultid="5127" heatid="7533" lane="3" entrytime="00:01:23.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="384" reactiontime="+82" swimtime="00:01:26.22" resultid="5128" heatid="7589" lane="2" entrytime="00:01:28.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="347" reactiontime="+85" swimtime="00:00:34.67" resultid="5129" heatid="7619" lane="1" entrytime="00:00:34.90" />
                <RESULT eventid="1645" points="410" swimtime="00:00:38.76" resultid="5130" heatid="7786" lane="5" entrytime="00:00:39.46" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="5131">
              <RESULTS>
                <RESULT eventid="1075" points="452" reactiontime="+70" swimtime="00:00:26.45" resultid="5132" heatid="7376" lane="1" entrytime="00:00:26.50" />
                <RESULT eventid="1109" points="416" reactiontime="+77" swimtime="00:02:27.35" resultid="5133" heatid="7405" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="150" swimtime="00:01:53.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="453" reactiontime="+64" swimtime="00:00:29.43" resultid="5134" heatid="7458" lane="1" entrytime="00:00:29.80" />
                <RESULT eventid="1302" points="453" reactiontime="+71" swimtime="00:01:06.07" resultid="5135" heatid="7558" lane="2" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1436" points="473" reactiontime="+76" swimtime="00:00:27.97" resultid="5136" heatid="7645" lane="6" entrytime="00:00:27.90" />
                <RESULT eventid="1504" points="433" reactiontime="+76" swimtime="00:02:11.25" resultid="5137" heatid="7705" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:04.74" />
                    <SPLIT distance="150" swimtime="00:01:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" reactiontime="+76" status="DNS" swimtime="00:00:00.00" resultid="5138" heatid="7751" lane="1" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="5139" heatid="8057" lane="5" entrytime="00:04:38.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-28" firstname="Paweł" gender="M" lastname="Rogosz" nation="POL" athleteid="5140">
              <RESULTS>
                <RESULT eventid="1109" points="340" swimtime="00:02:37.67" resultid="5141" heatid="7401" lane="5" entrytime="00:02:40.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                    <SPLIT distance="150" swimtime="00:02:02.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="299" swimtime="00:21:11.12" resultid="5142" heatid="7913" lane="5" entrytime="00:22:07.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="100" swimtime="00:01:20.16" />
                    <SPLIT distance="150" swimtime="00:02:03.17" />
                    <SPLIT distance="200" swimtime="00:02:45.96" />
                    <SPLIT distance="250" swimtime="00:03:29.00" />
                    <SPLIT distance="300" swimtime="00:04:11.60" />
                    <SPLIT distance="350" swimtime="00:04:53.95" />
                    <SPLIT distance="400" swimtime="00:05:36.62" />
                    <SPLIT distance="450" swimtime="00:06:18.79" />
                    <SPLIT distance="500" swimtime="00:07:01.54" />
                    <SPLIT distance="550" swimtime="00:07:43.78" />
                    <SPLIT distance="600" swimtime="00:08:26.01" />
                    <SPLIT distance="650" swimtime="00:09:07.98" />
                    <SPLIT distance="700" swimtime="00:09:49.47" />
                    <SPLIT distance="750" swimtime="00:10:31.18" />
                    <SPLIT distance="800" swimtime="00:11:13.21" />
                    <SPLIT distance="850" swimtime="00:11:55.54" />
                    <SPLIT distance="900" swimtime="00:12:37.69" />
                    <SPLIT distance="950" swimtime="00:13:19.82" />
                    <SPLIT distance="1000" swimtime="00:14:02.59" />
                    <SPLIT distance="1050" swimtime="00:14:45.89" />
                    <SPLIT distance="1100" swimtime="00:15:29.01" />
                    <SPLIT distance="1150" swimtime="00:16:11.72" />
                    <SPLIT distance="1200" swimtime="00:16:54.84" />
                    <SPLIT distance="1250" swimtime="00:17:38.07" />
                    <SPLIT distance="1300" swimtime="00:18:21.32" />
                    <SPLIT distance="1350" swimtime="00:19:04.54" />
                    <SPLIT distance="1400" swimtime="00:19:47.89" />
                    <SPLIT distance="1450" swimtime="00:20:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="347" swimtime="00:02:51.61" resultid="5143" heatid="7481" lane="5" entrytime="00:02:55.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                    <SPLIT distance="150" swimtime="00:02:08.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="303" reactiontime="+98" swimtime="00:02:42.43" resultid="5144" heatid="7569" lane="2" entrytime="00:02:48.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="100" swimtime="00:01:19.57" />
                    <SPLIT distance="150" swimtime="00:02:01.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="338" reactiontime="+105" swimtime="00:05:37.93" resultid="5145" heatid="7978" lane="1" entrytime="00:05:45.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:02:03.57" />
                    <SPLIT distance="200" swimtime="00:02:48.75" />
                    <SPLIT distance="250" swimtime="00:03:34.45" />
                    <SPLIT distance="300" swimtime="00:04:19.80" />
                    <SPLIT distance="350" swimtime="00:04:59.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="319" reactiontime="+94" swimtime="00:01:10.92" resultid="5146" heatid="7745" lane="3" entrytime="00:01:14.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="5147" heatid="8052" lane="1" entrytime="00:05:25.38" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-10-20" firstname="Norbert" gender="M" lastname="Stablewski" nation="POL" athleteid="5148">
              <RESULTS>
                <RESULT eventid="1268" points="300" reactiontime="+95" swimtime="00:01:07.07" resultid="5149" heatid="7510" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="283" reactiontime="+99" swimtime="00:01:24.70" resultid="5150" heatid="7607" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-09" firstname="Tomasz" gender="M" lastname="Makomaski" nation="POL" athleteid="5151">
              <RESULTS>
                <RESULT eventid="1234" points="347" reactiontime="+80" swimtime="00:02:51.63" resultid="5152" heatid="7483" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:22.40" />
                    <SPLIT distance="150" swimtime="00:02:07.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="367" swimtime="00:01:10.87" resultid="5153" heatid="7552" lane="5" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="392" reactiontime="+80" swimtime="00:01:15.95" resultid="5154" heatid="7609" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="345" reactiontime="+79" swimtime="00:00:31.07" resultid="5155" heatid="7636" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5156" heatid="7747" lane="5" entrytime="00:01:12.00" />
                <RESULT eventid="1662" points="413" reactiontime="+77" swimtime="00:00:33.89" resultid="5157" heatid="7808" lane="3" entrytime="00:00:34.34" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-21" firstname="Marianna" gender="F" lastname="Gajdus" nation="POL" athleteid="5158">
              <RESULTS>
                <RESULT eventid="1217" points="307" reactiontime="+76" swimtime="00:03:19.40" resultid="5159" heatid="7467" lane="2" entrytime="00:03:21.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                    <SPLIT distance="100" swimtime="00:01:36.06" />
                    <SPLIT distance="150" swimtime="00:02:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="352" reactiontime="+79" swimtime="00:01:21.74" resultid="5160" heatid="7534" lane="2" entrytime="00:01:20.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="296" reactiontime="+76" swimtime="00:01:34.02" resultid="5161" heatid="7587" lane="3" entrytime="00:01:33.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="319" reactiontime="+77" swimtime="00:02:42.54" resultid="5162" heatid="7682" lane="3" entrytime="00:02:37.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:01:18.03" />
                    <SPLIT distance="150" swimtime="00:02:00.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="314" reactiontime="+80" swimtime="00:01:20.96" resultid="5163" heatid="7734" lane="1" entrytime="00:01:22.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="301" reactiontime="+74" swimtime="00:05:50.20" resultid="5164" heatid="8023" lane="6" entrytime="00:05:45.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:22.85" />
                    <SPLIT distance="150" swimtime="00:02:08.28" />
                    <SPLIT distance="200" swimtime="00:02:53.89" />
                    <SPLIT distance="250" swimtime="00:03:39.23" />
                    <SPLIT distance="300" swimtime="00:04:24.81" />
                    <SPLIT distance="350" swimtime="00:05:09.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-28" firstname="Krzysztof" gender="M" lastname="Olszewski" nation="POL" athleteid="5165">
              <RESULTS>
                <RESULT eventid="1109" points="407" reactiontime="+83" swimtime="00:02:28.54" resultid="5166" heatid="7401" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                    <SPLIT distance="150" swimtime="00:01:54.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="386" reactiontime="+79" swimtime="00:02:45.70" resultid="5167" heatid="7482" lane="6" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                    <SPLIT distance="150" swimtime="00:02:03.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="469" swimtime="00:01:05.31" resultid="5168" heatid="7556" lane="5" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="419" reactiontime="+82" swimtime="00:01:14.27" resultid="5169" heatid="7609" lane="1" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="322" reactiontime="+83" swimtime="00:01:10.72" resultid="5170" heatid="7736" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="481" reactiontime="+78" swimtime="00:00:32.22" resultid="5171" heatid="7810" lane="1" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="F" lastname="Nawrocka" nation="POL" athleteid="5172">
              <RESULTS>
                <RESULT eventid="1092" points="402" reactiontime="+84" swimtime="00:02:48.79" resultid="5173" heatid="7389" lane="2" entrytime="00:02:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:02:06.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="484" reactiontime="+79" swimtime="00:01:13.54" resultid="5174" heatid="7536" lane="4" entrytime="00:01:13.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="388" reactiontime="+88" swimtime="00:01:25.91" resultid="5175" heatid="7591" lane="1" entrytime="00:01:22.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="347" reactiontime="+76" swimtime="00:01:18.58" resultid="5176" heatid="7657" lane="6" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="394" reactiontime="+86" swimtime="00:00:39.26" resultid="5177" heatid="7786" lane="1" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="Kozak" nation="POL" athleteid="5178">
              <RESULTS>
                <RESULT eventid="1075" points="322" swimtime="00:00:29.59" resultid="5179" heatid="7375" lane="4" entrytime="00:00:26.70" />
                <RESULT eventid="1234" points="414" reactiontime="+96" swimtime="00:02:41.78" resultid="5180" heatid="7484" lane="1" entrytime="00:02:39.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="150" swimtime="00:02:00.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="515" reactiontime="+92" swimtime="00:01:09.36" resultid="5181" heatid="7610" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="523" reactiontime="+90" swimtime="00:00:31.33" resultid="5182" heatid="7813" lane="6" entrytime="00:00:30.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="5183">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5184" heatid="7375" lane="2" entrytime="00:00:26.70" />
                <RESULT eventid="1200" points="404" reactiontime="+77" swimtime="00:00:30.58" resultid="5185" heatid="7456" lane="5" entrytime="00:00:30.90" />
                <RESULT eventid="1268" reactiontime="+75" status="DNF" swimtime="00:00:00.00" resultid="5186" heatid="7521" lane="2" entrytime="00:00:59.26" />
                <RESULT eventid="1436" points="434" reactiontime="+77" swimtime="00:00:28.78" resultid="5187" heatid="7641" lane="2" entrytime="00:00:29.30" />
                <RESULT eventid="1662" points="319" reactiontime="+71" swimtime="00:00:36.93" resultid="5188" heatid="7801" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-14" firstname="Wojciech" gender="M" lastname="Kałużyński" nation="POL" athleteid="5189">
              <RESULTS>
                <RESULT eventid="1268" points="283" reactiontime="+86" swimtime="00:01:08.38" resultid="5190" heatid="7512" lane="1" entrytime="00:01:07.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="264" reactiontime="+94" swimtime="00:01:19.11" resultid="5191" heatid="7547" lane="1" entrytime="00:01:18.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="240" swimtime="00:00:35.05" resultid="5192" heatid="7629" lane="5" entrytime="00:00:36.11" />
                <RESULT eventid="1504" points="277" reactiontime="+90" swimtime="00:02:32.34" resultid="5193" heatid="7696" lane="1" entrytime="00:02:34.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                    <SPLIT distance="150" swimtime="00:01:54.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="186" reactiontime="+91" swimtime="00:00:44.20" resultid="5194" heatid="7793" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1710" points="260" reactiontime="+86" swimtime="00:05:33.29" resultid="5195" heatid="8051" lane="4" entrytime="00:05:34.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:57.98" />
                    <SPLIT distance="150" swimtime="00:02:39.87" />
                    <SPLIT distance="200" swimtime="00:04:06.54" />
                    <SPLIT distance="250" swimtime="00:04:51.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="5196">
              <RESULTS>
                <RESULT eventid="1075" reactiontime="+75" status="DNS" swimtime="00:00:00.00" resultid="5197" heatid="7380" lane="2" entrytime="00:00:25.30" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="5198" heatid="7457" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1436" points="454" swimtime="00:00:28.35" resultid="5199" heatid="7644" lane="5" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1377" points="530" reactiontime="+65" swimtime="00:01:53.38" resultid="5203" heatid="7934" lane="3" entrytime="00:01:49.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:01.17" />
                    <SPLIT distance="150" swimtime="00:01:28.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5086" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="5178" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="5103" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="5183" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1528" points="497" reactiontime="+81" swimtime="00:01:41.93" resultid="5204" heatid="7716" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.04" />
                    <SPLIT distance="100" swimtime="00:00:51.79" />
                    <SPLIT distance="150" swimtime="00:01:16.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5196" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="5178" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="5103" number="3" reactiontime="+15" />
                    <RELAYPOSITION athleteid="5183" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1377" points="459" reactiontime="+73" swimtime="00:01:58.96" resultid="5205" heatid="7934" lane="6" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                    <SPLIT distance="100" swimtime="00:01:03.41" />
                    <SPLIT distance="150" swimtime="00:01:31.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4963" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="5025" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="5131" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="5038" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="1528" points="373" reactiontime="+71" swimtime="00:01:52.12" resultid="5206" heatid="7715" lane="2" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                    <SPLIT distance="100" swimtime="00:00:54.69" />
                    <SPLIT distance="150" swimtime="00:01:22.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5131" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5038" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4963" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="5148" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1528" points="420" reactiontime="+80" swimtime="00:01:47.78" resultid="5207" heatid="7715" lane="4" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                    <SPLIT distance="100" swimtime="00:00:54.42" />
                    <SPLIT distance="150" swimtime="00:01:21.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5079" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5025" number="2" reactiontime="+14" />
                    <RELAYPOSITION athleteid="5151" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="5086" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="1528" points="307" reactiontime="+91" swimtime="00:01:59.73" resultid="5208" heatid="7713" lane="2" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:00:58.82" />
                    <SPLIT distance="150" swimtime="00:01:28.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5140" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="5117" number="2" reactiontime="+88" />
                    <RELAYPOSITION athleteid="5021" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="5189" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1370" points="423" reactiontime="+80" swimtime="00:02:16.76" resultid="5200" heatid="7573" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:43.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5067" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5124" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4947" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="5158" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1370" points="243" reactiontime="+67" swimtime="00:02:44.52" resultid="5201" heatid="7572" lane="3" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:23.30" />
                    <SPLIT distance="150" swimtime="00:02:08.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5012" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="5034" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="5050" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="4984" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="3">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1521" points="450" reactiontime="+82" swimtime="00:02:01.62" resultid="5202" heatid="7708" lane="3" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                    <SPLIT distance="100" swimtime="00:01:04.38" />
                    <SPLIT distance="150" swimtime="00:01:33.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5124" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="5158" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="5067" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4947" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="10">
              <RESULTS>
                <RESULT eventid="1679" points="413" reactiontime="+74" swimtime="00:02:03.21" resultid="5209" heatid="7819" lane="3" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:01.99" />
                    <SPLIT distance="150" swimtime="00:01:31.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5183" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="5178" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="4947" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="5124" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="11">
              <RESULTS>
                <RESULT eventid="1679" points="358" reactiontime="+57" swimtime="00:02:09.17" resultid="5210" heatid="7819" lane="6" entrytime="00:02:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:01:04.61" />
                    <SPLIT distance="150" swimtime="00:01:40.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5086" number="1" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5151" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="5158" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="5067" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Start Wrocław" nation="POL" region="DOL">
          <CONTACT city="WROCŁAW" email="WZSSTART@POST.PL" fax="071 34 372 81" internet="www.start.wroclaw.pl" name="START WROCŁAW" phone="071 34 302 31" state="DOL" street="NOTECKA 12" zip="54-128" />
          <ATHLETES>
            <ATHLETE birthdate="1974-04-30" firstname="Sebastian" gender="M" lastname="Szymański" nation="POL" athleteid="5245">
              <RESULTS>
                <RESULT eventid="1200" points="277" reactiontime="+86" swimtime="00:00:34.68" resultid="5246" heatid="7451" lane="3" entrytime="00:00:34.34" entrycourse="SCM" />
                <RESULT eventid="1268" points="387" reactiontime="+87" swimtime="00:01:01.63" resultid="5247" heatid="7517" lane="3" entrytime="00:01:02.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="372" reactiontime="+88" swimtime="00:00:30.30" resultid="5248" heatid="7638" lane="3" entrytime="00:00:30.50" entrycourse="SCM" />
                <RESULT eventid="1504" points="356" reactiontime="+94" swimtime="00:02:20.18" resultid="5249" heatid="7699" lane="1" entrytime="00:02:24.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:08.77" />
                    <SPLIT distance="150" swimtime="00:01:45.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="364" reactiontime="+93" swimtime="00:01:07.88" resultid="5250" heatid="7748" lane="4" entrytime="00:01:09.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Sinnet Warszawa" nation="POL">
          <CONTACT email="piotrbarski@uw.edu.pl" name="Besler" />
          <ATHLETES>
            <ATHLETE birthdate="1978-09-25" firstname="Agnieszka" gender="F" lastname="Besler" nation="POL" athleteid="5419">
              <RESULTS>
                <RESULT eventid="1217" status="DNS" swimtime="00:00:00.00" resultid="5420" heatid="7466" lane="3" entrytime="00:03:28.95" />
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="5421" heatid="7588" lane="1" entrytime="00:01:33.15" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5422" heatid="7783" lane="4" entrytime="00:00:43.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Aquapark Wrocław" nation="POL">
          <CONTACT name="Dudek" />
          <ATHLETES>
            <ATHLETE birthdate="1987-05-13" firstname="Marcin" gender="M" lastname="Gajewski" nation="POL" athleteid="5648">
              <RESULTS>
                <RESULT eventid="1302" points="352" reactiontime="+87" swimtime="00:01:11.86" resultid="5649" heatid="7552" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="349" reactiontime="+83" swimtime="00:00:30.95" resultid="5650" heatid="7640" lane="6" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-13" firstname="Maciej" gender="M" lastname="Dąbrowski" nation="POL" athleteid="5651">
              <RESULTS>
                <RESULT eventid="1075" points="284" reactiontime="+97" swimtime="00:00:30.88" resultid="5652" heatid="7363" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1109" points="260" swimtime="00:02:52.39" resultid="5653" heatid="7399" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:18.79" />
                    <SPLIT distance="150" swimtime="00:02:11.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="255" reactiontime="+75" swimtime="00:00:35.64" resultid="5654" heatid="7451" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="281" reactiontime="+95" swimtime="00:01:17.43" resultid="5655" heatid="7547" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="240" reactiontime="+80" swimtime="00:01:18.73" resultid="5656" heatid="7666" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="5657" heatid="7768" lane="5" entrytime="00:02:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-04-05" firstname="Krzysztof" gender="M" lastname="Makowski" nation="POL" athleteid="5658">
              <RESULTS>
                <RESULT eventid="1268" points="458" reactiontime="+83" swimtime="00:00:58.30" resultid="5659" heatid="7524" lane="2" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="497" reactiontime="+86" swimtime="00:00:27.52" resultid="5660" heatid="7646" lane="3" entrytime="00:00:26.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="5661">
              <RESULTS>
                <RESULT eventid="1058" points="239" reactiontime="+87" swimtime="00:00:37.45" resultid="5662" heatid="7335" lane="4" entrytime="00:00:38.31" />
                <RESULT eventid="1148" points="162" reactiontime="+99" swimtime="00:14:48.31" resultid="5663" heatid="7903" lane="1" entrytime="00:14:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                    <SPLIT distance="100" swimtime="00:01:35.40" />
                    <SPLIT distance="150" swimtime="00:02:30.21" />
                    <SPLIT distance="200" swimtime="00:03:25.15" />
                    <SPLIT distance="250" swimtime="00:04:20.86" />
                    <SPLIT distance="300" swimtime="00:05:16.19" />
                    <SPLIT distance="350" swimtime="00:06:13.56" />
                    <SPLIT distance="400" swimtime="00:07:11.33" />
                    <SPLIT distance="450" swimtime="00:08:08.98" />
                    <SPLIT distance="500" swimtime="00:09:07.20" />
                    <SPLIT distance="550" swimtime="00:10:04.54" />
                    <SPLIT distance="600" swimtime="00:11:02.40" />
                    <SPLIT distance="650" swimtime="00:11:58.93" />
                    <SPLIT distance="700" swimtime="00:12:57.71" />
                    <SPLIT distance="750" swimtime="00:13:55.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="206" reactiontime="+93" swimtime="00:01:26.25" resultid="5664" heatid="7489" lane="2" entrytime="00:01:34.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="213" reactiontime="+90" swimtime="00:01:36.68" resultid="5665" heatid="7529" lane="6" entrytime="00:01:37.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="5666" heatid="7586" lane="6" entrytime="00:01:44.58" />
                <RESULT eventid="1487" status="DNS" swimtime="00:00:00.00" resultid="5667" heatid="7677" lane="3" entrytime="00:03:24.16" />
                <RESULT eventid="1645" points="256" reactiontime="+89" swimtime="00:00:45.33" resultid="5668" heatid="7782" lane="1" entrytime="00:00:46.38" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-14" firstname="Mateusz" gender="M" lastname="Kwaśniewski" nation="POL" athleteid="5670">
              <RESULTS>
                <RESULT eventid="1268" points="536" reactiontime="+70" swimtime="00:00:55.29" resultid="5671" heatid="7524" lane="3" entrytime="00:00:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="526" reactiontime="+72" swimtime="00:00:27.00" resultid="5672" heatid="7646" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1504" points="484" reactiontime="+71" swimtime="00:02:06.55" resultid="5673" heatid="7705" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                    <SPLIT distance="100" swimtime="00:01:00.31" />
                    <SPLIT distance="150" swimtime="00:01:33.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" gender="F" lastname="Mongiało" nation="POL" athleteid="5674">
              <RESULTS>
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="5675" heatid="7498" lane="2" entrytime="00:01:02.50" />
                <RESULT eventid="1285" status="WDR" swimtime="00:00:00.00" resultid="5676" entrytime="00:01:12.80" />
                <RESULT eventid="1419" status="DNS" swimtime="00:00:00.00" resultid="5677" heatid="7621" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1487" status="DNS" swimtime="00:00:00.00" resultid="5678" heatid="7685" lane="6" entrytime="00:02:18.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-10-10" firstname="Marek" gender="M" lastname="Rother" nation="POL" athleteid="5679">
              <RESULTS>
                <RESULT eventid="1200" points="446" reactiontime="+64" swimtime="00:00:29.59" resultid="5680" heatid="7458" lane="3" entrytime="00:00:29.50" />
                <RESULT eventid="1302" points="446" reactiontime="+79" swimtime="00:01:06.41" resultid="5681" heatid="7552" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="451" reactiontime="+68" swimtime="00:01:03.80" resultid="5682" heatid="7673" lane="6" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="436" reactiontime="+69" swimtime="00:02:19.86" resultid="5683" heatid="7773" lane="4" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:08.56" />
                    <SPLIT distance="150" swimtime="00:01:44.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-10-10" firstname="Marta" gender="F" lastname="Frank" nation="POL" athleteid="5684">
              <RESULTS>
                <RESULT eventid="1453" points="364" reactiontime="+66" swimtime="00:01:17.31" resultid="5685" heatid="7657" lane="5" entrytime="00:01:16.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" status="DNS" swimtime="00:00:00.00" resultid="5686" heatid="7680" lane="5" entrytime="00:02:52.00" />
                <RESULT eventid="1611" points="313" reactiontime="+71" swimtime="00:02:56.72" resultid="5687" heatid="7760" lane="6" entrytime="00:02:52.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:24.78" />
                    <SPLIT distance="150" swimtime="00:02:11.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-21" firstname="Mateusz" gender="M" lastname="Dudek" nation="POL" athleteid="5688">
              <RESULTS>
                <RESULT eventid="1234" points="462" reactiontime="+76" swimtime="00:02:35.99" resultid="5689" heatid="7484" lane="2" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:01:54.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="525" reactiontime="+73" swimtime="00:01:08.91" resultid="5690" heatid="7610" lane="2" entrytime="00:01:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="533" reactiontime="+75" swimtime="00:00:31.13" resultid="5691" heatid="7812" lane="6" entrytime="00:00:31.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-11-17" firstname="Michał" gender="M" lastname="Stasiaczek" nation="POL" athleteid="5692">
              <RESULTS>
                <RESULT eventid="1302" points="479" reactiontime="+81" swimtime="00:01:04.84" resultid="5693" heatid="7558" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="517" reactiontime="+84" swimtime="00:01:09.28" resultid="5694" heatid="7609" lane="3" entrytime="00:01:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="501" reactiontime="+77" swimtime="00:00:31.78" resultid="5695" heatid="7811" lane="3" entrytime="00:00:31.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-23" firstname="Agnieszka" gender="F" lastname="Bystrzycka" nation="POL" athleteid="5696">
              <RESULTS>
                <RESULT eventid="1217" status="DNS" swimtime="00:00:00.00" resultid="5697" heatid="7469" lane="5" entrytime="00:02:55.00" />
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="5698" heatid="7591" lane="4" entrytime="00:01:18.00" />
                <RESULT eventid="1419" status="DNS" swimtime="00:00:00.00" resultid="5699" heatid="7620" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5700" heatid="7787" lane="2" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-10" firstname="Sebastian" gender="M" lastname="Figarski" nation="POL" athleteid="5701">
              <RESULTS>
                <RESULT eventid="1200" points="448" reactiontime="+68" swimtime="00:00:29.53" resultid="5702" heatid="7459" lane="1" entrytime="00:00:29.20" />
                <RESULT eventid="1302" points="486" reactiontime="+92" swimtime="00:01:04.54" resultid="5703" heatid="7559" lane="1" entrytime="00:01:04.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="481" reactiontime="+65" swimtime="00:01:02.46" resultid="5704" heatid="7673" lane="2" entrytime="00:01:03.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="454" reactiontime="+73" swimtime="00:02:18.00" resultid="5705" heatid="7774" lane="1" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:04.92" />
                    <SPLIT distance="150" swimtime="00:01:41.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-11" firstname="Anna" gender="F" lastname="Głowiak" nation="POL" athleteid="5706">
              <RESULTS>
                <RESULT eventid="1058" points="176" reactiontime="+122" swimtime="00:00:41.48" resultid="5707" heatid="7335" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1183" points="223" reactiontime="+90" swimtime="00:00:42.37" resultid="5708" heatid="7434" lane="1" entrytime="00:00:46.00" />
                <RESULT eventid="1285" points="223" reactiontime="+94" swimtime="00:01:35.10" resultid="5709" heatid="7528" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="197" reactiontime="+93" swimtime="00:01:34.84" resultid="5710" heatid="7650" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-07" firstname="Radosław" gender="M" lastname="Stefurak" nation="POL" athleteid="5711">
              <RESULTS>
                <RESULT eventid="1234" points="233" swimtime="00:03:16.03" resultid="5712" heatid="7480" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                    <SPLIT distance="100" swimtime="00:01:31.39" />
                    <SPLIT distance="150" swimtime="00:02:24.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="227" reactiontime="+99" swimtime="00:01:31.03" resultid="5713" heatid="7603" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="5714" heatid="7693" lane="1" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-01" firstname="Ernest" gender="M" lastname="Hudziak" nation="POL" athleteid="5715">
              <RESULTS>
                <RESULT eventid="1200" points="410" reactiontime="+72" swimtime="00:00:30.42" resultid="5716" heatid="7459" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1302" points="377" reactiontime="+87" swimtime="00:01:10.26" resultid="5717" heatid="7555" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="371" reactiontime="+84" swimtime="00:01:08.06" resultid="5718" heatid="7673" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5719" heatid="7747" lane="2" entrytime="00:01:11.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="512" reactiontime="+62" swimtime="00:01:54.74" resultid="5720" heatid="7934" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:00.96" />
                    <SPLIT distance="150" swimtime="00:01:27.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5701" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="5688" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="5670" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="5648" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="5723" heatid="7714" lane="1" entrytime="00:01:54.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5651" number="1" />
                    <RELAYPOSITION athleteid="5701" number="2" />
                    <RELAYPOSITION athleteid="5679" number="3" />
                    <RELAYPOSITION athleteid="5711" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1377" points="359" reactiontime="+69" swimtime="00:02:09.14" resultid="5721" heatid="7933" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="100" swimtime="00:01:09.80" />
                    <SPLIT distance="150" swimtime="00:01:38.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5679" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="5692" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="5711" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="5651" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="5724" heatid="7716" lane="4" entrytime="00:01:43.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5692" number="1" />
                    <RELAYPOSITION athleteid="5688" number="2" />
                    <RELAYPOSITION athleteid="5670" number="3" />
                    <RELAYPOSITION athleteid="5658" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1370" status="DNS" swimtime="00:00:00.00" resultid="5722" heatid="7573" lane="3" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5684" number="1" />
                    <RELAYPOSITION athleteid="5696" number="2" />
                    <RELAYPOSITION athleteid="5674" number="3" />
                    <RELAYPOSITION athleteid="5706" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1679" points="346" reactiontime="+64" swimtime="00:02:10.66" resultid="5725" heatid="7818" lane="5" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:05.26" />
                    <SPLIT distance="150" swimtime="00:01:34.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5684" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5688" number="2" />
                    <RELAYPOSITION athleteid="5679" number="3" />
                    <RELAYPOSITION athleteid="5661" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="5726" heatid="7819" lane="2" entrytime="00:02:08.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5701" number="1" />
                    <RELAYPOSITION athleteid="5688" number="2" />
                    <RELAYPOSITION athleteid="5674" number="3" />
                    <RELAYPOSITION athleteid="5696" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="IGAN" name="IGAN Mława" nation="POL" region="MAZ">
          <CONTACT city="Mława" name="Szlagor" phone="609621127" state="MAZ" zip="06-500" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Ewa" gender="F" lastname="Szlagor" nation="POL" athleteid="5745">
              <RESULTS>
                <RESULT eventid="1058" points="502" reactiontime="+85" swimtime="00:00:29.25" resultid="5746" heatid="7343" lane="2" entrytime="00:00:29.30" entrycourse="SCM" />
                <RESULT eventid="1285" points="477" swimtime="00:01:13.88" resultid="5747" heatid="7536" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="478" reactiontime="+85" swimtime="00:00:31.17" resultid="5748" heatid="7621" lane="6" entrytime="00:00:31.50" />
                <RESULT eventid="1645" points="514" reactiontime="+83" swimtime="00:00:35.93" resultid="5749" heatid="7787" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" name="UKS Wodnik 29 Katowice" nation="POL" region="SLA">
          <CONTACT email="skoczyt@gmail.com" name="Skoczylas" />
          <ATHLETES>
            <ATHLETE birthdate="1952-01-19" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="5751">
              <RESULTS>
                <RESULT eventid="1075" points="251" reactiontime="+95" swimtime="00:00:32.16" resultid="5752" heatid="7359" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="1268" points="230" reactiontime="+97" swimtime="00:01:13.31" resultid="5753" heatid="7508" lane="1" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="112" swimtime="00:03:46.28" resultid="5754" heatid="7567" lane="5" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                    <SPLIT distance="100" swimtime="00:01:42.75" />
                    <SPLIT distance="150" swimtime="00:02:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="243" reactiontime="+93" swimtime="00:00:34.91" resultid="5755" heatid="7632" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1504" points="162" reactiontime="+101" swimtime="00:03:02.12" resultid="5756" heatid="7691" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                    <SPLIT distance="150" swimtime="00:02:14.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="173" reactiontime="+96" swimtime="00:01:26.97" resultid="5757" heatid="7741" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="5759">
              <RESULTS>
                <RESULT eventid="1075" points="357" reactiontime="+92" swimtime="00:00:28.59" resultid="5760" heatid="7366" lane="4" entrytime="00:00:29.20" />
                <RESULT eventid="1165" points="303" reactiontime="+105" swimtime="00:21:04.70" resultid="5761" heatid="7915" lane="6" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:11.87" />
                    <SPLIT distance="150" swimtime="00:01:50.72" />
                    <SPLIT distance="200" swimtime="00:02:31.01" />
                    <SPLIT distance="250" swimtime="00:03:13.03" />
                    <SPLIT distance="300" swimtime="00:03:54.76" />
                    <SPLIT distance="350" swimtime="00:04:36.83" />
                    <SPLIT distance="400" swimtime="00:05:18.44" />
                    <SPLIT distance="450" swimtime="00:06:00.60" />
                    <SPLIT distance="500" swimtime="00:06:42.70" />
                    <SPLIT distance="550" swimtime="00:07:25.56" />
                    <SPLIT distance="600" swimtime="00:08:07.16" />
                    <SPLIT distance="650" swimtime="00:08:49.34" />
                    <SPLIT distance="700" swimtime="00:09:31.89" />
                    <SPLIT distance="750" swimtime="00:10:13.98" />
                    <SPLIT distance="800" swimtime="00:10:56.01" />
                    <SPLIT distance="850" swimtime="00:11:38.01" />
                    <SPLIT distance="900" swimtime="00:12:20.59" />
                    <SPLIT distance="950" swimtime="00:13:03.22" />
                    <SPLIT distance="1000" swimtime="00:13:45.53" />
                    <SPLIT distance="1050" swimtime="00:14:28.26" />
                    <SPLIT distance="1100" swimtime="00:15:10.41" />
                    <SPLIT distance="1150" swimtime="00:15:53.10" />
                    <SPLIT distance="1200" swimtime="00:16:35.83" />
                    <SPLIT distance="1250" swimtime="00:17:19.45" />
                    <SPLIT distance="1300" swimtime="00:18:04.35" />
                    <SPLIT distance="1350" swimtime="00:18:49.62" />
                    <SPLIT distance="1400" swimtime="00:19:35.31" />
                    <SPLIT distance="1450" swimtime="00:20:20.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="264" reactiontime="+85" swimtime="00:00:35.24" resultid="5762" heatid="7450" lane="5" entrytime="00:00:35.50" />
                <RESULT eventid="1268" points="358" reactiontime="+100" swimtime="00:01:03.24" resultid="5763" heatid="7516" lane="3" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="327" reactiontime="+104" swimtime="00:02:24.15" resultid="5764" heatid="7698" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="150" swimtime="00:01:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="332" swimtime="00:05:07.09" resultid="5765" heatid="8052" lane="5" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:10.56" />
                    <SPLIT distance="150" swimtime="00:01:49.71" />
                    <SPLIT distance="200" swimtime="00:02:29.61" />
                    <SPLIT distance="250" swimtime="00:03:09.37" />
                    <SPLIT distance="300" swimtime="00:03:49.52" />
                    <SPLIT distance="350" swimtime="00:04:28.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-15" firstname="Andrzej" gender="M" lastname="Porszke" nation="POL" athleteid="5766">
              <RESULTS>
                <RESULT eventid="1075" points="174" reactiontime="+94" swimtime="00:00:36.34" resultid="5767" heatid="7352" lane="1" entrytime="00:00:35.50" />
                <RESULT eventid="1234" points="229" reactiontime="+88" swimtime="00:03:17.16" resultid="5768" heatid="7476" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.87" />
                    <SPLIT distance="100" swimtime="00:01:32.86" />
                    <SPLIT distance="150" swimtime="00:02:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="244" reactiontime="+92" swimtime="00:01:28.91" resultid="5769" heatid="7600" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="251" reactiontime="+82" swimtime="00:00:40.02" resultid="5770" heatid="7797" lane="1" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="5771">
              <RESULTS>
                <RESULT eventid="1075" points="339" reactiontime="+98" swimtime="00:00:29.11" resultid="5772" heatid="7367" lane="4" entrytime="00:00:28.65" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="5773" heatid="7511" lane="6" entrytime="00:01:09.21" />
                <RESULT eventid="1436" points="323" reactiontime="+95" swimtime="00:00:31.77" resultid="5774" heatid="7636" lane="1" entrytime="00:00:31.61" />
                <RESULT eventid="1594" points="273" reactiontime="+95" swimtime="00:01:14.65" resultid="5775" heatid="7746" lane="4" entrytime="00:01:12.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="5776">
              <RESULTS>
                <RESULT eventid="1109" points="243" reactiontime="+94" swimtime="00:02:56.38" resultid="5777" heatid="7398" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:23.21" />
                    <SPLIT distance="150" swimtime="00:02:11.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="293" reactiontime="+84" swimtime="00:03:01.63" resultid="5778" heatid="7478" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:25.43" />
                    <SPLIT distance="150" swimtime="00:02:13.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="274" reactiontime="+90" swimtime="00:01:18.11" resultid="5779" heatid="7548" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="325" reactiontime="+91" swimtime="00:01:20.87" resultid="5780" heatid="7605" lane="3" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="5781" heatid="7982" lane="5" entrytime="00:06:40.00" />
                <RESULT eventid="1662" points="363" reactiontime="+85" swimtime="00:00:35.37" resultid="5782" heatid="7805" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-09" firstname="Krystyna" gender="F" lastname="Nicpoń" nation="POL" athleteid="5783">
              <RESULTS>
                <RESULT eventid="1183" points="105" reactiontime="+83" swimtime="00:00:54.43" resultid="5784" heatid="7433" lane="1" entrytime="00:00:54.00" />
                <RESULT eventid="1453" points="103" reactiontime="+80" swimtime="00:01:57.51" resultid="5785" heatid="7649" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.49" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G-3 - Wynurzenie głowy spod lustra wody po starcie poza 15m" eventid="1611" reactiontime="+83" status="DSQ" swimtime="00:04:09.15" resultid="5786" heatid="7755" lane="6" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.47" />
                    <SPLIT distance="100" swimtime="00:02:00.84" />
                    <SPLIT distance="150" swimtime="00:03:05.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-05" firstname="Marcin" gender="M" lastname="Szczypiński" nation="POL" athleteid="5787">
              <RESULTS>
                <RESULT eventid="1075" points="555" reactiontime="+79" swimtime="00:00:24.70" resultid="5788" heatid="7380" lane="4" entrytime="00:00:24.50" />
                <RESULT eventid="1200" points="506" reactiontime="+70" swimtime="00:00:28.36" resultid="5789" heatid="7458" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="1268" points="597" reactiontime="+80" swimtime="00:00:53.36" resultid="5790" heatid="7499" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="577" reactiontime="+78" swimtime="00:00:58.23" resultid="5791" heatid="7752" lane="6" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="545" reactiontime="+84" swimtime="00:04:20.44" resultid="5792" heatid="8058" lane="2" entrytime="00:04:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:02.06" />
                    <SPLIT distance="150" swimtime="00:01:35.63" />
                    <SPLIT distance="200" swimtime="00:02:09.31" />
                    <SPLIT distance="250" swimtime="00:02:42.57" />
                    <SPLIT distance="300" swimtime="00:03:15.71" />
                    <SPLIT distance="350" swimtime="00:03:48.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-11-14" firstname="Aleksander" gender="M" lastname="Aleksandrowicz" nation="POL" athleteid="5793">
              <RESULTS>
                <RESULT eventid="1075" points="94" reactiontime="+104" swimtime="00:00:44.49" resultid="5794" heatid="7349" lane="4" entrytime="00:00:41.18" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="5795" heatid="7443" lane="3" entrytime="00:00:55.66" />
                <RESULT eventid="1234" points="63" reactiontime="+111" swimtime="00:05:02.18" resultid="5796" heatid="7471" lane="3" entrytime="00:04:50.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.74" />
                    <SPLIT distance="100" swimtime="00:02:24.23" />
                    <SPLIT distance="150" swimtime="00:03:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="65" reactiontime="+117" swimtime="00:02:17.99" resultid="5797" heatid="7594" lane="4" entrytime="00:02:13.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="60" reactiontime="+80" swimtime="00:02:04.86" resultid="5798" heatid="7661" lane="4" entrytime="00:02:01.55" />
                <RESULT eventid="1662" points="73" swimtime="00:01:00.31" resultid="5799" heatid="7790" lane="5" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-08-30" firstname="Aleksandra" gender="F" lastname="Kącki" nation="POL" athleteid="5800">
              <RESULTS>
                <RESULT eventid="1058" points="185" reactiontime="+104" swimtime="00:00:40.79" resultid="5801" heatid="7334" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1251" points="157" reactiontime="+108" swimtime="00:01:34.52" resultid="5802" heatid="7488" lane="1" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-05-18" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="5803">
              <RESULTS>
                <RESULT eventid="1453" points="42" reactiontime="+82" swimtime="00:02:38.46" resultid="5804" heatid="7649" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="37" reactiontime="+122" swimtime="00:05:31.78" resultid="5805" heatid="7675" lane="2" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.96" />
                    <SPLIT distance="100" swimtime="00:02:43.03" />
                    <SPLIT distance="150" swimtime="00:04:13.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="41" reactiontime="+96" swimtime="00:05:48.05" resultid="5806" heatid="7754" lane="2" entrytime="00:05:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.66" />
                    <SPLIT distance="100" swimtime="00:02:51.07" />
                    <SPLIT distance="150" swimtime="00:04:23.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-08-07" firstname="Marzena" gender="F" lastname="Fligier" nation="POL" athleteid="5808">
              <RESULTS>
                <RESULT eventid="1217" points="174" reactiontime="+100" swimtime="00:04:01.00" resultid="5809" heatid="7464" lane="3" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.76" />
                    <SPLIT distance="100" swimtime="00:01:53.09" />
                    <SPLIT distance="150" swimtime="00:02:57.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="205" swimtime="00:01:46.19" resultid="5810" heatid="7585" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-10" firstname="Sandra" gender="F" lastname="Pietrzak" nation="POL" athleteid="5811">
              <RESULTS>
                <RESULT eventid="1058" points="537" swimtime="00:00:28.59" resultid="5812" heatid="7341" lane="5" entrytime="00:00:32.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1148" points="537" reactiontime="+81" swimtime="00:09:55.78" resultid="5813" heatid="7906" lane="2" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:07.34" />
                    <SPLIT distance="150" swimtime="00:01:42.78" />
                    <SPLIT distance="200" swimtime="00:02:19.40" />
                    <SPLIT distance="250" swimtime="00:02:55.82" />
                    <SPLIT distance="300" swimtime="00:03:33.13" />
                    <SPLIT distance="350" swimtime="00:04:10.46" />
                    <SPLIT distance="400" swimtime="00:04:48.58" />
                    <SPLIT distance="450" swimtime="00:05:26.69" />
                    <SPLIT distance="500" swimtime="00:06:04.62" />
                    <SPLIT distance="550" swimtime="00:06:43.26" />
                    <SPLIT distance="600" swimtime="00:07:21.53" />
                    <SPLIT distance="650" swimtime="00:08:00.01" />
                    <SPLIT distance="700" swimtime="00:08:39.09" />
                    <SPLIT distance="750" swimtime="00:09:17.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="450" reactiontime="+69" swimtime="00:00:33.53" resultid="5814" heatid="7440" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1251" points="560" reactiontime="+79" swimtime="00:01:01.85" resultid="5815" heatid="7495" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="457" reactiontime="+76" swimtime="00:00:31.63" resultid="5816" heatid="7619" lane="3" entrytime="00:00:34.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1542" points="506" swimtime="00:05:27.52" resultid="5817" heatid="7718" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="150" swimtime="00:01:54.57" />
                    <SPLIT distance="200" swimtime="00:02:37.32" />
                    <SPLIT distance="250" swimtime="00:03:23.34" />
                    <SPLIT distance="300" swimtime="00:04:11.26" />
                    <SPLIT distance="350" swimtime="00:04:50.20" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1693" points="545" swimtime="00:04:47.59" resultid="5818" heatid="8023" lane="5" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:07.56" />
                    <SPLIT distance="150" swimtime="00:01:43.17" />
                    <SPLIT distance="200" swimtime="00:02:19.41" />
                    <SPLIT distance="250" swimtime="00:02:55.91" />
                    <SPLIT distance="300" swimtime="00:03:33.12" />
                    <SPLIT distance="350" swimtime="00:04:10.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-26" firstname="Piotr" gender="M" lastname="Klepacki" nation="POL" athleteid="5819">
              <RESULTS>
                <RESULT eventid="1075" points="235" swimtime="00:00:32.87" resultid="5820" heatid="7351" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1200" points="111" reactiontime="+70" swimtime="00:00:47.02" resultid="5821" heatid="7445" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1268" points="155" reactiontime="+77" swimtime="00:01:23.52" resultid="5822" heatid="7504" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="5823" heatid="7662" lane="6" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-08" firstname="Paweł" gender="M" lastname="Dygdoń" nation="POL" athleteid="5824">
              <RESULTS>
                <RESULT eventid="1109" points="278" reactiontime="+80" swimtime="00:02:48.52" resultid="5825" heatid="7401" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:02:06.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="252" reactiontime="+93" swimtime="00:22:24.85" resultid="5826" heatid="7914" lane="2" entrytime="00:21:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:57.24" />
                    <SPLIT distance="200" swimtime="00:02:40.04" />
                    <SPLIT distance="250" swimtime="00:03:23.91" />
                    <SPLIT distance="300" swimtime="00:04:08.57" />
                    <SPLIT distance="350" swimtime="00:04:53.91" />
                    <SPLIT distance="400" swimtime="00:05:39.77" />
                    <SPLIT distance="450" swimtime="00:06:26.27" />
                    <SPLIT distance="500" swimtime="00:07:13.53" />
                    <SPLIT distance="550" swimtime="00:08:00.69" />
                    <SPLIT distance="600" swimtime="00:08:48.25" />
                    <SPLIT distance="650" swimtime="00:09:35.49" />
                    <SPLIT distance="700" swimtime="00:10:22.62" />
                    <SPLIT distance="750" swimtime="00:11:10.25" />
                    <SPLIT distance="800" swimtime="00:11:58.27" />
                    <SPLIT distance="850" swimtime="00:12:45.82" />
                    <SPLIT distance="900" swimtime="00:13:33.80" />
                    <SPLIT distance="950" swimtime="00:14:21.58" />
                    <SPLIT distance="1000" swimtime="00:15:09.79" />
                    <SPLIT distance="1050" swimtime="00:15:58.01" />
                    <SPLIT distance="1100" swimtime="00:16:47.06" />
                    <SPLIT distance="1150" swimtime="00:17:35.28" />
                    <SPLIT distance="1200" swimtime="00:18:23.26" />
                    <SPLIT distance="1250" swimtime="00:19:11.96" />
                    <SPLIT distance="1300" swimtime="00:20:00.01" />
                    <SPLIT distance="1350" swimtime="00:20:48.03" />
                    <SPLIT distance="1400" swimtime="00:21:35.59" />
                    <SPLIT distance="1450" swimtime="00:22:22.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="5827" heatid="7454" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="5828" heatid="7550" lane="5" entrytime="00:01:14.00" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="5829" heatid="7667" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1594" points="372" reactiontime="+83" swimtime="00:01:07.37" resultid="5831" heatid="7747" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="263" reactiontime="+73" swimtime="00:02:45.48" resultid="5832" heatid="7769" lane="3" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:18.71" />
                    <SPLIT distance="150" swimtime="00:02:03.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-12-22" firstname="Sylwia" gender="F" lastname="Kornaś" nation="POL" athleteid="5833">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="5834" heatid="7338" lane="1" entrytime="00:00:35.85" />
                <RESULT eventid="1183" status="DNS" swimtime="00:00:00.00" resultid="5835" heatid="7435" lane="6" entrytime="00:00:44.79" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="5836" heatid="7490" lane="4" entrytime="00:01:26.05" />
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="5837" heatid="7651" lane="1" entrytime="00:01:38.12" />
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="5838" heatid="7756" lane="5" entrytime="00:03:28.79" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5839" heatid="7781" lane="6" entrytime="00:00:48.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-16" firstname="Michał" gender="M" lastname="Spławiński " nation="POL" athleteid="6450">
              <RESULTS>
                <RESULT eventid="1075" points="525" reactiontime="+77" swimtime="00:00:25.15" resultid="6451" heatid="7379" lane="4" entrytime="00:00:25.10" />
                <RESULT eventid="1302" points="504" reactiontime="+76" swimtime="00:01:03.78" resultid="6452" heatid="7560" lane="6" entrytime="00:01:02.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="6453" heatid="7610" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="1436" points="547" reactiontime="+75" swimtime="00:00:26.65" resultid="6454" heatid="7645" lane="2" entrytime="00:00:27.30" />
                <RESULT eventid="1662" points="571" reactiontime="+77" swimtime="00:00:30.42" resultid="6455" heatid="7813" lane="1" entrytime="00:00:30.84" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-24" firstname="Paulina" gender="F" lastname="Szuła" nation="POL" athleteid="6456">
              <RESULTS>
                <RESULT eventid="1058" points="538" swimtime="00:00:28.57" resultid="6457" heatid="7344" lane="5" entrytime="00:00:28.10" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="6458" heatid="7498" lane="5" entrytime="00:01:02.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Michał" gender="M" lastname="Sapoń" nation="POL" athleteid="6459">
              <RESULTS>
                <RESULT eventid="1268" points="360" swimtime="00:01:03.17" resultid="6460" heatid="7515" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="388" reactiontime="+86" swimtime="00:00:29.88" resultid="6461" heatid="7643" lane="6" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="Marek" gender="M" lastname="Mróz " nation="POL" athleteid="6463">
              <RESULTS>
                <RESULT eventid="1075" points="485" reactiontime="+80" swimtime="00:00:25.82" resultid="6464" heatid="7378" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1268" points="504" reactiontime="+90" swimtime="00:00:56.47" resultid="6465" heatid="7523" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="472" reactiontime="+83" swimtime="00:00:27.99" resultid="6466" heatid="7644" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1504" points="432" swimtime="00:02:11.38" resultid="6467" heatid="7696" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:04.68" />
                    <SPLIT distance="150" swimtime="00:01:38.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Adam" gender="M" lastname="Krzystolik" nation="POL" athleteid="6468">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="6469" heatid="7356" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="6470" heatid="7543" lane="5" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Joanna" gender="F" lastname="Ziółkowska" nation="POL" athleteid="6471">
              <RESULTS>
                <RESULT eventid="1645" points="231" reactiontime="+81" swimtime="00:00:46.89" resultid="6472" heatid="7782" lane="2" entrytime="00:00:46.00" />
                <RESULT eventid="1487" points="131" reactiontime="+82" swimtime="00:03:38.81" resultid="7943" heatid="7675" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.70" />
                    <SPLIT distance="100" swimtime="00:01:40.92" />
                    <SPLIT distance="150" swimtime="00:02:41.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="295" reactiontime="+85" swimtime="00:02:17.89" resultid="5840" heatid="7931" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:12.00" />
                    <SPLIT distance="150" swimtime="00:01:47.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5759" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="5776" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="5751" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="5771" number="4" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="5841" heatid="7712" lane="6" entrytime="00:02:06.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5759" number="1" />
                    <RELAYPOSITION athleteid="5776" number="2" />
                    <RELAYPOSITION athleteid="5751" number="3" />
                    <RELAYPOSITION athleteid="5771" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="6462" heatid="7715" lane="3" entrytime="00:01:48.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6459" number="1" />
                    <RELAYPOSITION athleteid="6450" number="2" />
                    <RELAYPOSITION athleteid="5787" number="3" />
                    <RELAYPOSITION athleteid="6463" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="5842" heatid="7410" lane="4" entrytime="00:02:03.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5811" number="1" />
                    <RELAYPOSITION athleteid="5819" number="2" />
                    <RELAYPOSITION athleteid="5833" number="3" />
                    <RELAYPOSITION athleteid="5787" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="5843" heatid="7817" lane="3" entrytime="00:02:18.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5811" number="1" />
                    <RELAYPOSITION athleteid="5833" number="2" />
                    <RELAYPOSITION athleteid="5787" number="3" />
                    <RELAYPOSITION athleteid="5819" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TOTOR" name="Toruńczyk Masters Toruń" nation="POL" region="KUJ">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="5850">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="5851" heatid="7385" lane="3" entrytime="00:03:15.00" />
                <RESULT eventid="1217" points="233" reactiontime="+82" swimtime="00:03:38.46" resultid="5853" heatid="7465" lane="1" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.04" />
                    <SPLIT distance="100" swimtime="00:01:46.21" />
                    <SPLIT distance="150" swimtime="00:02:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1319" points="156" reactiontime="+84" swimtime="00:03:44.35" resultid="5854" heatid="7562" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                    <SPLIT distance="100" swimtime="00:01:41.79" />
                    <SPLIT distance="150" swimtime="00:02:42.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="5855" heatid="7586" lane="3" entrytime="00:01:38.00" />
                <RESULT eventid="1542" points="291" reactiontime="+80" swimtime="00:06:33.79" resultid="5856" heatid="7717" lane="1" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:01:37.78" />
                    <SPLIT distance="150" swimtime="00:02:26.85" />
                    <SPLIT distance="200" swimtime="00:03:15.08" />
                    <SPLIT distance="250" swimtime="00:04:09.22" />
                    <SPLIT distance="300" swimtime="00:05:03.79" />
                    <SPLIT distance="350" swimtime="00:05:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="287" reactiontime="+74" swimtime="00:03:01.82" resultid="5857" heatid="7757" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:01:30.52" />
                    <SPLIT distance="150" swimtime="00:02:16.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" status="DNS" swimtime="00:00:00.00" resultid="5858" heatid="8021" lane="3" entrytime="00:06:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-10-22" firstname="Maciej" gender="M" lastname="Muszyński" nation="POL" athleteid="5859">
              <RESULTS>
                <RESULT eventid="1075" points="376" reactiontime="+96" swimtime="00:00:28.11" resultid="5860" heatid="7369" lane="4" entrytime="00:00:28.09" />
                <RESULT eventid="1200" points="289" reactiontime="+79" swimtime="00:00:34.19" resultid="5861" heatid="7452" lane="6" entrytime="00:00:34.25" />
                <RESULT eventid="1268" points="330" reactiontime="+99" swimtime="00:01:05.02" resultid="5862" heatid="7513" lane="2" entrytime="00:01:06.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="314" reactiontime="+98" swimtime="00:00:32.07" resultid="5863" heatid="7634" lane="6" entrytime="00:00:32.60" />
                <RESULT eventid="1594" points="162" reactiontime="+90" swimtime="00:01:28.81" resultid="5864" heatid="7736" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-06" firstname="Arkadiusz" gender="M" lastname="Doliński" nation="POL" athleteid="5865">
              <RESULTS>
                <RESULT eventid="1075" points="382" reactiontime="+90" swimtime="00:00:27.96" resultid="5866" heatid="7370" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1165" points="245" swimtime="00:22:38.16" resultid="5867" heatid="7912" lane="5" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                    <SPLIT distance="150" swimtime="00:02:00.99" />
                    <SPLIT distance="200" swimtime="00:02:44.45" />
                    <SPLIT distance="250" swimtime="00:03:28.26" />
                    <SPLIT distance="300" swimtime="00:04:12.34" />
                    <SPLIT distance="350" swimtime="00:04:56.62" />
                    <SPLIT distance="400" swimtime="00:05:41.52" />
                    <SPLIT distance="450" swimtime="00:06:26.54" />
                    <SPLIT distance="500" swimtime="00:07:12.05" />
                    <SPLIT distance="550" swimtime="00:07:57.94" />
                    <SPLIT distance="600" swimtime="00:08:43.82" />
                    <SPLIT distance="650" swimtime="00:09:29.67" />
                    <SPLIT distance="700" swimtime="00:10:15.48" />
                    <SPLIT distance="750" swimtime="00:11:01.83" />
                    <SPLIT distance="800" swimtime="00:11:49.01" />
                    <SPLIT distance="850" swimtime="00:12:35.98" />
                    <SPLIT distance="900" swimtime="00:13:22.89" />
                    <SPLIT distance="950" swimtime="00:14:09.55" />
                    <SPLIT distance="1000" swimtime="00:14:56.13" />
                    <SPLIT distance="1050" swimtime="00:15:42.94" />
                    <SPLIT distance="1100" swimtime="00:16:29.28" />
                    <SPLIT distance="1150" swimtime="00:17:16.21" />
                    <SPLIT distance="1200" swimtime="00:18:02.39" />
                    <SPLIT distance="1250" swimtime="00:18:48.54" />
                    <SPLIT distance="1300" swimtime="00:19:35.47" />
                    <SPLIT distance="1350" swimtime="00:20:21.77" />
                    <SPLIT distance="1400" swimtime="00:21:08.08" />
                    <SPLIT distance="1450" swimtime="00:21:53.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="329" reactiontime="+76" swimtime="00:00:32.73" resultid="5868" heatid="7454" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1336" points="232" reactiontime="+103" swimtime="00:02:57.33" resultid="5869" heatid="7568" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                    <SPLIT distance="100" swimtime="00:01:23.82" />
                    <SPLIT distance="150" swimtime="00:02:09.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="312" reactiontime="+92" swimtime="00:00:32.13" resultid="5870" heatid="7633" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1470" points="286" reactiontime="+79" swimtime="00:01:14.28" resultid="5871" heatid="7669" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="5872" heatid="7770" lane="4" entrytime="00:02:40.00" />
                <RESULT eventid="1710" points="277" reactiontime="+104" swimtime="00:05:26.28" resultid="5873" heatid="8052" lane="6" entrytime="00:05:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:12.33" />
                    <SPLIT distance="150" swimtime="00:01:53.53" />
                    <SPLIT distance="200" swimtime="00:02:36.03" />
                    <SPLIT distance="250" swimtime="00:03:19.23" />
                    <SPLIT distance="300" swimtime="00:04:02.35" />
                    <SPLIT distance="350" swimtime="00:04:45.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="5874">
              <RESULTS>
                <RESULT eventid="1200" points="72" reactiontime="+73" swimtime="00:00:54.19" resultid="5875" heatid="7444" lane="3" entrytime="00:00:51.20" />
                <RESULT eventid="1234" points="93" reactiontime="+110" swimtime="00:04:25.75" resultid="5876" heatid="7472" lane="4" entrytime="00:04:15.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.02" />
                    <SPLIT distance="100" swimtime="00:02:00.59" />
                    <SPLIT distance="150" swimtime="00:03:13.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="104" reactiontime="+101" swimtime="00:01:58.14" resultid="5877" heatid="7595" lane="6" entrytime="00:01:50.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="52" reactiontime="+82" swimtime="00:02:10.88" resultid="5878" heatid="7661" lane="2" entrytime="00:02:05.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="5879" heatid="7792" lane="2" entrytime="00:00:48.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowki" nation="POL" athleteid="5880">
              <RESULTS>
                <RESULT eventid="1234" points="63" reactiontime="+124" swimtime="00:05:02.44" resultid="5881" heatid="7472" lane="2" entrytime="00:04:16.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.18" />
                    <SPLIT distance="100" swimtime="00:02:31.40" />
                    <SPLIT distance="150" swimtime="00:03:47.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="73" reactiontime="+112" swimtime="00:03:57.71" resultid="5883" heatid="7689" lane="1" entrytime="00:03:29.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.16" />
                    <SPLIT distance="100" swimtime="00:01:53.44" />
                    <SPLIT distance="150" swimtime="00:02:56.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" status="DNS" swimtime="00:00:00.00" resultid="5884" heatid="7975" lane="1" entrytime="00:09:31.51" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5885" heatid="7737" lane="6" entrytime="00:02:09.68" />
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="5886" heatid="7762" lane="5" entrytime="00:04:52.58" />
                <RESULT eventid="1336" status="DNS" swimtime="00:00:00.00" resultid="7937" heatid="7564" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="Osóbka" nation="POL" athleteid="5887">
              <RESULTS>
                <RESULT eventid="1268" points="13" reactiontime="+115" swimtime="00:03:10.36" resultid="5888" heatid="7500" lane="3" entrytime="00:02:50.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K-12 - zmiana pozycji ciała (odbicie od dna)" eventid="1402" reactiontime="+119" status="DSQ" swimtime="00:03:53.07" resultid="5889" heatid="7593" lane="3" entrytime="00:03:10.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="5890" heatid="7789" lane="3" entrytime="00:01:24.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="5891">
              <RESULTS>
                <RESULT eventid="1200" points="43" reactiontime="+83" swimtime="00:01:04.10" resultid="5892" heatid="7443" lane="5" entrytime="00:00:59.42" />
                <RESULT eventid="1268" points="97" reactiontime="+112" swimtime="00:01:37.56" resultid="5893" heatid="7502" lane="2" entrytime="00:01:35.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="5894" heatid="7624" lane="1" entrytime="00:00:59.64" />
                <RESULT eventid="1470" points="45" reactiontime="+76" swimtime="00:02:16.65" resultid="5895" heatid="7661" lane="5" entrytime="00:02:12.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="5896" heatid="7762" lane="1" entrytime="00:04:58.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="5897">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5898" heatid="7354" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="5899" heatid="7393" lane="3" entrytime="00:03:55.00" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="5900" heatid="7473" lane="4" entrytime="00:03:45.00" />
                <RESULT eventid="1336" status="DNS" swimtime="00:00:00.00" resultid="5901" heatid="7568" lane="6" entrytime="00:03:15.00" />
                <RESULT eventid="1436" points="279" reactiontime="+90" swimtime="00:00:33.33" resultid="5902" heatid="7629" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5904" heatid="7742" lane="3" entrytime="00:01:22.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-03" firstname="Artur" gender="M" lastname="Kłosiński" nation="POL" athleteid="5906">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5907" heatid="7346" lane="3" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="5908" heatid="7403" lane="1" entrytime="00:02:38.00" />
                <RESULT eventid="1200" points="292" reactiontime="+76" swimtime="00:00:34.05" resultid="5909" heatid="7442" lane="5" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="5910" heatid="7481" lane="2" entrytime="00:02:55.00" />
                <RESULT eventid="1402" points="300" reactiontime="+87" swimtime="00:01:22.98" resultid="5911" heatid="7592" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="263" reactiontime="+72" swimtime="00:01:16.38" resultid="5912" heatid="7670" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="5913" heatid="7762" lane="4" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="5914" heatid="7807" lane="2" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-27" firstname="Magdalena" gender="F" lastname="Rogozińska" nation="POL" athleteid="5915">
              <RESULTS>
                <RESULT eventid="1217" points="280" reactiontime="+99" swimtime="00:03:25.65" resultid="5916" heatid="7466" lane="1" entrytime="00:03:34.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.48" />
                    <SPLIT distance="100" swimtime="00:01:40.52" />
                    <SPLIT distance="150" swimtime="00:02:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="305" reactiontime="+101" swimtime="00:01:25.77" resultid="5917" heatid="7529" lane="3" entrytime="00:01:30.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="286" reactiontime="+104" swimtime="00:01:35.09" resultid="5918" heatid="7587" lane="2" entrytime="00:01:37.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="210" reactiontime="+113" swimtime="00:00:40.96" resultid="5919" heatid="7614" lane="3" entrytime="00:00:42.70" />
                <RESULT eventid="1645" points="302" reactiontime="+97" swimtime="00:00:42.89" resultid="5920" heatid="7783" lane="1" entrytime="00:00:44.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-10-22" firstname="Magdalena" gender="F" lastname="Bolewska" nation="POL" athleteid="5921">
              <RESULTS>
                <RESULT eventid="1217" points="440" reactiontime="+88" swimtime="00:02:56.88" resultid="5922" heatid="7469" lane="2" entrytime="00:02:54.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:24.28" />
                    <SPLIT distance="150" swimtime="00:02:10.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="429" reactiontime="+83" swimtime="00:01:16.51" resultid="5923" heatid="7535" lane="2" entrytime="00:01:16.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="459" swimtime="00:01:21.26" resultid="5924" heatid="7591" lane="5" entrytime="00:01:21.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="395" reactiontime="+82" swimtime="00:00:33.22" resultid="5925" heatid="7620" lane="3" entrytime="00:00:32.80" />
                <RESULT eventid="1577" points="377" reactiontime="+88" swimtime="00:01:16.14" resultid="5926" heatid="7734" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="459" swimtime="00:00:37.33" resultid="5927" heatid="7787" lane="5" entrytime="00:00:37.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Jarosław" gender="M" lastname="Wysocki" nation="POL" athleteid="5928">
              <RESULTS>
                <RESULT eventid="1109" points="145" reactiontime="+89" swimtime="00:03:29.09" resultid="5929" heatid="7390" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:38.75" />
                    <SPLIT distance="150" swimtime="00:02:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="173" reactiontime="+90" swimtime="00:03:36.52" resultid="5930" heatid="7470" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                    <SPLIT distance="100" swimtime="00:01:43.38" />
                    <SPLIT distance="150" swimtime="00:02:40.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="129" reactiontime="+93" swimtime="00:03:35.84" resultid="5931" heatid="7565" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.26" />
                    <SPLIT distance="100" swimtime="00:01:39.13" />
                    <SPLIT distance="150" swimtime="00:02:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="171" reactiontime="+88" swimtime="00:01:40.07" resultid="5932" heatid="7593" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="134" reactiontime="+85" swimtime="00:07:39.39" resultid="5933" heatid="7974" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                    <SPLIT distance="100" swimtime="00:01:40.77" />
                    <SPLIT distance="150" swimtime="00:02:45.16" />
                    <SPLIT distance="200" swimtime="00:03:46.50" />
                    <SPLIT distance="250" swimtime="00:04:48.57" />
                    <SPLIT distance="300" swimtime="00:05:50.76" />
                    <SPLIT distance="350" swimtime="00:06:47.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="208" reactiontime="+86" swimtime="00:00:42.55" resultid="5934" heatid="7788" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="5935">
              <RESULTS>
                <RESULT eventid="1075" points="253" swimtime="00:00:32.09" resultid="5936" heatid="7358" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1109" points="166" swimtime="00:03:19.91" resultid="5937" heatid="7396" lane="5" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:39.78" />
                    <SPLIT distance="150" swimtime="00:02:38.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="238" reactiontime="+80" swimtime="00:01:12.51" resultid="5938" heatid="7508" lane="4" entrytime="00:01:11.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="205" swimtime="00:01:26.07" resultid="5939" heatid="7545" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="210" swimtime="00:00:36.67" resultid="5940" heatid="7631" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1504" points="206" reactiontime="+83" swimtime="00:02:48.13" resultid="5941" heatid="7691" lane="3" entrytime="00:02:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:01:22.80" />
                    <SPLIT distance="150" swimtime="00:02:07.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="158" swimtime="00:01:29.60" resultid="5942" heatid="7741" lane="5" entrytime="00:01:27.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="189" reactiontime="+94" swimtime="00:06:10.73" resultid="5943" heatid="8048" lane="1" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:24.64" />
                    <SPLIT distance="150" swimtime="00:02:11.83" />
                    <SPLIT distance="200" swimtime="00:03:00.14" />
                    <SPLIT distance="250" swimtime="00:03:49.58" />
                    <SPLIT distance="300" swimtime="00:04:38.62" />
                    <SPLIT distance="350" swimtime="00:05:27.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-19" firstname="Tomasz" gender="M" lastname="Zasadowski" nation="POL" athleteid="5944">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5945" heatid="7364" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1200" points="273" reactiontime="+69" swimtime="00:00:34.85" resultid="5946" heatid="7454" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1302" points="298" reactiontime="+93" swimtime="00:01:15.91" resultid="5947" heatid="7538" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="308" reactiontime="+91" swimtime="00:00:32.28" resultid="5948" heatid="7634" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="5949" heatid="7665" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1594" points="234" reactiontime="+93" swimtime="00:01:18.61" resultid="5950" heatid="7743" lane="3" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-04" firstname="Karol" gender="M" lastname="Twarowski" nation="POL" athleteid="5951">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5952" heatid="7345" lane="3" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="5953" heatid="7391" lane="5" />
                <RESULT eventid="1200" points="378" reactiontime="+82" swimtime="00:00:31.27" resultid="5954" heatid="7442" lane="4" />
                <RESULT eventid="1268" points="458" reactiontime="+87" swimtime="00:00:58.26" resultid="5955" heatid="7500" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="376" reactiontime="+72" swimtime="00:01:07.78" resultid="5956" heatid="7660" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="5958" heatid="7737" lane="5" />
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="5959" heatid="7762" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-06" firstname="Andzrej" gender="M" lastname="Szufarski" nation="POL" athleteid="5960">
              <RESULTS>
                <RESULT eventid="1109" points="118" reactiontime="+84" swimtime="00:03:43.94" resultid="5961" heatid="7394" lane="3" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:01:42.83" />
                    <SPLIT distance="150" swimtime="00:02:45.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="86" reactiontime="+85" swimtime="00:00:51.14" resultid="5962" heatid="7445" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1302" points="138" reactiontime="+103" swimtime="00:01:38.20" resultid="5963" heatid="7541" lane="2" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="128" reactiontime="+104" swimtime="00:00:43.19" resultid="5964" heatid="7626" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1559" points="109" reactiontime="+103" swimtime="00:08:12.04" resultid="5965" heatid="7976" lane="1" entrytime="00:07:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.79" />
                    <SPLIT distance="100" swimtime="00:01:54.86" />
                    <SPLIT distance="150" swimtime="00:03:02.55" />
                    <SPLIT distance="200" swimtime="00:04:05.58" />
                    <SPLIT distance="250" swimtime="00:05:10.27" />
                    <SPLIT distance="300" swimtime="00:06:17.71" />
                    <SPLIT distance="350" swimtime="00:07:16.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="84" reactiontime="+105" swimtime="00:01:50.53" resultid="5966" heatid="7740" lane="1" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="139" reactiontime="+101" swimtime="00:00:48.67" resultid="5967" heatid="7793" lane="1" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="5968">
              <RESULTS>
                <RESULT eventid="1058" points="446" reactiontime="+92" swimtime="00:00:30.42" resultid="5969" heatid="7342" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1092" points="414" reactiontime="+90" swimtime="00:02:47.10" resultid="5970" heatid="7387" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:01:18.27" />
                    <SPLIT distance="150" swimtime="00:02:05.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="382" reactiontime="+92" swimtime="00:03:05.34" resultid="5971" heatid="7466" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                    <SPLIT distance="100" swimtime="00:01:30.20" />
                    <SPLIT distance="150" swimtime="00:02:17.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="430" reactiontime="+92" swimtime="00:01:16.46" resultid="5972" heatid="7533" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="402" reactiontime="+84" swimtime="00:01:24.92" resultid="5973" heatid="7588" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="377" reactiontime="+85" swimtime="00:00:33.73" resultid="5974" heatid="7620" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1577" points="368" reactiontime="+78" swimtime="00:01:16.77" resultid="5975" heatid="7734" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="395" reactiontime="+68" swimtime="00:00:39.25" resultid="5976" heatid="7784" lane="3" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-07-25" firstname="Sławomir" gender="M" lastname="Prędki" nation="POL" athleteid="5977">
              <RESULTS>
                <RESULT eventid="1075" points="520" reactiontime="+79" swimtime="00:00:25.24" resultid="5978" heatid="7345" lane="4" />
                <RESULT eventid="1109" points="531" reactiontime="+86" swimtime="00:02:15.87" resultid="5979" heatid="7390" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                    <SPLIT distance="150" swimtime="00:01:43.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="508" reactiontime="+87" swimtime="00:02:31.14" resultid="5980" heatid="7471" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                    <SPLIT distance="150" swimtime="00:01:50.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="545" reactiontime="+85" swimtime="00:01:02.14" resultid="5981" heatid="7538" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1402" points="535" swimtime="00:01:08.46" resultid="5982" heatid="7593" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="520" swimtime="00:02:03.57" resultid="5983" heatid="7686" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                    <SPLIT distance="100" swimtime="00:01:00.14" />
                    <SPLIT distance="150" swimtime="00:01:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1662" points="519" reactiontime="+84" swimtime="00:00:31.41" resultid="5984" heatid="7788" lane="3" />
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="5985" heatid="8044" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="319" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="76" reactiontime="+80" swimtime="00:03:35.85" resultid="5986" heatid="7929" lane="4" entrytime="00:03:41.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.45" />
                    <SPLIT distance="100" swimtime="00:01:19.25" />
                    <SPLIT distance="150" swimtime="00:02:36.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5874" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5887" number="2" reactiontime="+121" />
                    <RELAYPOSITION athleteid="5880" number="3" />
                    <RELAYPOSITION athleteid="5891" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1528" points="57" swimtime="00:03:28.78" resultid="7997" heatid="7709" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.89" />
                    <SPLIT distance="100" swimtime="00:01:59.77" />
                    <SPLIT distance="150" swimtime="00:02:04.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1377" points="372" reactiontime="+72" swimtime="00:02:07.56" resultid="5989" heatid="7933" lane="6" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:03.42" />
                    <SPLIT distance="150" swimtime="00:01:39.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5906" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="5977" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="5935" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5951" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="5990" heatid="7714" lane="6" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5906" number="1" />
                    <RELAYPOSITION athleteid="5935" number="2" />
                    <RELAYPOSITION athleteid="5951" number="3" />
                    <RELAYPOSITION athleteid="5977" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1377" points="305" reactiontime="+74" swimtime="00:02:16.34" resultid="5991" heatid="7932" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:01:48.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5865" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="5897" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="5944" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="5859" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="5992" heatid="7713" lane="4" entrytime="00:01:57.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5897" number="1" />
                    <RELAYPOSITION athleteid="5944" number="2" />
                    <RELAYPOSITION athleteid="5859" number="3" />
                    <RELAYPOSITION athleteid="5865" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1679" points="379" reactiontime="+72" swimtime="00:02:06.81" resultid="5988" heatid="7819" lane="4" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:03.29" />
                    <SPLIT distance="150" swimtime="00:01:36.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5865" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="5977" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="5968" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="5921" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Redeco Wrocław" nation="POL" region="DOL">
          <CONTACT city="Wrocław" name="Wolny Dariusz" phone="603630870" state="DOL" street="Rogowska 52a" zip="54-440" />
          <ATHLETES>
            <ATHLETE birthdate="1960-03-21" firstname="Dariusz" gender="M" lastname="Wolny" nation="POL" athleteid="6016">
              <RESULTS>
                <RESULT eventid="1109" points="429" reactiontime="+83" swimtime="00:02:25.94" resultid="6017" heatid="7404" lane="2" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:07.52" />
                    <SPLIT distance="150" swimtime="00:01:51.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="406" reactiontime="+67" swimtime="00:00:30.52" resultid="6018" heatid="7455" lane="2" entrytime="00:00:31.31" />
                <RESULT eventid="1302" points="420" reactiontime="+77" swimtime="00:01:07.73" resultid="6019" heatid="7555" lane="6" entrytime="00:01:08.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="396" reactiontime="+66" swimtime="00:01:06.63" resultid="6020" heatid="7671" lane="2" entrytime="00:01:08.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-13" firstname="Kazimiera" gender="F" lastname="Syguła" nation="POL" athleteid="6021">
              <RESULTS>
                <RESULT eventid="1092" points="126" reactiontime="+108" swimtime="00:04:08.43" resultid="6022" heatid="7384" lane="6" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.22" />
                    <SPLIT distance="100" swimtime="00:01:56.90" />
                    <SPLIT distance="150" swimtime="00:03:08.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="127" reactiontime="+115" swimtime="00:01:54.70" resultid="6023" heatid="7527" lane="1" entrytime="00:01:57.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="110" reactiontime="+70" swimtime="00:01:54.94" resultid="6024" heatid="7650" lane="2" entrytime="00:01:53.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="121" reactiontime="+78" swimtime="00:04:02.05" resultid="6025" heatid="7756" lane="6" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.08" />
                    <SPLIT distance="100" swimtime="00:01:57.43" />
                    <SPLIT distance="150" swimtime="00:03:00.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-11-30" firstname="Ryszard" gender="M" lastname="Sowiński" nation="POL" athleteid="6026">
              <RESULTS>
                <RESULT eventid="1165" points="81" swimtime="00:32:40.87" resultid="6027" heatid="7908" lane="1" entrytime="00:31:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.17" />
                    <SPLIT distance="100" swimtime="00:02:17.41" />
                    <SPLIT distance="150" swimtime="00:03:22.25" />
                    <SPLIT distance="200" swimtime="00:04:26.97" />
                    <SPLIT distance="250" swimtime="00:05:31.13" />
                    <SPLIT distance="300" swimtime="00:06:36.82" />
                    <SPLIT distance="350" swimtime="00:07:40.97" />
                    <SPLIT distance="400" swimtime="00:08:47.36" />
                    <SPLIT distance="450" swimtime="00:09:53.90" />
                    <SPLIT distance="500" swimtime="00:10:59.91" />
                    <SPLIT distance="550" swimtime="00:12:04.82" />
                    <SPLIT distance="600" swimtime="00:13:12.11" />
                    <SPLIT distance="650" swimtime="00:14:18.56" />
                    <SPLIT distance="700" swimtime="00:15:22.50" />
                    <SPLIT distance="750" swimtime="00:16:26.43" />
                    <SPLIT distance="800" swimtime="00:17:32.73" />
                    <SPLIT distance="850" swimtime="00:18:37.63" />
                    <SPLIT distance="900" swimtime="00:19:41.64" />
                    <SPLIT distance="950" swimtime="00:20:48.14" />
                    <SPLIT distance="1000" swimtime="00:21:53.84" />
                    <SPLIT distance="1050" swimtime="00:22:58.46" />
                    <SPLIT distance="1100" swimtime="00:24:03.63" />
                    <SPLIT distance="1150" swimtime="00:25:07.33" />
                    <SPLIT distance="1200" swimtime="00:26:13.55" />
                    <SPLIT distance="1250" swimtime="00:27:18.07" />
                    <SPLIT distance="1300" swimtime="00:28:22.56" />
                    <SPLIT distance="1350" swimtime="00:29:28.34" />
                    <SPLIT distance="1400" swimtime="00:30:33.45" />
                    <SPLIT distance="1450" swimtime="00:31:39.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-09-26" firstname="Rafał" gender="M" lastname="Rogoza" nation="POL" athleteid="6028">
              <RESULTS>
                <RESULT eventid="1075" points="270" reactiontime="+83" swimtime="00:00:31.39" resultid="6029" heatid="7354" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1268" points="214" reactiontime="+87" swimtime="00:01:15.10" resultid="6030" heatid="7507" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="212" reactiontime="+84" swimtime="00:01:25.05" resultid="6031" heatid="7547" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="268" reactiontime="+89" swimtime="00:00:33.79" resultid="6032" heatid="7628" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1594" points="182" reactiontime="+106" swimtime="00:01:25.42" resultid="6033" heatid="7742" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="145" swimtime="00:00:47.96" resultid="6034" heatid="7794" lane="5" entrytime="00:00:44.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-13" firstname="Małgorzata" gender="F" lastname="Bołtuć" nation="POL" athleteid="6035">
              <RESULTS>
                <RESULT eventid="1058" points="163" reactiontime="+101" swimtime="00:00:42.50" resultid="6036" heatid="7334" lane="1" entrytime="00:00:46.88" />
                <RESULT eventid="1092" points="179" reactiontime="+102" swimtime="00:03:40.72" resultid="6037" heatid="7384" lane="2" entrytime="00:03:44.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.85" />
                    <SPLIT distance="100" swimtime="00:02:51.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="183" reactiontime="+101" swimtime="00:03:56.68" resultid="6038" heatid="7464" lane="2" entrytime="00:04:01.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.36" />
                    <SPLIT distance="100" swimtime="00:01:58.84" />
                    <SPLIT distance="150" swimtime="00:02:58.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="164" swimtime="00:01:33.10" resultid="6039" heatid="7488" lane="5" entrytime="00:01:41.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="174" swimtime="00:01:52.15" resultid="6040" heatid="7584" lane="5" entrytime="00:01:52.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="110" reactiontime="+182" swimtime="00:00:50.83" resultid="6041" heatid="7614" lane="2" entrytime="00:00:48.88" />
                <RESULT eventid="1645" points="178" reactiontime="+103" swimtime="00:00:51.11" resultid="6042" heatid="7780" lane="6" entrytime="00:00:49.75" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-12-13" firstname="Agata" gender="F" lastname="Grochowska" nation="POL" athleteid="6043">
              <RESULTS>
                <RESULT eventid="1092" points="187" reactiontime="+82" swimtime="00:03:37.87" resultid="6044" heatid="7384" lane="4" entrytime="00:03:39.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:42.24" />
                    <SPLIT distance="150" swimtime="00:02:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="194" reactiontime="+60" swimtime="00:00:44.37" resultid="6045" heatid="7434" lane="2" entrytime="00:00:45.07" />
                <RESULT eventid="1285" points="214" reactiontime="+87" swimtime="00:01:36.51" resultid="6046" heatid="7528" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="187" reactiontime="+88" swimtime="00:01:49.53" resultid="6047" heatid="7588" lane="6" entrytime="00:01:33.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="170" reactiontime="+61" swimtime="00:01:39.66" resultid="6048" heatid="7651" lane="6" entrytime="00:01:38.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:39.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="6049" heatid="7784" lane="6" entrytime="00:00:43.43" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-27" firstname="Hanna" gender="F" lastname="Sikacz" nation="POL" athleteid="6051">
              <RESULTS>
                <RESULT eventid="1058" points="297" reactiontime="+83" swimtime="00:00:34.83" resultid="6052" heatid="7336" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1148" points="256" reactiontime="+89" swimtime="00:12:42.36" resultid="6053" heatid="7904" lane="2" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:27.31" />
                    <SPLIT distance="150" swimtime="00:02:13.89" />
                    <SPLIT distance="200" swimtime="00:03:00.66" />
                    <SPLIT distance="250" swimtime="00:03:49.54" />
                    <SPLIT distance="300" swimtime="00:04:37.74" />
                    <SPLIT distance="350" swimtime="00:05:26.48" />
                    <SPLIT distance="400" swimtime="00:06:15.19" />
                    <SPLIT distance="450" swimtime="00:07:03.73" />
                    <SPLIT distance="500" swimtime="00:07:52.19" />
                    <SPLIT distance="550" swimtime="00:08:42.27" />
                    <SPLIT distance="600" swimtime="00:09:30.55" />
                    <SPLIT distance="650" swimtime="00:10:20.47" />
                    <SPLIT distance="700" swimtime="00:11:09.29" />
                    <SPLIT distance="750" swimtime="00:11:57.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="279" reactiontime="+82" swimtime="00:01:17.98" resultid="6054" heatid="7493" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="288" reactiontime="+89" swimtime="00:01:27.36" resultid="6055" heatid="7530" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="280" reactiontime="+81" swimtime="00:02:49.73" resultid="6056" heatid="7681" lane="4" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="100" swimtime="00:01:19.76" />
                    <SPLIT distance="150" swimtime="00:02:05.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" status="DNS" swimtime="00:00:00.00" resultid="6058" heatid="7757" lane="4" entrytime="00:03:13.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-01" firstname="Wojciech" gender="M" lastname="Dobrowolski" nation="POL" athleteid="6060">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="6061" heatid="7370" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="6062" heatid="7517" lane="4" entrytime="00:01:03.00" />
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="6063" heatid="7635" lane="1" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-03-25" firstname="Krzysztof" gender="M" lastname="Gajewski" nation="POL" athleteid="6064">
              <RESULTS>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start), Przekroczony limit czasu." eventid="1165" reactiontime="+73" status="DSQ" swimtime="00:23:50.62" resultid="6065" heatid="7912" lane="4" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:17.04" />
                    <SPLIT distance="150" swimtime="00:02:02.10" />
                    <SPLIT distance="200" swimtime="00:02:47.14" />
                    <SPLIT distance="250" swimtime="00:03:32.95" />
                    <SPLIT distance="300" swimtime="00:04:19.44" />
                    <SPLIT distance="350" swimtime="00:05:06.63" />
                    <SPLIT distance="400" swimtime="00:05:54.41" />
                    <SPLIT distance="450" swimtime="00:06:42.29" />
                    <SPLIT distance="500" swimtime="00:07:30.68" />
                    <SPLIT distance="550" swimtime="00:08:19.14" />
                    <SPLIT distance="600" swimtime="00:09:07.79" />
                    <SPLIT distance="650" swimtime="00:09:56.79" />
                    <SPLIT distance="700" swimtime="00:10:46.04" />
                    <SPLIT distance="750" swimtime="00:11:35.39" />
                    <SPLIT distance="800" swimtime="00:12:24.56" />
                    <SPLIT distance="850" swimtime="00:13:13.29" />
                    <SPLIT distance="900" swimtime="00:14:02.32" />
                    <SPLIT distance="950" swimtime="00:14:51.01" />
                    <SPLIT distance="1000" swimtime="00:15:40.03" />
                    <SPLIT distance="1050" swimtime="00:16:29.49" />
                    <SPLIT distance="1100" swimtime="00:17:19.21" />
                    <SPLIT distance="1150" swimtime="00:18:08.26" />
                    <SPLIT distance="1200" swimtime="00:18:58.67" />
                    <SPLIT distance="1250" swimtime="00:19:47.14" />
                    <SPLIT distance="1300" swimtime="00:20:36.98" />
                    <SPLIT distance="1350" swimtime="00:21:26.15" />
                    <SPLIT distance="1400" swimtime="00:22:15.14" />
                    <SPLIT distance="1450" swimtime="00:23:03.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-14" firstname="Anna" gender="F" lastname="Jaśkiewicz" nation="POL" athleteid="7067">
              <RESULTS>
                <RESULT eventid="1092" points="241" swimtime="00:03:20.12" resultid="7068" heatid="7385" lane="5" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                    <SPLIT distance="100" swimtime="00:01:37.08" />
                    <SPLIT distance="150" swimtime="00:02:34.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="213" reactiontime="+90" swimtime="00:13:31.28" resultid="7069" heatid="7903" lane="3" entrytime="00:13:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:01:29.10" />
                    <SPLIT distance="150" swimtime="00:02:19.08" />
                    <SPLIT distance="200" swimtime="00:03:09.58" />
                    <SPLIT distance="250" swimtime="00:04:01.21" />
                    <SPLIT distance="300" swimtime="00:04:53.21" />
                    <SPLIT distance="350" swimtime="00:05:45.78" />
                    <SPLIT distance="400" swimtime="00:06:38.09" />
                    <SPLIT distance="450" swimtime="00:07:30.11" />
                    <SPLIT distance="500" swimtime="00:08:22.41" />
                    <SPLIT distance="550" swimtime="00:09:14.83" />
                    <SPLIT distance="600" swimtime="00:10:07.37" />
                    <SPLIT distance="650" swimtime="00:10:59.84" />
                    <SPLIT distance="700" swimtime="00:11:51.79" />
                    <SPLIT distance="750" swimtime="00:12:43.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="269" reactiontime="+98" swimtime="00:03:28.37" resultid="7070" heatid="7467" lane="6" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                    <SPLIT distance="100" swimtime="00:01:39.86" />
                    <SPLIT distance="150" swimtime="00:02:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="271" reactiontime="+91" swimtime="00:01:18.80" resultid="7071" heatid="7491" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="286" reactiontime="+87" swimtime="00:01:35.09" resultid="7072" heatid="7587" lane="1" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="241" reactiontime="+83" swimtime="00:02:58.48" resultid="7073" heatid="7679" lane="3" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:25.56" />
                    <SPLIT distance="150" swimtime="00:02:08.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="290" swimtime="00:00:43.51" resultid="7074" heatid="7782" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="1693" points="219" reactiontime="+82" swimtime="00:06:29.71" resultid="7075" heatid="8021" lane="6" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:01:26.37" />
                    <SPLIT distance="150" swimtime="00:02:16.74" />
                    <SPLIT distance="200" swimtime="00:03:07.17" />
                    <SPLIT distance="250" swimtime="00:03:58.29" />
                    <SPLIT distance="300" swimtime="00:04:49.30" />
                    <SPLIT distance="350" swimtime="00:05:40.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-25" firstname="Marlena" gender="F" lastname="Jakubów" nation="POL" athleteid="7243">
              <RESULTS>
                <RESULT eventid="1092" points="207" reactiontime="+115" swimtime="00:03:30.36" resultid="7244" heatid="7385" lane="1" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:40.21" />
                    <SPLIT distance="150" swimtime="00:02:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="196" reactiontime="+119" swimtime="00:13:53.96" resultid="7245" heatid="7903" lane="6" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="100" swimtime="00:01:36.09" />
                    <SPLIT distance="150" swimtime="00:02:28.26" />
                    <SPLIT distance="200" swimtime="00:03:21.08" />
                    <SPLIT distance="250" swimtime="00:04:15.44" />
                    <SPLIT distance="300" swimtime="00:05:07.36" />
                    <SPLIT distance="350" swimtime="00:05:59.93" />
                    <SPLIT distance="400" swimtime="00:06:53.26" />
                    <SPLIT distance="450" swimtime="00:07:45.86" />
                    <SPLIT distance="500" swimtime="00:08:38.90" />
                    <SPLIT distance="550" swimtime="00:09:33.38" />
                    <SPLIT distance="600" swimtime="00:10:26.89" />
                    <SPLIT distance="650" swimtime="00:11:19.58" />
                    <SPLIT distance="700" swimtime="00:12:11.57" />
                    <SPLIT distance="750" swimtime="00:13:03.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="189" reactiontime="+97" swimtime="00:00:44.71" resultid="7246" heatid="7435" lane="1" entrytime="00:00:44.40" />
                <RESULT eventid="1251" points="237" reactiontime="+121" swimtime="00:01:22.39" resultid="7247" heatid="7492" lane="3" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="179" reactiontime="+104" swimtime="00:01:37.86" resultid="7248" heatid="7651" lane="5" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="198" reactiontime="+119" swimtime="00:03:10.67" resultid="7249" heatid="7679" lane="6" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:01:28.98" />
                    <SPLIT distance="150" swimtime="00:02:21.05" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G-3 - Wynurzenie głowy spod lustra wody po starcie poza 15m" eventid="1611" reactiontime="+108" status="DSQ" swimtime="00:03:46.10" resultid="7250" heatid="7756" lane="1" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                    <SPLIT distance="100" swimtime="00:01:47.12" />
                    <SPLIT distance="150" swimtime="00:02:47.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1693" points="185" reactiontime="+126" swimtime="00:06:52.18" resultid="7251" heatid="8021" lane="1" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                    <SPLIT distance="100" swimtime="00:01:33.09" />
                    <SPLIT distance="150" swimtime="00:02:26.34" />
                    <SPLIT distance="200" swimtime="00:03:20.95" />
                    <SPLIT distance="250" swimtime="00:04:17.61" />
                    <SPLIT distance="300" swimtime="00:05:11.67" />
                    <SPLIT distance="350" swimtime="00:06:04.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Masters rzeszów" nation="POL">
          <CONTACT city="Rzeszów" email="wieslawcieklinski@wp.pl" name="Ciekliński Wiesław" phone="602682904" state="PODK" street="Jagiellońska 7/3" zip="35-25" />
          <ATHLETES>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="6067">
              <RESULTS>
                <RESULT eventid="1075" points="264" reactiontime="+91" swimtime="00:00:31.61" resultid="6068" heatid="7358" lane="4" entrytime="00:00:32.00" />
                <RESULT comment="K-14" eventid="1109" reactiontime="+124" status="DSQ" swimtime="00:03:26.70" resultid="6069" heatid="7396" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                    <SPLIT distance="100" swimtime="00:01:44.97" />
                    <SPLIT distance="150" swimtime="00:02:45.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="249" reactiontime="+96" swimtime="00:01:11.38" resultid="6070" heatid="7508" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="171" reactiontime="+92" swimtime="00:01:31.29" resultid="6071" heatid="7543" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="175" reactiontime="+86" swimtime="00:00:38.92" resultid="6072" heatid="7628" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1504" points="209" reactiontime="+107" swimtime="00:02:47.24" resultid="6073" heatid="7693" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:20.81" />
                    <SPLIT distance="150" swimtime="00:02:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="184" reactiontime="+114" swimtime="00:06:13.53" resultid="6074" heatid="8049" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:03:52.28" />
                    <SPLIT distance="150" swimtime="00:04:40.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="AQUA Masters Kiev" nation="UKR">
          <ATHLETES>
            <ATHLETE birthdate="1959-01-01" firstname="Sergii" gender="M" lastname="Fesenko " nation="POL" athleteid="6103">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1200" points="369" reactiontime="+71" swimtime="00:00:31.51" resultid="6104" heatid="7454" lane="6" entrytime="00:00:33.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1302" points="407" reactiontime="+89" swimtime="00:01:08.48" resultid="6105" heatid="7554" lane="1" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1436" points="386" reactiontime="+89" swimtime="00:00:29.93" resultid="6106" heatid="7639" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1504" points="356" reactiontime="+85" swimtime="00:02:20.16" resultid="6107" heatid="7700" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="336" reactiontime="+86" swimtime="00:01:09.70" resultid="6108" heatid="7748" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="319" reactiontime="+76" swimtime="00:02:35.24" resultid="6109" heatid="7770" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                    <SPLIT distance="100" swimtime="00:01:17.43" />
                    <SPLIT distance="150" swimtime="00:01:56.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Volodymyr " gender="M" lastname="Brykov " nation="UKR" athleteid="6110">
              <RESULTS>
                <RESULT comment="K-2 - Brak wynurzenia głowy po rozpoczeciu ruchuramion do wewnątrz z jego najszerszego położenia w drugim cyklu ruchu ramion po starcie" eventid="1402" reactiontime="+139" status="DSQ" swimtime="00:02:25.83" resultid="6111" heatid="7592" lane="1" entrytime="00:01:00.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="6112" heatid="7485" lane="3" entrytime="00:02:00.30" />
                <RESULT eventid="1662" points="64" reactiontime="+124" swimtime="00:01:03.01" resultid="8005" heatid="7788" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Petro " gender="M" lastname="Gemba" nation="UKR" athleteid="6113">
              <RESULTS>
                <RESULT eventid="1165" points="237" reactiontime="+99" swimtime="00:22:53.11" resultid="6114" heatid="7912" lane="6" entrytime="00:23:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:24.92" />
                    <SPLIT distance="150" swimtime="00:02:10.36" />
                    <SPLIT distance="200" swimtime="00:02:55.69" />
                    <SPLIT distance="250" swimtime="00:03:42.25" />
                    <SPLIT distance="300" swimtime="00:04:28.67" />
                    <SPLIT distance="350" swimtime="00:05:14.96" />
                    <SPLIT distance="400" swimtime="00:06:00.98" />
                    <SPLIT distance="450" swimtime="00:06:47.53" />
                    <SPLIT distance="500" swimtime="00:07:34.48" />
                    <SPLIT distance="550" swimtime="00:08:21.53" />
                    <SPLIT distance="600" swimtime="00:09:07.44" />
                    <SPLIT distance="650" swimtime="00:09:55.02" />
                    <SPLIT distance="700" swimtime="00:10:41.25" />
                    <SPLIT distance="750" swimtime="00:11:27.56" />
                    <SPLIT distance="800" swimtime="00:12:13.80" />
                    <SPLIT distance="850" swimtime="00:13:00.32" />
                    <SPLIT distance="900" swimtime="00:13:46.03" />
                    <SPLIT distance="950" swimtime="00:14:32.21" />
                    <SPLIT distance="1000" swimtime="00:15:19.15" />
                    <SPLIT distance="1050" swimtime="00:16:03.91" />
                    <SPLIT distance="1100" swimtime="00:16:49.84" />
                    <SPLIT distance="1150" swimtime="00:17:36.00" />
                    <SPLIT distance="1200" swimtime="00:18:22.47" />
                    <SPLIT distance="1250" swimtime="00:19:09.03" />
                    <SPLIT distance="1300" swimtime="00:19:55.01" />
                    <SPLIT distance="1350" swimtime="00:20:39.86" />
                    <SPLIT distance="1400" swimtime="00:21:26.47" />
                    <SPLIT distance="1450" swimtime="00:22:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="206" reactiontime="+87" swimtime="00:01:25.88" resultid="6115" heatid="7543" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="213" swimtime="00:02:46.28" resultid="6116" heatid="7693" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:21.29" />
                    <SPLIT distance="150" swimtime="00:02:04.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="225" swimtime="00:05:49.71" resultid="8060" heatid="8043" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:26.04" />
                    <SPLIT distance="150" swimtime="00:02:10.90" />
                    <SPLIT distance="200" swimtime="00:02:55.68" />
                    <SPLIT distance="250" swimtime="00:03:41.12" />
                    <SPLIT distance="300" swimtime="00:04:25.27" />
                    <SPLIT distance="350" swimtime="00:05:09.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="PK Haviřov" nation="CZE">
          <ATHLETES>
            <ATHLETE birthdate="1972-01-01" firstname="Libor " gender="M" lastname="Hracki  " nation="POL" athleteid="6119">
              <RESULTS>
                <RESULT eventid="1234" points="291" swimtime="00:03:01.96" resultid="6120" heatid="7479" lane="5" entrytime="00:03:02.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:25.85" />
                    <SPLIT distance="150" swimtime="00:02:14.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="304" reactiontime="+82" swimtime="00:01:06.78" resultid="6121" heatid="7511" lane="4" entrytime="00:01:07.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="300" swimtime="00:01:23.04" resultid="6122" heatid="7604" lane="5" entrytime="00:01:23.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="287" reactiontime="+85" swimtime="00:02:30.55" resultid="6123" heatid="7696" lane="3" entrytime="00:02:30.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:10.38" />
                    <SPLIT distance="150" swimtime="00:01:50.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="UKS Jagiellonka Warszawa" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1982-06-03" firstname="Piotr" gender="M" lastname="Fuliński" nation="POL" athleteid="3954">
              <RESULTS>
                <RESULT eventid="1075" points="439" swimtime="00:00:26.71" resultid="3955" heatid="7378" lane="5" entrytime="00:00:26.00" />
                <RESULT eventid="1268" points="432" reactiontime="+83" swimtime="00:00:59.41" resultid="3956" heatid="7500" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="376" reactiontime="+87" swimtime="00:01:10.32" resultid="3957" heatid="7555" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="418" reactiontime="+88" swimtime="00:02:12.86" resultid="3958" heatid="7704" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="150" swimtime="00:01:37.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Zvezdy Rossii" nation="RUS">
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Natalia" gender="F" lastname="Aleshchenko " nation="RUS" athleteid="6185">
              <RESULTS>
                <RESULT eventid="1058" points="314" reactiontime="+89" swimtime="00:00:34.19" resultid="6186" heatid="7339" lane="1" entrytime="00:00:34.80" />
                <RESULT eventid="1251" points="292" swimtime="00:01:16.81" resultid="6188" heatid="7493" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="313" reactiontime="+96" swimtime="00:01:24.99" resultid="6189" heatid="7531" lane="6" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="287" reactiontime="+87" swimtime="00:00:36.92" resultid="6190" heatid="7617" lane="3" entrytime="00:00:37.80" />
                <RESULT eventid="1487" points="272" reactiontime="+97" swimtime="00:02:51.54" resultid="6191" heatid="7681" lane="1" entrytime="00:02:49.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:23.28" />
                    <SPLIT distance="150" swimtime="00:02:09.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="254" reactiontime="+88" swimtime="00:01:26.85" resultid="6192" heatid="7733" lane="2" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Irina" gender="F" lastname="Titova " nation="RUS" athleteid="6195">
              <RESULTS>
                <RESULT eventid="1058" points="293" swimtime="00:00:34.97" resultid="6196" heatid="7338" lane="5" entrytime="00:00:35.80" />
                <RESULT eventid="1251" points="304" reactiontime="+108" swimtime="00:01:15.79" resultid="6197" heatid="7493" lane="6" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="310" swimtime="00:02:44.12" resultid="6198" heatid="7681" lane="5" entrytime="00:02:49.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:01.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Marina" gender="F" lastname="Kilina " nation="RUS" athleteid="6200">
              <RESULTS>
                <RESULT eventid="1058" points="326" reactiontime="+100" swimtime="00:00:33.76" resultid="6201" heatid="7340" lane="1" entrytime="00:00:33.80" />
                <RESULT eventid="1285" points="319" reactiontime="+95" swimtime="00:01:24.46" resultid="6202" heatid="7531" lane="4" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="260" reactiontime="+75" swimtime="00:01:26.48" resultid="6203" heatid="7653" lane="2" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="255" swimtime="00:00:45.36" resultid="6204" heatid="7783" lane="5" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Elena" gender="F" lastname="Dautova " nation="RUS" athleteid="6205">
              <RESULTS>
                <RESULT eventid="1058" points="385" reactiontime="+66" swimtime="00:00:31.95" resultid="6206" heatid="7340" lane="3" entrytime="00:00:32.60" />
                <RESULT eventid="1183" points="283" swimtime="00:00:39.13" resultid="6207" heatid="7438" lane="5" entrytime="00:00:38.70" />
                <RESULT eventid="1453" points="279" reactiontime="+50" swimtime="00:01:24.45" resultid="6208" heatid="7654" lane="3" entrytime="00:01:24.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="243" reactiontime="+67" swimtime="00:03:12.32" resultid="6209" heatid="7757" lane="2" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.20" />
                    <SPLIT distance="100" swimtime="00:01:35.17" />
                    <SPLIT distance="150" swimtime="00:02:25.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Aleksandr" gender="M" lastname="Tervinskiy " nation="RUS" athleteid="6217">
              <RESULTS>
                <RESULT eventid="1200" points="172" reactiontime="+74" swimtime="00:00:40.63" resultid="6219" heatid="7446" lane="1" entrytime="00:00:42.90" />
                <RESULT eventid="1075" points="236" reactiontime="+87" swimtime="00:00:32.81" resultid="6220" heatid="7354" lane="3" entrytime="00:00:33.80" />
                <RESULT eventid="1302" points="213" swimtime="00:01:24.99" resultid="6221" heatid="7544" lane="5" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="217" reactiontime="+88" swimtime="00:01:32.53" resultid="6222" heatid="7597" lane="3" entrytime="00:01:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="266" reactiontime="+88" swimtime="00:00:39.23" resultid="6223" heatid="7795" lane="4" entrytime="00:00:42.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Sergey" gender="M" lastname="Mikhaylov " nation="RUS" athleteid="6224">
              <RESULTS>
                <RESULT eventid="1075" points="120" swimtime="00:00:41.13" resultid="6225" heatid="7350" lane="5" entrytime="00:00:39.50" />
                <RESULT eventid="1165" points="156" reactiontime="+98" swimtime="00:26:18.41" resultid="6226" heatid="7909" lane="3" entrytime="00:26:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                    <SPLIT distance="100" swimtime="00:01:35.84" />
                    <SPLIT distance="150" swimtime="00:02:27.61" />
                    <SPLIT distance="200" swimtime="00:03:19.24" />
                    <SPLIT distance="250" swimtime="00:04:10.81" />
                    <SPLIT distance="300" swimtime="00:05:02.62" />
                    <SPLIT distance="350" swimtime="00:05:55.33" />
                    <SPLIT distance="400" swimtime="00:06:47.97" />
                    <SPLIT distance="450" swimtime="00:07:39.94" />
                    <SPLIT distance="500" swimtime="00:08:32.18" />
                    <SPLIT distance="550" swimtime="00:09:25.42" />
                    <SPLIT distance="600" swimtime="00:10:18.53" />
                    <SPLIT distance="650" swimtime="00:11:10.85" />
                    <SPLIT distance="700" swimtime="00:12:03.65" />
                    <SPLIT distance="750" swimtime="00:12:56.55" />
                    <SPLIT distance="800" swimtime="00:13:50.30" />
                    <SPLIT distance="850" swimtime="00:14:43.09" />
                    <SPLIT distance="900" swimtime="00:15:36.64" />
                    <SPLIT distance="950" swimtime="00:16:30.84" />
                    <SPLIT distance="1000" swimtime="00:17:25.36" />
                    <SPLIT distance="1050" swimtime="00:18:20.13" />
                    <SPLIT distance="1100" swimtime="00:19:14.23" />
                    <SPLIT distance="1150" swimtime="00:20:09.12" />
                    <SPLIT distance="1200" swimtime="00:21:01.81" />
                    <SPLIT distance="1250" swimtime="00:21:56.32" />
                    <SPLIT distance="1300" swimtime="00:22:49.68" />
                    <SPLIT distance="1350" swimtime="00:23:43.22" />
                    <SPLIT distance="1400" swimtime="00:24:34.96" />
                    <SPLIT distance="1450" swimtime="00:25:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="128" reactiontime="+88" swimtime="00:01:29.08" resultid="6227" heatid="7503" lane="3" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="146" reactiontime="+98" swimtime="00:03:08.32" resultid="6228" heatid="7689" lane="3" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                    <SPLIT distance="100" swimtime="00:01:30.37" />
                    <SPLIT distance="150" swimtime="00:02:20.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="6229" heatid="8046" lane="3" entrytime="00:06:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Vladlen" gender="M" lastname="Nesvetaev " nation="RUS" athleteid="6230">
              <RESULTS>
                <RESULT eventid="1165" points="437" swimtime="00:18:39.77" resultid="6231" heatid="7916" lane="5" entrytime="00:18:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                    <SPLIT distance="150" swimtime="00:01:44.64" />
                    <SPLIT distance="200" swimtime="00:02:21.20" />
                    <SPLIT distance="250" swimtime="00:02:58.11" />
                    <SPLIT distance="300" swimtime="00:03:35.01" />
                    <SPLIT distance="350" swimtime="00:04:12.52" />
                    <SPLIT distance="400" swimtime="00:04:50.07" />
                    <SPLIT distance="450" swimtime="00:05:27.44" />
                    <SPLIT distance="500" swimtime="00:06:05.43" />
                    <SPLIT distance="550" swimtime="00:06:43.04" />
                    <SPLIT distance="600" swimtime="00:07:20.77" />
                    <SPLIT distance="650" swimtime="00:07:58.74" />
                    <SPLIT distance="700" swimtime="00:08:36.70" />
                    <SPLIT distance="750" swimtime="00:09:14.58" />
                    <SPLIT distance="800" swimtime="00:09:52.38" />
                    <SPLIT distance="850" swimtime="00:10:30.20" />
                    <SPLIT distance="900" swimtime="00:11:07.89" />
                    <SPLIT distance="950" swimtime="00:11:46.03" />
                    <SPLIT distance="1000" swimtime="00:12:24.02" />
                    <SPLIT distance="1050" swimtime="00:13:01.66" />
                    <SPLIT distance="1100" swimtime="00:13:39.21" />
                    <SPLIT distance="1150" swimtime="00:14:16.98" />
                    <SPLIT distance="1200" swimtime="00:14:54.95" />
                    <SPLIT distance="1250" swimtime="00:15:33.07" />
                    <SPLIT distance="1300" swimtime="00:16:11.34" />
                    <SPLIT distance="1350" swimtime="00:16:49.29" />
                    <SPLIT distance="1400" swimtime="00:17:27.22" />
                    <SPLIT distance="1450" swimtime="00:18:04.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="360" reactiontime="+80" swimtime="00:01:11.30" resultid="6232" heatid="7552" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="340" reactiontime="+85" swimtime="00:02:36.28" resultid="6233" heatid="7571" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="341" reactiontime="+76" swimtime="00:00:31.18" resultid="6234" heatid="7638" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="1559" points="384" swimtime="00:05:23.99" resultid="6235" heatid="7980" lane="5" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:54.64" />
                    <SPLIT distance="200" swimtime="00:02:36.38" />
                    <SPLIT distance="250" swimtime="00:03:24.65" />
                    <SPLIT distance="300" swimtime="00:04:11.83" />
                    <SPLIT distance="350" swimtime="00:04:48.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="389" swimtime="00:01:06.40" resultid="6236" heatid="7749" lane="5" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="6237" heatid="8056" lane="3" entrytime="00:04:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Grigoriy" gender="M" lastname="Lopin " nation="RUS" athleteid="6238">
              <RESULTS>
                <RESULT eventid="1075" points="272" reactiontime="+97" swimtime="00:00:31.30" resultid="6239" heatid="7360" lane="6" entrytime="00:00:31.40" />
                <RESULT eventid="1234" points="217" reactiontime="+98" swimtime="00:03:20.69" resultid="6240" heatid="7476" lane="6" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                    <SPLIT distance="100" swimtime="00:01:34.30" />
                    <SPLIT distance="150" swimtime="00:02:26.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="250" reactiontime="+100" swimtime="00:01:28.16" resultid="6241" heatid="7599" lane="4" entrytime="00:01:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="130" reactiontime="+70" swimtime="00:03:29.24" resultid="6243" heatid="7765" lane="5" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.45" />
                    <SPLIT distance="100" swimtime="00:01:42.05" />
                    <SPLIT distance="150" swimtime="00:02:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="272" reactiontime="+100" swimtime="00:00:38.94" resultid="6244" heatid="7798" lane="6" entrytime="00:00:40.30" />
                <RESULT eventid="1559" points="180" reactiontime="+107" swimtime="00:06:56.63" resultid="7987" heatid="7974" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                    <SPLIT distance="100" swimtime="00:01:33.73" />
                    <SPLIT distance="150" swimtime="00:02:30.45" />
                    <SPLIT distance="200" swimtime="00:03:27.25" />
                    <SPLIT distance="250" swimtime="00:04:26.89" />
                    <SPLIT distance="300" swimtime="00:05:24.88" />
                    <SPLIT distance="350" swimtime="00:06:11.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Sergey" gender="M" lastname="Dirindyaev " nation="RUS" athleteid="6245">
              <RESULTS>
                <RESULT eventid="1075" points="324" reactiontime="+76" swimtime="00:00:29.55" resultid="6246" heatid="7362" lane="1" entrytime="00:00:30.30" />
                <RESULT eventid="1200" points="146" reactiontime="+64" swimtime="00:00:42.88" resultid="6247" heatid="7447" lane="5" entrytime="00:00:40.80" />
                <RESULT eventid="1268" points="332" reactiontime="+77" swimtime="00:01:04.85" resultid="6248" heatid="7510" lane="2" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="247" reactiontime="+74" swimtime="00:00:34.70" resultid="6249" heatid="7632" lane="6" entrytime="00:00:34.50" />
                <RESULT eventid="1662" points="263" swimtime="00:00:39.39" resultid="6250" heatid="7796" lane="5" entrytime="00:00:41.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Vadim" gender="M" lastname="Ezhkov " nation="RUS" athleteid="6251">
              <RESULTS>
                <RESULT eventid="1075" points="277" reactiontime="+72" swimtime="00:00:31.12" resultid="6252" heatid="7360" lane="1" entrytime="00:00:31.30" />
                <RESULT eventid="1234" points="289" reactiontime="+74" swimtime="00:03:02.46" resultid="6253" heatid="7478" lane="2" entrytime="00:03:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:25.02" />
                    <SPLIT distance="150" swimtime="00:02:13.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="313" reactiontime="+72" swimtime="00:01:21.85" resultid="6254" heatid="7604" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="269" reactiontime="+70" swimtime="00:00:33.73" resultid="6255" heatid="7631" lane="3" entrytime="00:00:34.50" />
                <RESULT comment="K-4" eventid="1662" status="DSQ" swimtime="00:00:36.14" resultid="8077" heatid="7804" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Viktor" gender="M" lastname="Liubavin " nation="RUS" athleteid="6257">
              <RESULTS>
                <RESULT eventid="1075" points="397" reactiontime="+84" swimtime="00:00:27.60" resultid="6258" heatid="7368" lane="3" entrytime="00:00:28.30" />
                <RESULT eventid="1268" points="412" reactiontime="+86" swimtime="00:01:00.37" resultid="6259" heatid="7520" lane="2" entrytime="00:01:00.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="354" reactiontime="+86" swimtime="00:01:18.54" resultid="6260" heatid="7605" lane="1" entrytime="00:01:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="362" reactiontime="+80" swimtime="00:02:19.41" resultid="6261" heatid="7701" lane="2" entrytime="00:02:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:09.48" />
                    <SPLIT distance="150" swimtime="00:01:45.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1594" points="266" reactiontime="+89" swimtime="00:01:15.34" resultid="6262" heatid="7746" lane="1" entrytime="00:01:13.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="365" reactiontime="+83" swimtime="00:00:35.31" resultid="6263" heatid="7804" lane="4" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Aleksandr" gender="M" lastname="Smirnov  " nation="RUS" athleteid="6264">
              <RESULTS>
                <RESULT eventid="1504" points="426" reactiontime="+98" swimtime="00:02:12.02" resultid="6266" heatid="7702" lane="4" entrytime="00:02:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:01:03.59" />
                    <SPLIT distance="150" swimtime="00:01:38.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" points="419" reactiontime="+97" swimtime="00:04:44.21" resultid="6267" heatid="8056" lane="2" entrytime="00:04:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:07.65" />
                    <SPLIT distance="150" swimtime="00:01:43.67" />
                    <SPLIT distance="200" swimtime="00:02:19.76" />
                    <SPLIT distance="250" swimtime="00:02:56.07" />
                    <SPLIT distance="300" swimtime="00:03:32.32" />
                    <SPLIT distance="350" swimtime="00:04:08.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="386" reactiontime="+99" swimtime="00:19:27.46" resultid="7158" heatid="7915" lane="3" entrytime="00:19:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:11.71" />
                    <SPLIT distance="150" swimtime="00:01:49.88" />
                    <SPLIT distance="200" swimtime="00:02:27.98" />
                    <SPLIT distance="250" swimtime="00:03:06.37" />
                    <SPLIT distance="300" swimtime="00:03:44.42" />
                    <SPLIT distance="350" swimtime="00:04:23.00" />
                    <SPLIT distance="400" swimtime="00:05:01.92" />
                    <SPLIT distance="450" swimtime="00:05:40.69" />
                    <SPLIT distance="500" swimtime="00:06:19.68" />
                    <SPLIT distance="550" swimtime="00:06:58.67" />
                    <SPLIT distance="600" swimtime="00:07:37.69" />
                    <SPLIT distance="650" swimtime="00:08:16.49" />
                    <SPLIT distance="700" swimtime="00:08:56.07" />
                    <SPLIT distance="750" swimtime="00:09:35.42" />
                    <SPLIT distance="800" swimtime="00:10:15.27" />
                    <SPLIT distance="850" swimtime="00:10:55.03" />
                    <SPLIT distance="900" swimtime="00:11:35.39" />
                    <SPLIT distance="950" swimtime="00:12:15.46" />
                    <SPLIT distance="1000" swimtime="00:12:55.13" />
                    <SPLIT distance="1050" swimtime="00:13:34.91" />
                    <SPLIT distance="1100" swimtime="00:14:15.09" />
                    <SPLIT distance="1150" swimtime="00:14:54.82" />
                    <SPLIT distance="1200" swimtime="00:15:34.17" />
                    <SPLIT distance="1250" swimtime="00:16:13.78" />
                    <SPLIT distance="1300" swimtime="00:16:53.22" />
                    <SPLIT distance="1350" swimtime="00:17:32.59" />
                    <SPLIT distance="1400" swimtime="00:18:12.06" />
                    <SPLIT distance="1450" swimtime="00:18:50.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="336" reactiontime="+69" swimtime="00:02:11.92" resultid="6281" heatid="7931" lane="5" entrytime="00:02:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:42.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6257" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="6251" number="2" />
                    <RELAYPOSITION athleteid="6230" number="3" />
                    <RELAYPOSITION athleteid="6245" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="344" reactiontime="+92" swimtime="00:01:55.22" resultid="6282" heatid="7712" lane="3" entrytime="00:02:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="100" swimtime="00:00:55.38" />
                    <SPLIT distance="150" swimtime="00:01:23.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6264" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="6257" number="2" reactiontime="+8" />
                    <RELAYPOSITION athleteid="6230" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="6217" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1521" points="302" reactiontime="+96" swimtime="00:02:18.87" resultid="6284" heatid="7707" lane="3" entrytime="00:02:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:07.93" />
                    <SPLIT distance="150" swimtime="00:01:43.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6200" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="6185" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="6205" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="6195" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1370" points="302" reactiontime="+56" swimtime="00:02:33.05" resultid="6280" heatid="7572" lane="4" entrytime="00:02:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:22.31" />
                    <SPLIT distance="150" swimtime="00:01:58.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6200" number="1" reactiontime="+56" />
                    <RELAYPOSITION athleteid="6185" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="6205" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="6195" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1126" points="272" reactiontime="+98" swimtime="00:02:04.54" resultid="6278" heatid="7409" lane="2" entrytime="00:02:14.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6200" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="6238" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="6245" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="6185" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="6285" heatid="7817" lane="6" entrytime="00:02:25.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6200" number="1" />
                    <RELAYPOSITION athleteid="6251" number="2" />
                    <RELAYPOSITION athleteid="6230" number="3" />
                    <RELAYPOSITION athleteid="6185" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="6279" heatid="7410" lane="3" entrytime="00:02:01.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6264" number="1" />
                    <RELAYPOSITION athleteid="6257" number="2" />
                    <RELAYPOSITION athleteid="6205" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="6286" heatid="7817" lane="4" entrytime="00:02:18.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6205" number="1" />
                    <RELAYPOSITION athleteid="6257" number="2" />
                    <RELAYPOSITION athleteid="6264" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Kaliningrad" nation="RUS">
          <ATHLETES>
            <ATHLETE birthdate="1970-01-01" firstname="Svetlana" gender="F" lastname="Smirnova  " nation="RUS" athleteid="6270">
              <RESULTS>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="6271" heatid="7779" lane="6" entrytime="00:00:52.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Moskow" nation="RUS">
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Aleksandr" gender="M" lastname="Zelenov " nation="RUS" athleteid="6273">
              <RESULTS>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="6275" heatid="7502" lane="5" entrytime="00:01:37.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="6276" heatid="7688" lane="4" entrytime="00:03:37.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Swimmers Stowarzyszenie Pływackie" nation="POL" region="MAZ" shortname="Swimmers Stowarzyszenie Pływac">
          <CONTACT city="WARSZAWA" email="INFO@SWIMMERSTEAM.PL" name="GOŁĘBIOWSKI REMIGIUSZ" phone="601333782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1976-07-07" firstname="Remigiusz" gender="M" lastname="Gołębiowski" nation="POL" athleteid="6291">
              <RESULTS>
                <RESULT eventid="1075" points="445" reactiontime="+76" swimtime="00:00:26.58" resultid="6292" heatid="7373" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="6294" heatid="7521" lane="4" entrytime="00:00:59.00" />
                <RESULT eventid="1436" points="460" reactiontime="+79" swimtime="00:00:28.24" resultid="6295" heatid="7644" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="6296" heatid="7704" lane="1" entrytime="00:02:10.00" />
                <RESULT eventid="1594" status="DNS" swimtime="00:00:00.00" resultid="6297" heatid="7749" lane="2" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-14" firstname="Hubert" gender="M" lastname="Lis" nation="POL" athleteid="6299">
              <RESULTS>
                <RESULT eventid="1075" points="406" reactiontime="+85" swimtime="00:00:27.41" resultid="6300" heatid="7373" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1200" points="349" reactiontime="+65" swimtime="00:00:32.10" resultid="6301" heatid="7457" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1436" points="388" reactiontime="+88" swimtime="00:00:29.88" resultid="6302" heatid="7642" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1662" points="335" reactiontime="+83" swimtime="00:00:36.34" resultid="6303" heatid="7810" lane="3" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-10-21" firstname="Piotr" gender="M" lastname="Macioszek" nation="POL" athleteid="6304">
              <RESULTS>
                <RESULT eventid="1268" points="144" reactiontime="+98" swimtime="00:01:25.72" resultid="6305" heatid="7507" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="125" reactiontime="+93" swimtime="00:01:41.36" resultid="6306" heatid="7540" lane="3" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="6307" heatid="7626" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="6308" heatid="7691" lane="2" entrytime="00:02:55.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="6309" heatid="7793" lane="6" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-12" firstname="Jan" gender="M" lastname="Rekowski" nation="POL" athleteid="6310">
              <RESULTS>
                <RESULT eventid="1075" points="499" reactiontime="+72" swimtime="00:00:25.59" resultid="6311" heatid="7378" lane="3" entrytime="00:00:25.60" />
                <RESULT eventid="1268" points="481" reactiontime="+80" swimtime="00:00:57.33" resultid="6312" heatid="7522" lane="2" entrytime="00:00:58.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="363" swimtime="00:01:11.13" resultid="6313" heatid="7554" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="412" reactiontime="+87" swimtime="00:00:29.28" resultid="6314" heatid="7641" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1470" status="DNS" swimtime="00:00:00.00" resultid="6315" heatid="7669" lane="6" entrytime="00:01:14.00" />
                <RESULT eventid="1662" points="333" swimtime="00:00:36.42" resultid="6316" heatid="7802" lane="5" entrytime="00:00:37.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-03" firstname="Bolesław" gender="M" lastname="Porolniczak" nation="POL" athleteid="6317">
              <RESULTS>
                <RESULT eventid="1075" points="425" reactiontime="+87" swimtime="00:00:26.98" resultid="6318" heatid="7374" lane="3" entrytime="00:00:26.90" />
                <RESULT eventid="1268" points="384" reactiontime="+90" swimtime="00:01:01.78" resultid="6319" heatid="7518" lane="1" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="350" reactiontime="+95" swimtime="00:00:30.91" resultid="6320" heatid="7640" lane="3" entrytime="00:00:29.78" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-05-27" firstname="Mariusz" gender="M" lastname="Bartczak" nation="POL" athleteid="6321">
              <RESULTS>
                <RESULT eventid="1075" points="234" reactiontime="+115" swimtime="00:00:32.90" resultid="6322" heatid="7353" lane="3" entrytime="00:00:34.50" />
                <RESULT eventid="1268" points="204" reactiontime="+98" swimtime="00:01:16.32" resultid="6323" heatid="7506" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="187" reactiontime="+112" swimtime="00:02:53.70" resultid="6324" heatid="7694" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                    <SPLIT distance="150" swimtime="00:02:08.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-07" firstname="Paweł" gender="M" lastname="Witkowski" nation="POL" athleteid="6326">
              <RESULTS>
                <RESULT eventid="1075" points="230" reactiontime="+102" swimtime="00:00:33.13" resultid="6327" heatid="7356" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1268" points="211" reactiontime="+92" swimtime="00:01:15.44" resultid="6328" heatid="7509" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="213" swimtime="00:01:33.08" resultid="6329" heatid="7598" lane="5" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="237" reactiontime="+96" swimtime="00:00:40.77" resultid="6330" heatid="7796" lane="4" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-12-11" firstname="Mikołaj" gender="M" lastname="Tusiński" nation="POL" athleteid="6331">
              <RESULTS>
                <RESULT eventid="1075" points="420" reactiontime="+86" swimtime="00:00:27.10" resultid="6332" heatid="7374" lane="4" entrytime="00:00:26.90" />
                <RESULT eventid="1200" points="277" reactiontime="+62" swimtime="00:00:34.67" resultid="6333" heatid="7456" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1268" points="436" reactiontime="+86" swimtime="00:00:59.25" resultid="6334" heatid="7521" lane="6" entrytime="00:00:59.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="410" reactiontime="+79" swimtime="00:00:29.33" resultid="6335" heatid="7641" lane="6" entrytime="00:00:29.50" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="6336" heatid="7808" lane="5" entrytime="00:00:34.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-12-20" firstname="Arkadiusz" gender="M" lastname="Aptewicz" nation="POL" athleteid="6337">
              <RESULTS>
                <RESULT eventid="1109" points="549" reactiontime="+72" swimtime="00:02:14.39" resultid="6338" heatid="7407" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                    <SPLIT distance="100" swimtime="00:01:04.55" />
                    <SPLIT distance="150" swimtime="00:01:42.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="591" reactiontime="+68" swimtime="00:02:23.75" resultid="6339" heatid="7485" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="599" reactiontime="+78" swimtime="00:01:00.21" resultid="6340" heatid="7560" lane="4" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="606" reactiontime="+74" swimtime="00:01:05.71" resultid="6341" heatid="7611" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="6342" heatid="7706" lane="5" entrytime="00:01:59.50" />
                <RESULT eventid="1594" points="533" swimtime="00:00:59.78" resultid="6343" heatid="7752" lane="5" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="595" reactiontime="+72" swimtime="00:00:30.02" resultid="6344" heatid="7813" lane="2" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brożyna" nation="POL" athleteid="6345">
              <RESULTS>
                <RESULT eventid="1109" points="266" reactiontime="+88" swimtime="00:02:51.13" resultid="6346" heatid="7401" lane="1" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:16.78" />
                    <SPLIT distance="150" swimtime="00:02:09.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="288" reactiontime="+66" swimtime="00:00:34.21" resultid="6347" heatid="7452" lane="3" entrytime="00:00:33.90" />
                <RESULT eventid="1470" points="277" reactiontime="+75" swimtime="00:01:15.05" resultid="6348" heatid="7668" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" status="DNS" swimtime="00:00:00.00" resultid="6349" heatid="7768" lane="3" entrytime="00:02:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-07" firstname="Mariusz" gender="M" lastname="Iller" nation="POL" athleteid="6350">
              <RESULTS>
                <RESULT eventid="1075" points="94" reactiontime="+111" swimtime="00:00:44.64" resultid="6351" heatid="7348" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="6352" heatid="7791" lane="5" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-05-13" firstname="Michał" gender="M" lastname="Witkowski" nation="POL" athleteid="6353">
              <RESULTS>
                <RESULT eventid="1075" points="440" reactiontime="+70" swimtime="00:00:26.68" resultid="6354" heatid="7377" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="6355" heatid="7455" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1268" points="443" swimtime="00:00:58.95" resultid="6356" heatid="7523" lane="5" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="474" reactiontime="+70" swimtime="00:00:27.95" resultid="6357" heatid="7644" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1594" points="418" reactiontime="+69" swimtime="00:01:04.81" resultid="6358" heatid="7750" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-21" firstname="Anna" gender="F" lastname="Jabłońska" nation="POL" athleteid="6359">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="6360" heatid="7339" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1183" points="233" reactiontime="+90" swimtime="00:00:41.72" resultid="6361" heatid="7438" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1285" points="193" swimtime="00:01:39.89" resultid="6362" heatid="7532" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="6363" heatid="7653" lane="6" entrytime="00:01:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-29" firstname="Urszula" gender="F" lastname="Jakubowska-Cłapińska" nation="POL" athleteid="6364">
              <RESULTS>
                <RESULT eventid="1058" points="287" reactiontime="+86" swimtime="00:00:35.21" resultid="6365" heatid="7339" lane="6" entrytime="00:00:34.80" />
                <RESULT eventid="1092" points="244" reactiontime="+90" swimtime="00:03:19.24" resultid="6366" heatid="7386" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                    <SPLIT distance="100" swimtime="00:01:31.42" />
                    <SPLIT distance="150" swimtime="00:02:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" status="DNS" swimtime="00:00:00.00" resultid="6367" heatid="7436" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1285" points="279" reactiontime="+85" swimtime="00:01:28.26" resultid="6368" heatid="7531" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="6369" heatid="7655" lane="1" entrytime="00:01:23.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-12" firstname="Katarzyna" gender="F" lastname="Blajer" nation="POL" athleteid="6370">
              <RESULTS>
                <RESULT eventid="1058" points="176" swimtime="00:00:41.48" resultid="6371" heatid="7335" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="1251" points="136" reactiontime="+106" swimtime="00:01:39.12" resultid="6372" heatid="7490" lane="2" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="152" reactiontime="+87" swimtime="00:01:57.30" resultid="6373" heatid="7585" lane="2" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="174" reactiontime="+97" swimtime="00:00:51.55" resultid="6374" heatid="7781" lane="3" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-11" firstname="Ewa" gender="F" lastname="Gałązka" nation="POL" athleteid="6375">
              <RESULTS>
                <RESULT eventid="1058" points="201" reactiontime="+115" swimtime="00:00:39.65" resultid="6376" heatid="7334" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="1251" points="136" reactiontime="+127" swimtime="00:01:38.99" resultid="6377" heatid="7488" lane="3" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-18" firstname="Małgorzata" gender="F" lastname="Wietrzykowska" nation="POL" athleteid="6378">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="6379" heatid="7333" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1183" points="88" reactiontime="+103" swimtime="00:00:57.62" resultid="6380" heatid="7433" lane="6" entrytime="00:00:55.00" />
                <RESULT eventid="1645" points="149" reactiontime="+123" swimtime="00:00:54.27" resultid="6381" heatid="7777" lane="1" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-01" firstname="Katarzyna" gender="F" lastname="Koba" nation="POL" athleteid="6382">
              <RESULTS>
                <RESULT eventid="1058" points="400" swimtime="00:00:31.53" resultid="6383" heatid="7342" lane="5" entrytime="00:00:31.49" />
                <RESULT eventid="1251" points="353" reactiontime="+90" swimtime="00:01:12.14" resultid="6384" heatid="7495" lane="1" entrytime="00:01:12.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="311" reactiontime="+92" swimtime="00:02:43.97" resultid="6385" heatid="7683" lane="1" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                    <SPLIT distance="150" swimtime="00:02:00.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-07-31" firstname="Katarzyna" gender="F" lastname="Herczyńska" nation="POL" athleteid="6386">
              <RESULTS>
                <RESULT eventid="1285" points="286" reactiontime="+91" swimtime="00:01:27.54" resultid="6387" heatid="7533" lane="4" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="263" reactiontime="+91" swimtime="00:00:38.03" resultid="6388" heatid="7618" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1377" points="403" reactiontime="+67" swimtime="00:02:04.23" resultid="6395" heatid="7929" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:38.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6345" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="6299" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="6291" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="6310" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1528" points="466" reactiontime="+85" swimtime="00:01:44.17" resultid="6396" heatid="7709" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.55" />
                    <SPLIT distance="100" swimtime="00:00:51.70" />
                    <SPLIT distance="150" swimtime="00:01:17.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6317" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="6331" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="6291" number="3" reactiontime="+8" />
                    <RELAYPOSITION athleteid="6310" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT comment="K-15" eventid="1377" reactiontime="+61" status="DSQ" swimtime="00:02:26.28" resultid="6397" heatid="7928" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:20.01" />
                    <SPLIT distance="150" swimtime="00:01:59.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6321" number="1" reactiontime="+61" status="DSQ" />
                    <RELAYPOSITION athleteid="6326" number="2" reactiontime="+44" status="DSQ" />
                    <RELAYPOSITION athleteid="6331" number="3" reactiontime="+66" status="DSQ" />
                    <RELAYPOSITION athleteid="6317" number="4" reactiontime="+21" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="6398" heatid="7710" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6350" number="1" />
                    <RELAYPOSITION athleteid="6304" number="2" />
                    <RELAYPOSITION athleteid="6321" number="3" />
                    <RELAYPOSITION athleteid="6326" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1370" points="248" reactiontime="+70" swimtime="00:02:43.42" resultid="6393" heatid="7572" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                    <SPLIT distance="100" swimtime="00:01:34.65" />
                    <SPLIT distance="150" swimtime="00:02:11.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6359" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="6364" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="6386" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="6382" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1521" points="299" reactiontime="+91" swimtime="00:02:19.31" resultid="6394" heatid="7707" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:11.97" />
                    <SPLIT distance="150" swimtime="00:01:47.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6364" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="6359" number="2" reactiontime="+87" />
                    <RELAYPOSITION athleteid="6386" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="6382" number="4" reactiontime="+86" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1126" points="321" swimtime="00:01:57.91" resultid="6389" heatid="7408" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:00:57.53" />
                    <SPLIT distance="150" swimtime="00:01:32.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6310" number="1" />
                    <RELAYPOSITION athleteid="6359" number="2" />
                    <RELAYPOSITION athleteid="6331" number="3" />
                    <RELAYPOSITION athleteid="6382" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" points="261" reactiontime="+72" swimtime="00:02:23.61" resultid="6390" heatid="7814" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:01:47.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6364" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="6326" number="2" reactiontime="+79" />
                    <RELAYPOSITION athleteid="6386" number="3" reactiontime="+12" />
                    <RELAYPOSITION athleteid="6331" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1126" points="217" reactiontime="+104" swimtime="00:02:14.31" resultid="6391" heatid="7408" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.28" />
                    <SPLIT distance="150" swimtime="00:01:47.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6364" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="6317" number="2" reactiontime="+3" />
                    <RELAYPOSITION athleteid="6370" number="3" />
                    <RELAYPOSITION athleteid="6291" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1679" points="294" reactiontime="+67" swimtime="00:02:18.03" resultid="6392" heatid="7815" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:46.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6345" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="6310" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="6386" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="6382" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1679" points="211" reactiontime="+68" swimtime="00:02:34.08" resultid="6399" heatid="7816" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:01:21.90" />
                    <SPLIT distance="150" swimtime="00:01:57.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6359" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="6299" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="6310" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="6378" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="KPS Nereus Zilina" nation="SVK">
          <ATHLETES>
            <ATHLETE birthdate="1989-01-01" firstname="Lukas" gender="M" lastname="Smiesko " nation="POL" athleteid="6426">
              <RESULTS>
                <RESULT eventid="1200" points="485" reactiontime="+66" swimtime="00:00:28.77" resultid="6427" heatid="7459" lane="6" entrytime="00:00:29.23" />
                <RESULT eventid="1302" points="586" reactiontime="+76" swimtime="00:01:00.64" resultid="6428" heatid="7560" lane="1" entrytime="00:01:01.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="564" reactiontime="+76" swimtime="00:00:26.38" resultid="6429" heatid="7647" lane="6" entrytime="00:00:26.37" />
                <RESULT eventid="1470" points="468" reactiontime="+61" swimtime="00:01:03.00" resultid="6430" heatid="7674" lane="2" entrytime="00:01:00.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Rastislav" gender="M" lastname="Pavlik " nation="SVK" athleteid="6431">
              <RESULTS>
                <RESULT eventid="1075" points="443" reactiontime="+83" swimtime="00:00:26.62" resultid="6432" heatid="7374" lane="2" entrytime="00:00:26.96" />
                <RESULT eventid="1200" points="397" reactiontime="+73" swimtime="00:00:30.74" resultid="6433" heatid="7456" lane="4" entrytime="00:00:30.89" />
                <RESULT eventid="1302" points="455" reactiontime="+82" swimtime="00:01:05.98" resultid="6434" heatid="7557" lane="4" entrytime="00:01:06.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="409" swimtime="00:01:05.92" resultid="6435" heatid="7672" lane="2" entrytime="00:01:05.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1662" points="429" reactiontime="+88" swimtime="00:00:33.47" resultid="6436" heatid="7809" lane="6" entrytime="00:00:34.11" />
                <RESULT eventid="1710" points="313" reactiontime="+72" swimtime="00:05:13.10" resultid="6437" heatid="8052" lane="3" entrytime="00:05:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:01:51.13" />
                    <SPLIT distance="200" swimtime="00:02:30.78" />
                    <SPLIT distance="250" swimtime="00:03:11.83" />
                    <SPLIT distance="300" swimtime="00:03:52.71" />
                    <SPLIT distance="350" swimtime="00:04:34.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="WOPR Kędzierzyn-Koźle" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1958-01-01" firstname="RYSZARD" gender="M" lastname="TATARCZUK " nation="POL" athleteid="6441">
              <RESULTS>
                <RESULT eventid="1165" points="171" swimtime="00:25:30.11" resultid="6442" heatid="7909" lane="5" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:01:27.91" />
                    <SPLIT distance="150" swimtime="00:02:15.26" />
                    <SPLIT distance="200" swimtime="00:03:02.73" />
                    <SPLIT distance="250" swimtime="00:03:51.62" />
                    <SPLIT distance="300" swimtime="00:04:41.14" />
                    <SPLIT distance="350" swimtime="00:05:30.30" />
                    <SPLIT distance="400" swimtime="00:06:20.08" />
                    <SPLIT distance="450" swimtime="00:07:10.33" />
                    <SPLIT distance="500" swimtime="00:08:00.45" />
                    <SPLIT distance="550" swimtime="00:08:50.68" />
                    <SPLIT distance="600" swimtime="00:09:43.04" />
                    <SPLIT distance="650" swimtime="00:10:34.24" />
                    <SPLIT distance="700" swimtime="00:11:26.74" />
                    <SPLIT distance="750" swimtime="00:12:18.48" />
                    <SPLIT distance="800" swimtime="00:13:10.60" />
                    <SPLIT distance="850" swimtime="00:14:03.43" />
                    <SPLIT distance="900" swimtime="00:14:55.81" />
                    <SPLIT distance="950" swimtime="00:15:48.21" />
                    <SPLIT distance="1000" swimtime="00:16:41.00" />
                    <SPLIT distance="1050" swimtime="00:17:33.21" />
                    <SPLIT distance="1100" swimtime="00:18:25.62" />
                    <SPLIT distance="1150" swimtime="00:19:18.15" />
                    <SPLIT distance="1200" swimtime="00:20:11.85" />
                    <SPLIT distance="1250" swimtime="00:21:05.87" />
                    <SPLIT distance="1300" swimtime="00:21:58.83" />
                    <SPLIT distance="1350" swimtime="00:22:52.61" />
                    <SPLIT distance="1400" swimtime="00:23:46.83" />
                    <SPLIT distance="1450" swimtime="00:24:39.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="245" reactiontime="+95" swimtime="00:00:32.43" resultid="6443" heatid="7352" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" name="KU AZS UAM Poznań" nation="POL" region="PO">
          <CONTACT city="Poznań" email="kukowalazs@gmail.com" name="Kowalik" phone="603965223" state="WLKP" street="Zagajnikowa 9" zip="61-602" />
          <ATHLETES>
            <ATHLETE birthdate="1977-03-14" firstname="Jarosław" gender="M" lastname="Bystry" nation="POL" athleteid="7126">
              <RESULTS>
                <RESULT eventid="1075" points="368" swimtime="00:00:28.32" resultid="7127" heatid="7369" lane="5" entrytime="00:00:28.20" />
                <RESULT eventid="1268" points="357" reactiontime="+86" swimtime="00:01:03.31" resultid="7128" heatid="7518" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="278" reactiontime="+84" swimtime="00:01:17.74" resultid="7129" heatid="7550" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="7130" heatid="7637" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="7131" heatid="7701" lane="1" entrytime="00:02:20.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="7132" heatid="7801" lane="3" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="Stadnik" nation="POL" license="103315100003" athleteid="7133">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1058" points="618" reactiontime="+61" swimtime="00:00:27.29" resultid="7134" heatid="7344" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="1183" points="482" reactiontime="+81" swimtime="00:00:32.77" resultid="7135" heatid="7441" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1251" points="638" reactiontime="+80" swimtime="00:00:59.25" resultid="7136" heatid="7498" lane="3" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="482" reactiontime="+70" swimtime="00:01:10.43" resultid="7137" heatid="7658" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="531" swimtime="00:02:17.25" resultid="7138" heatid="7685" lane="5" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:01:07.08" />
                    <SPLIT distance="150" swimtime="00:01:42.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="412" reactiontime="+77" swimtime="00:02:41.22" resultid="7139" heatid="7761" lane="2" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:16.93" />
                    <SPLIT distance="150" swimtime="00:02:00.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="495" reactiontime="+73" swimtime="00:00:36.39" resultid="7140" heatid="7786" lane="4" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="Sterczyński" nation="POL" license="103315200002" athleteid="7141">
              <RESULTS>
                <RESULT eventid="1109" points="489" reactiontime="+74" swimtime="00:02:19.68" resultid="7142" heatid="7406" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="100" swimtime="00:01:04.71" />
                    <SPLIT distance="150" swimtime="00:01:45.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="426" reactiontime="+65" swimtime="00:00:30.03" resultid="7143" heatid="7458" lane="5" entrytime="00:00:29.60" />
                <RESULT eventid="1302" points="508" swimtime="00:01:03.60" resultid="7144" heatid="7559" lane="5" entrytime="00:01:03.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="455" reactiontime="+69" swimtime="00:01:03.62" resultid="7145" heatid="7673" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="451" reactiontime="+77" swimtime="00:05:06.88" resultid="7146" heatid="7980" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="100" swimtime="00:01:04.57" />
                    <SPLIT distance="150" swimtime="00:01:44.31" />
                    <SPLIT distance="200" swimtime="00:02:24.00" />
                    <SPLIT distance="250" swimtime="00:03:07.58" />
                    <SPLIT distance="300" swimtime="00:03:52.25" />
                    <SPLIT distance="350" swimtime="00:04:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="440" reactiontime="+69" swimtime="00:02:19.45" resultid="7147" heatid="7774" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:06.17" />
                    <SPLIT distance="150" swimtime="00:01:42.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZSWSB" name="AZS WSB Dąbrowa Górnicza" nation="POL" region="KA">
          <CONTACT city="Dąbrowa Górnicza" email="kacperkapron@wp.pl" name="Kaproń Kacper" phone="791512012" state="ŚLĄSK" zip="41-300" />
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="7149">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="7150" heatid="7379" lane="3" entrytime="00:00:25.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="7151" heatid="7402" lane="1" entrytime="00:02:40.00" />
                <RESULT eventid="1200" status="DNS" swimtime="00:00:00.00" resultid="7152" heatid="7455" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="7153" heatid="7481" lane="4" entrytime="00:02:55.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="7154" heatid="7606" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1504" status="DNS" swimtime="00:00:00.00" resultid="7155" heatid="7703" lane="4" entrytime="00:02:10.00" />
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="7157" heatid="8054" lane="3" entrytime="00:04:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" name="AZS AWF Katowice" nation="POL" region="SLA">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1931-04-27" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" athleteid="7177">
              <RESULTS>
                <RESULT eventid="1165" points="30" reactiontime="+93" swimtime="00:45:14.39" resultid="7178" heatid="7907" lane="4" entrytime="00:44:50.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.81" />
                    <SPLIT distance="100" swimtime="00:02:46.61" />
                    <SPLIT distance="150" swimtime="00:04:16.25" />
                    <SPLIT distance="200" swimtime="00:05:40.67" />
                    <SPLIT distance="250" swimtime="00:07:09.98" />
                    <SPLIT distance="300" swimtime="00:08:36.79" />
                    <SPLIT distance="350" swimtime="00:10:09.06" />
                    <SPLIT distance="400" swimtime="00:11:37.39" />
                    <SPLIT distance="450" swimtime="00:13:12.41" />
                    <SPLIT distance="500" swimtime="00:14:41.64" />
                    <SPLIT distance="550" swimtime="00:16:15.95" />
                    <SPLIT distance="600" swimtime="00:17:44.55" />
                    <SPLIT distance="650" swimtime="00:19:18.03" />
                    <SPLIT distance="700" swimtime="00:20:48.83" />
                    <SPLIT distance="750" swimtime="00:22:24.74" />
                    <SPLIT distance="800" swimtime="00:23:52.50" />
                    <SPLIT distance="850" swimtime="00:25:30.72" />
                    <SPLIT distance="900" swimtime="00:26:58.43" />
                    <SPLIT distance="950" swimtime="00:28:33.01" />
                    <SPLIT distance="1000" swimtime="00:30:01.93" />
                    <SPLIT distance="1050" swimtime="00:31:34.93" />
                    <SPLIT distance="1100" swimtime="00:33:07.02" />
                    <SPLIT distance="1150" swimtime="00:34:41.05" />
                    <SPLIT distance="1200" swimtime="00:36:16.00" />
                    <SPLIT distance="1250" swimtime="00:37:49.03" />
                    <SPLIT distance="1300" swimtime="00:39:19.97" />
                    <SPLIT distance="1350" swimtime="00:40:52.90" />
                    <SPLIT distance="1400" swimtime="00:42:25.27" />
                    <SPLIT distance="1450" swimtime="00:43:56.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="46" reactiontime="+103" swimtime="00:05:34.62" resultid="7179" heatid="7471" lane="2" entrytime="00:05:23.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.74" />
                    <SPLIT distance="100" swimtime="00:02:43.93" />
                    <SPLIT distance="150" swimtime="00:04:10.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="30" reactiontime="+96" swimtime="00:05:19.06" resultid="7180" heatid="7687" lane="2" entrytime="00:05:03.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.28" />
                    <SPLIT distance="100" swimtime="00:02:35.13" />
                    <SPLIT distance="150" swimtime="00:04:00.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1710" reactiontime="+65" status="DSQ" swimtime="00:10:57.36" resultid="7181" heatid="8044" lane="2" entrytime="00:10:46.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.50" />
                    <SPLIT distance="100" swimtime="00:02:34.79" />
                    <SPLIT distance="150" swimtime="00:03:58.96" />
                    <SPLIT distance="200" swimtime="00:05:22.15" />
                    <SPLIT distance="250" swimtime="00:06:46.67" />
                    <SPLIT distance="300" swimtime="00:08:10.07" />
                    <SPLIT distance="350" swimtime="00:09:33.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-08-05" firstname="Tomasz" gender="M" lastname="Polewka" nation="POL" license="100611200220" athleteid="7182">
              <RESULTS>
                <RESULT eventid="1200" points="790" reactiontime="+51" swimtime="00:00:24.45" resultid="7183" heatid="7460" lane="3" entrytime="00:00:23.62" />
                <RESULT eventid="1268" points="648" reactiontime="+76" swimtime="00:00:51.92" resultid="7184" heatid="7525" lane="4" entrytime="00:00:50.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="622" reactiontime="+79" swimtime="00:00:25.53" resultid="7185" heatid="7622" lane="4" />
                <RESULT eventid="1470" points="723" reactiontime="+62" swimtime="00:00:54.51" resultid="7186" heatid="7674" lane="3" entrytime="00:00:52.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.96" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="3 start w bloku." eventid="1504" points="600" reactiontime="+80" status="EXH" swimtime="00:01:57.77" resultid="7187" heatid="7686" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                    <SPLIT distance="100" swimtime="00:00:57.68" />
                    <SPLIT distance="150" swimtime="00:01:28.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-05-08" firstname="Marlena" gender="F" lastname="Dudek" nation="POL" license="100611100198" athleteid="7188">
              <RESULTS>
                <RESULT eventid="1058" points="533" swimtime="00:00:28.66" resultid="7189" heatid="7331" lane="5" />
                <RESULT eventid="1217" points="600" reactiontime="+77" swimtime="00:02:39.50" resultid="7190" heatid="7469" lane="3" entrytime="00:02:30.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:16.42" />
                    <SPLIT distance="150" swimtime="00:01:58.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="546" reactiontime="+83" swimtime="00:01:10.63" resultid="7191" heatid="7526" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-05-27" firstname="Wojciech" gender="M" lastname="Głyk" nation="POL" license="100611200202" athleteid="7192">
              <RESULTS>
                <RESULT eventid="1165" points="747" reactiontime="+85" swimtime="00:15:36.79" resultid="7193" heatid="7917" lane="3" entrytime="00:15:27.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="100" swimtime="00:01:01.27" />
                    <SPLIT distance="150" swimtime="00:01:33.10" />
                    <SPLIT distance="200" swimtime="00:02:04.78" />
                    <SPLIT distance="250" swimtime="00:02:36.63" />
                    <SPLIT distance="300" swimtime="00:03:08.38" />
                    <SPLIT distance="350" swimtime="00:03:39.70" />
                    <SPLIT distance="400" swimtime="00:04:11.15" />
                    <SPLIT distance="450" swimtime="00:04:42.65" />
                    <SPLIT distance="500" swimtime="00:05:13.72" />
                    <SPLIT distance="550" swimtime="00:05:44.86" />
                    <SPLIT distance="600" swimtime="00:06:15.87" />
                    <SPLIT distance="650" swimtime="00:06:47.03" />
                    <SPLIT distance="700" swimtime="00:07:18.16" />
                    <SPLIT distance="750" swimtime="00:07:49.29" />
                    <SPLIT distance="800" swimtime="00:08:20.48" />
                    <SPLIT distance="850" swimtime="00:08:51.91" />
                    <SPLIT distance="900" swimtime="00:09:23.31" />
                    <SPLIT distance="950" swimtime="00:09:54.75" />
                    <SPLIT distance="1000" swimtime="00:10:25.90" />
                    <SPLIT distance="1050" swimtime="00:10:57.29" />
                    <SPLIT distance="1100" swimtime="00:11:28.53" />
                    <SPLIT distance="1150" swimtime="00:11:59.85" />
                    <SPLIT distance="1200" swimtime="00:12:31.35" />
                    <SPLIT distance="1250" swimtime="00:13:02.70" />
                    <SPLIT distance="1300" swimtime="00:13:33.98" />
                    <SPLIT distance="1350" swimtime="00:14:05.05" />
                    <SPLIT distance="1400" swimtime="00:14:36.64" />
                    <SPLIT distance="1450" swimtime="00:15:07.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="689" reactiontime="+84" swimtime="00:01:52.49" resultid="7194" heatid="7706" lane="3" entrytime="00:01:51.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.00" />
                    <SPLIT distance="100" swimtime="00:00:55.74" />
                    <SPLIT distance="150" swimtime="00:01:24.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="7195" heatid="8058" lane="3" entrytime="00:03:54.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-05-19" firstname="Łukasz" gender="M" lastname="Chmiel" nation="POL" license="100611200212" athleteid="7196">
              <RESULTS>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1075" reactiontime="+48" status="DSQ" swimtime="00:00:23.71" resultid="7197" heatid="7381" lane="2" entrytime="00:00:23.71" />
                <RESULT eventid="1109" points="601" reactiontime="+85" swimtime="00:02:10.38" resultid="7198" heatid="7407" lane="3" entrytime="00:02:05.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                    <SPLIT distance="100" swimtime="00:01:00.86" />
                    <SPLIT distance="150" swimtime="00:01:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="574" reactiontime="+65" swimtime="00:00:27.20" resultid="7199" heatid="7460" lane="2" entrytime="00:00:26.02" />
                <RESULT eventid="1302" points="625" reactiontime="+77" swimtime="00:00:59.34" resultid="7200" heatid="7560" lane="3" entrytime="00:00:53.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="539" reactiontime="+84" swimtime="00:01:08.33" resultid="7201" heatid="7593" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" status="DNS" swimtime="00:00:00.00" resultid="7202" heatid="7647" lane="3" entrytime="00:00:24.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="7203" heatid="7788" lane="4" />
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="7204" heatid="8044" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-06-20" firstname="Mateusz" gender="M" lastname="Szewczyk" nation="POL" athleteid="7205">
              <RESULTS>
                <RESULT eventid="1075" points="567" reactiontime="+63" swimtime="00:00:24.52" resultid="7206" heatid="7380" lane="3" entrytime="00:00:24.50" />
                <RESULT eventid="1200" points="511" reactiontime="+53" swimtime="00:00:28.28" resultid="7208" heatid="7459" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1302" points="506" reactiontime="+62" swimtime="00:01:03.66" resultid="7209" heatid="7558" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="512" reactiontime="+50" swimtime="00:01:01.14" resultid="7210" heatid="7674" lane="1" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1559" points="402" reactiontime="+69" swimtime="00:05:19.08" resultid="7211" heatid="7983" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="100" swimtime="00:01:05.53" />
                    <SPLIT distance="150" swimtime="00:01:46.22" />
                    <SPLIT distance="200" swimtime="00:02:25.70" />
                    <SPLIT distance="250" swimtime="00:03:13.55" />
                    <SPLIT distance="300" swimtime="00:04:02.30" />
                    <SPLIT distance="350" swimtime="00:04:41.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1628" points="442" reactiontime="+54" swimtime="00:02:19.21" resultid="7212" heatid="7774" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:06.20" />
                    <SPLIT distance="150" swimtime="00:01:43.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="7213" heatid="8057" lane="3" entrytime="00:04:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-27" firstname="Aleksandra" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="7214">
              <RESULTS>
                <RESULT eventid="1058" points="541" reactiontime="+69" swimtime="00:00:28.53" resultid="7215" heatid="7344" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1183" points="565" reactiontime="+69" swimtime="00:00:31.08" resultid="7216" heatid="7441" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1251" points="540" reactiontime="+70" swimtime="00:01:02.63" resultid="7217" heatid="7497" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="535" reactiontime="+67" swimtime="00:01:08.03" resultid="7218" heatid="7658" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1487" points="450" reactiontime="+75" swimtime="00:02:25.02" resultid="7219" heatid="7685" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1611" points="523" reactiontime="+71" swimtime="00:02:28.92" resultid="7220" heatid="7761" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:12.95" />
                    <SPLIT distance="150" swimtime="00:01:52.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-01" firstname="Robert" gender="M" lastname="Wilk" nation="POL" license="100611200111" athleteid="7221">
              <RESULTS>
                <RESULT eventid="1075" points="609" reactiontime="+72" swimtime="00:00:23.94" resultid="7222" heatid="7381" lane="3" entrytime="00:00:22.89" />
                <RESULT eventid="1268" points="608" swimtime="00:00:53.04" resultid="7223" heatid="7525" lane="5" entrytime="00:00:52.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="592" reactiontime="+71" swimtime="00:00:25.96" resultid="7224" heatid="7647" lane="2" entrytime="00:00:24.53" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-09-13" firstname="Tomasz" gender="M" lastname="Czermak" nation="POL" license="100611200197" athleteid="7225">
              <RESULTS>
                <RESULT eventid="1075" points="484" reactiontime="+75" swimtime="00:00:25.85" resultid="7226" heatid="7380" lane="1" entrytime="00:00:24.90" />
                <RESULT eventid="1109" points="520" reactiontime="+78" swimtime="00:02:16.86" resultid="7227" heatid="7407" lane="1" entrytime="00:02:16.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:06.30" />
                    <SPLIT distance="150" swimtime="00:01:43.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="555" reactiontime="+83" swimtime="00:02:26.83" resultid="7228" heatid="7485" lane="2" entrytime="00:02:23.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:11.14" />
                    <SPLIT distance="150" swimtime="00:01:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="464" swimtime="00:02:20.87" resultid="7229" heatid="7571" lane="5" entrytime="00:02:27.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:06.97" />
                    <SPLIT distance="150" swimtime="00:01:43.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="565" swimtime="00:01:07.24" resultid="7230" heatid="7611" lane="5" entrytime="00:01:05.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1436" points="446" swimtime="00:00:28.53" resultid="7231" heatid="7645" lane="5" entrytime="00:00:27.40" />
                <RESULT eventid="1662" points="549" swimtime="00:00:30.82" resultid="7232" heatid="7813" lane="5" entrytime="00:00:29.85" />
                <RESULT eventid="1710" points="499" reactiontime="+81" swimtime="00:04:28.23" resultid="7233" heatid="8058" lane="6" entrytime="00:04:27.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                    <SPLIT distance="100" swimtime="00:01:03.10" />
                    <SPLIT distance="150" swimtime="00:01:36.69" />
                    <SPLIT distance="200" swimtime="00:02:10.78" />
                    <SPLIT distance="250" swimtime="00:02:45.41" />
                    <SPLIT distance="300" swimtime="00:03:20.30" />
                    <SPLIT distance="350" swimtime="00:03:54.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Sylwia" gender="F" lastname="Wnuk " nation="POL" license="100611100197" athleteid="7252">
              <RESULTS>
                <RESULT eventid="1058" points="548" reactiontime="+77" swimtime="00:00:28.41" resultid="7253" heatid="7332" lane="6" />
                <RESULT eventid="1285" points="614" reactiontime="+72" swimtime="00:01:07.93" resultid="7254" heatid="7537" lane="3" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="547" reactiontime="+91" swimtime="00:01:16.63" resultid="7255" heatid="7581" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1419" points="509" reactiontime="+74" swimtime="00:00:30.52" resultid="7256" heatid="7621" lane="4" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-10-09" firstname="Arkadiusz" gender="M" lastname="Kula" nation="POL" athleteid="7944">
              <RESULTS>
                <RESULT eventid="1165" points="446" reactiontime="+83" swimtime="00:18:32.33" resultid="7945" heatid="7917" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="100" swimtime="00:01:04.10" />
                    <SPLIT distance="150" swimtime="00:01:39.67" />
                    <SPLIT distance="200" swimtime="00:02:15.99" />
                    <SPLIT distance="250" swimtime="00:02:52.73" />
                    <SPLIT distance="300" swimtime="00:03:29.63" />
                    <SPLIT distance="350" swimtime="00:04:06.53" />
                    <SPLIT distance="400" swimtime="00:04:43.65" />
                    <SPLIT distance="450" swimtime="00:05:21.15" />
                    <SPLIT distance="500" swimtime="00:05:58.35" />
                    <SPLIT distance="550" swimtime="00:06:36.74" />
                    <SPLIT distance="600" swimtime="00:07:14.96" />
                    <SPLIT distance="650" swimtime="00:07:53.63" />
                    <SPLIT distance="700" swimtime="00:08:32.31" />
                    <SPLIT distance="750" swimtime="00:09:11.00" />
                    <SPLIT distance="800" swimtime="00:09:48.70" />
                    <SPLIT distance="850" swimtime="00:10:26.39" />
                    <SPLIT distance="900" swimtime="00:11:04.05" />
                    <SPLIT distance="950" swimtime="00:11:41.17" />
                    <SPLIT distance="1000" swimtime="00:12:19.84" />
                    <SPLIT distance="1050" swimtime="00:12:57.69" />
                    <SPLIT distance="1100" swimtime="00:13:35.02" />
                    <SPLIT distance="1150" swimtime="00:14:12.24" />
                    <SPLIT distance="1200" swimtime="00:14:49.71" />
                    <SPLIT distance="1250" swimtime="00:15:27.57" />
                    <SPLIT distance="1300" swimtime="00:16:04.72" />
                    <SPLIT distance="1350" swimtime="00:16:42.96" />
                    <SPLIT distance="1400" swimtime="00:17:20.24" />
                    <SPLIT distance="1450" swimtime="00:17:57.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="AZS UŚ Katowice" nation="POL" region="SLA">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1950-09-19" firstname="Wiesław" gender="M" lastname="Majcher" nation="POL" athleteid="7235">
              <RESULTS>
                <RESULT comment="O-4 - Start wykonany przed sygnałem (Przedwczesny start)" eventid="1075" reactiontime="+56" status="DSQ" swimtime="00:00:41.14" resultid="7236" heatid="7347" lane="6" />
                <RESULT eventid="1165" points="61" reactiontime="+115" swimtime="00:35:56.33" resultid="7237" heatid="7907" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.49" />
                    <SPLIT distance="100" swimtime="00:03:06.97" />
                    <SPLIT distance="150" swimtime="00:04:15.19" />
                    <SPLIT distance="200" swimtime="00:05:26.80" />
                    <SPLIT distance="250" swimtime="00:06:39.23" />
                    <SPLIT distance="300" swimtime="00:07:43.52" />
                    <SPLIT distance="350" swimtime="00:09:01.57" />
                    <SPLIT distance="400" swimtime="00:10:21.28" />
                    <SPLIT distance="450" swimtime="00:11:32.57" />
                    <SPLIT distance="500" swimtime="00:12:51.56" />
                    <SPLIT distance="550" swimtime="00:14:03.33" />
                    <SPLIT distance="600" swimtime="00:15:21.67" />
                    <SPLIT distance="650" swimtime="00:19:02.95" />
                    <SPLIT distance="700" swimtime="00:20:16.34" />
                    <SPLIT distance="750" swimtime="00:21:27.52" />
                    <SPLIT distance="800" swimtime="00:22:47.40" />
                    <SPLIT distance="850" swimtime="00:23:56.23" />
                    <SPLIT distance="900" swimtime="00:25:03.53" />
                    <SPLIT distance="950" swimtime="00:26:12.63" />
                    <SPLIT distance="1000" swimtime="00:27:31.08" />
                    <SPLIT distance="1050" swimtime="00:28:39.90" />
                    <SPLIT distance="1100" swimtime="00:30:00.33" />
                    <SPLIT distance="1150" swimtime="00:31:17.18" />
                    <SPLIT distance="1200" swimtime="00:32:20.26" />
                    <SPLIT distance="1250" swimtime="00:33:37.47" />
                    <SPLIT distance="1300" swimtime="00:34:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="7238" heatid="7470" lane="5" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="7239" heatid="7538" lane="3" />
                <RESULT eventid="1436" points="64" reactiontime="+102" swimtime="00:00:54.40" resultid="7240" heatid="7622" lane="2" />
                <RESULT eventid="1504" points="87" reactiontime="+111" swimtime="00:03:43.45" resultid="7241" heatid="7686" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.99" />
                    <SPLIT distance="100" swimtime="00:01:45.53" />
                    <SPLIT distance="150" swimtime="00:02:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1710" status="DNS" swimtime="00:00:00.00" resultid="7242" heatid="8043" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Beskidzkie WOPR" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Przemysław " gender="M" lastname="Pobóg-Zarzecki " nation="POL" athleteid="7313">
              <RESULTS>
                <RESULT comment="O-15 - Brak kontaktu ze ścianą nawrotową (na 50 metrze)" eventid="1268" reactiontime="+81" status="DSQ" swimtime="00:01:13.30" resultid="7314" heatid="7504" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="7315" heatid="7600" lane="4" entrytime="00:01:30.00" />
                <RESULT eventid="1662" status="DNS" swimtime="00:00:00.00" resultid="7316" heatid="7803" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02711" name="CSiR MOS Dąbrowa Górnicza" nation="POL" region="SLA">
          <CONTACT name="Waliczek mariusz" phone="606448210" />
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

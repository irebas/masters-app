<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Warmińsko-Mazurski Okręgowy Związek Pływacki" version="11.45285">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" phone="+41 99 999 99 99" fax="+41 99 999 99 99" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Olsztyn" name="Zimowe Mistrzostwa Polski w Pływaniu w kategorii Masters" name.en="Letnie Mistrzostwa Polski w Plywaniu Masters" course="SCM" deadline="2016-10-10" nation="POL" organizer="Masters Olsztyn" result.url="http://www.megatiming.pl" startmethod="1" timing="AUTOMATIC">
      <AGEDATE value="2016-12-31" type="YEAR" />
      <POOL name="OSIR Aquasfera Olsztyn" lanemax="9" />
      <POINTTABLE pointtableid="3009" name="FINA Point Scoring" version="2016" />
      <CONTACT email="zawody.olsztyn@interia.pl" name="Elżbieta Chodyna" phone="600215732" />
      <FEES>
        <FEE currency="PLN" type="ATHLETE" value="10000" />
        <FEE currency="PLN" type="LATEENTRY.INDIVIDUAL" value="15000" />
      </FEES>
      <SESSIONS>
        <SESSION date="2016-10-21" daytime="14:00" number="1" warmupfrom="12:45" warmupuntil="13:40">
          <EVENTS>
            <EVENT eventid="98814" daytime="14:48" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99692" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107940" />
                    <RANKING order="2" place="2" resultid="108637" />
                    <RANKING order="3" place="3" resultid="107370" />
                    <RANKING order="4" place="4" resultid="108673" />
                    <RANKING order="5" place="5" resultid="110373" />
                    <RANKING order="6" place="-1" resultid="108955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99693" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108216" />
                    <RANKING order="2" place="2" resultid="109986" />
                    <RANKING order="3" place="3" resultid="110276" />
                    <RANKING order="4" place="4" resultid="108904" />
                    <RANKING order="5" place="-1" resultid="106798" />
                    <RANKING order="6" place="-1" resultid="108644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99694" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107226" />
                    <RANKING order="2" place="2" resultid="107482" />
                    <RANKING order="3" place="3" resultid="108622" />
                    <RANKING order="4" place="4" resultid="107870" />
                    <RANKING order="5" place="5" resultid="106987" />
                    <RANKING order="6" place="6" resultid="107836" />
                    <RANKING order="7" place="7" resultid="107031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99695" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108267" />
                    <RANKING order="2" place="2" resultid="107705" />
                    <RANKING order="3" place="3" resultid="108680" />
                    <RANKING order="4" place="4" resultid="109016" />
                    <RANKING order="5" place="5" resultid="109927" />
                    <RANKING order="6" place="6" resultid="106593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99696" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108084" />
                    <RANKING order="2" place="2" resultid="106982" />
                    <RANKING order="3" place="3" resultid="106425" />
                    <RANKING order="4" place="4" resultid="110135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99697" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108078" />
                    <RANKING order="2" place="2" resultid="108432" />
                    <RANKING order="3" place="3" resultid="109822" />
                    <RANKING order="4" place="4" resultid="107039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99698" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108525" />
                    <RANKING order="2" place="2" resultid="108040" />
                    <RANKING order="3" place="3" resultid="107987" />
                    <RANKING order="4" place="4" resultid="109544" />
                    <RANKING order="5" place="-1" resultid="106758" />
                    <RANKING order="6" place="-1" resultid="110102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99699" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107089" />
                    <RANKING order="2" place="2" resultid="109527" />
                    <RANKING order="3" place="3" resultid="106958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99700" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107903" />
                    <RANKING order="2" place="-1" resultid="106747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99701" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108092" />
                    <RANKING order="2" place="2" resultid="110094" />
                    <RANKING order="3" place="3" resultid="110472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99702" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99703" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99704" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99705" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99706" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110614" daytime="14:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110615" daytime="14:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110616" daytime="15:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110617" daytime="15:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110618" daytime="15:09" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="106256" daytime="18:41" gender="M" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="106257" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106258" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106398" />
                    <RANKING order="2" place="2" resultid="109003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106259" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107509" />
                    <RANKING order="2" place="2" resultid="110856" />
                    <RANKING order="3" place="-1" resultid="106638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106260" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109553" />
                    <RANKING order="2" place="2" resultid="108408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106261" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107743" />
                    <RANKING order="2" place="2" resultid="108996" />
                    <RANKING order="3" place="3" resultid="109139" />
                    <RANKING order="4" place="-1" resultid="109882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106262" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106877" />
                    <RANKING order="2" place="2" resultid="107686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106263" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106998" />
                    <RANKING order="2" place="2" resultid="109165" />
                    <RANKING order="3" place="3" resultid="106611" />
                    <RANKING order="4" place="4" resultid="110408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106264" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108022" />
                    <RANKING order="2" place="2" resultid="109855" />
                    <RANKING order="3" place="3" resultid="110489" />
                    <RANKING order="4" place="4" resultid="106831" />
                    <RANKING order="5" place="-1" resultid="106837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106265" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106411" />
                    <RANKING order="2" place="2" resultid="107097" />
                    <RANKING order="3" place="3" resultid="108155" />
                    <RANKING order="4" place="-1" resultid="110500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106266" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109378" />
                    <RANKING order="2" place="2" resultid="108164" />
                    <RANKING order="3" place="3" resultid="107789" />
                    <RANKING order="4" place="4" resultid="109996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106267" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="106268" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106269" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="106270" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="106271" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110641" daytime="18:41" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110642" daytime="19:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110643" daytime="19:27" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110644" daytime="20:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98798" daytime="14:16" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99677" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107111" />
                    <RANKING order="2" place="2" resultid="107541" />
                    <RANKING order="3" place="3" resultid="109212" />
                    <RANKING order="4" place="4" resultid="109534" />
                    <RANKING order="5" place="5" resultid="107104" />
                    <RANKING order="6" place="6" resultid="110530" />
                    <RANKING order="7" place="7" resultid="110551" />
                    <RANKING order="8" place="8" resultid="106672" />
                    <RANKING order="9" place="9" resultid="108702" />
                    <RANKING order="10" place="10" resultid="108689" />
                    <RANKING order="11" place="-1" resultid="107923" />
                    <RANKING order="12" place="-1" resultid="108945" />
                    <RANKING order="13" place="-1" resultid="109311" />
                    <RANKING order="14" place="-1" resultid="110507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99678" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107187" />
                    <RANKING order="2" place="2" resultid="109888" />
                    <RANKING order="3" place="3" resultid="106440" />
                    <RANKING order="4" place="4" resultid="107176" />
                    <RANKING order="5" place="5" resultid="106653" />
                    <RANKING order="6" place="6" resultid="110142" />
                    <RANKING order="7" place="7" resultid="107246" />
                    <RANKING order="8" place="8" resultid="109473" />
                    <RANKING order="9" place="9" resultid="107180" />
                    <RANKING order="10" place="9" resultid="107720" />
                    <RANKING order="11" place="11" resultid="110381" />
                    <RANKING order="12" place="12" resultid="107629" />
                    <RANKING order="13" place="13" resultid="107848" />
                    <RANKING order="14" place="14" resultid="107223" />
                    <RANKING order="15" place="15" resultid="106605" />
                    <RANKING order="16" place="16" resultid="107877" />
                    <RANKING order="17" place="17" resultid="109940" />
                    <RANKING order="18" place="18" resultid="108696" />
                    <RANKING order="19" place="19" resultid="110370" />
                    <RANKING order="20" place="20" resultid="107193" />
                    <RANKING order="21" place="21" resultid="107677" />
                    <RANKING order="22" place="-1" resultid="106648" />
                    <RANKING order="23" place="-1" resultid="107212" />
                    <RANKING order="24" place="-1" resultid="110578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99679" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107199" />
                    <RANKING order="2" place="2" resultid="107391" />
                    <RANKING order="3" place="3" resultid="107397" />
                    <RANKING order="4" place="3" resultid="107414" />
                    <RANKING order="5" place="5" resultid="108649" />
                    <RANKING order="6" place="6" resultid="107406" />
                    <RANKING order="7" place="7" resultid="108570" />
                    <RANKING order="8" place="8" resultid="107117" />
                    <RANKING order="9" place="9" resultid="108629" />
                    <RANKING order="10" place="10" resultid="107502" />
                    <RANKING order="11" place="10" resultid="107608" />
                    <RANKING order="12" place="12" resultid="110419" />
                    <RANKING order="13" place="13" resultid="109831" />
                    <RANKING order="14" place="14" resultid="109353" />
                    <RANKING order="15" place="15" resultid="106637" />
                    <RANKING order="16" place="16" resultid="110457" />
                    <RANKING order="17" place="17" resultid="109842" />
                    <RANKING order="18" place="18" resultid="107475" />
                    <RANKING order="19" place="19" resultid="108708" />
                    <RANKING order="20" place="20" resultid="108212" />
                    <RANKING order="21" place="21" resultid="107195" />
                    <RANKING order="22" place="-1" resultid="106945" />
                    <RANKING order="23" place="-1" resultid="107619" />
                    <RANKING order="24" place="-1" resultid="108710" />
                    <RANKING order="25" place="-1" resultid="109819" />
                    <RANKING order="26" place="-1" resultid="107021" />
                    <RANKING order="27" place="-1" resultid="109458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99680" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107663" />
                    <RANKING order="2" place="2" resultid="108048" />
                    <RANKING order="3" place="2" resultid="109440" />
                    <RANKING order="4" place="4" resultid="107183" />
                    <RANKING order="5" place="5" resultid="106579" />
                    <RANKING order="6" place="6" resultid="109561" />
                    <RANKING order="7" place="7" resultid="107724" />
                    <RANKING order="8" place="8" resultid="107553" />
                    <RANKING order="9" place="9" resultid="107570" />
                    <RANKING order="10" place="10" resultid="109148" />
                    <RANKING order="11" place="11" resultid="107598" />
                    <RANKING order="12" place="12" resultid="107580" />
                    <RANKING order="13" place="13" resultid="110244" />
                    <RANKING order="14" place="14" resultid="107625" />
                    <RANKING order="15" place="15" resultid="107436" />
                    <RANKING order="16" place="16" resultid="106631" />
                    <RANKING order="17" place="17" resultid="107603" />
                    <RANKING order="18" place="18" resultid="107615" />
                    <RANKING order="19" place="19" resultid="108591" />
                    <RANKING order="20" place="20" resultid="107948" />
                    <RANKING order="21" place="-1" resultid="107575" />
                    <RANKING order="22" place="-1" resultid="107589" />
                    <RANKING order="23" place="-1" resultid="107694" />
                    <RANKING order="24" place="-1" resultid="109073" />
                    <RANKING order="25" place="-1" resultid="109933" />
                    <RANKING order="26" place="-1" resultid="106889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99681" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109031" />
                    <RANKING order="2" place="2" resultid="109863" />
                    <RANKING order="3" place="3" resultid="108970" />
                    <RANKING order="4" place="4" resultid="107843" />
                    <RANKING order="5" place="5" resultid="106572" />
                    <RANKING order="6" place="6" resultid="108398" />
                    <RANKING order="7" place="7" resultid="110120" />
                    <RANKING order="8" place="8" resultid="108416" />
                    <RANKING order="9" place="9" resultid="107965" />
                    <RANKING order="10" place="10" resultid="108979" />
                    <RANKING order="11" place="11" resultid="108553" />
                    <RANKING order="12" place="12" resultid="108989" />
                    <RANKING order="13" place="13" resultid="108558" />
                    <RANKING order="14" place="14" resultid="108658" />
                    <RANKING order="15" place="14" resultid="110192" />
                    <RANKING order="16" place="16" resultid="108995" />
                    <RANKING order="17" place="17" resultid="109881" />
                    <RANKING order="18" place="18" resultid="109138" />
                    <RANKING order="19" place="19" resultid="107216" />
                    <RANKING order="20" place="20" resultid="108248" />
                    <RANKING order="21" place="21" resultid="109959" />
                    <RANKING order="22" place="22" resultid="107214" />
                    <RANKING order="23" place="-1" resultid="107251" />
                    <RANKING order="24" place="-1" resultid="110185" />
                    <RANKING order="25" place="-1" resultid="110393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99682" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110255" />
                    <RANKING order="2" place="2" resultid="110269" />
                    <RANKING order="3" place="3" resultid="107930" />
                    <RANKING order="4" place="4" resultid="108370" />
                    <RANKING order="5" place="5" resultid="108423" />
                    <RANKING order="6" place="6" resultid="109009" />
                    <RANKING order="7" place="7" resultid="110162" />
                    <RANKING order="8" place="8" resultid="107135" />
                    <RANKING order="9" place="9" resultid="109943" />
                    <RANKING order="10" place="10" resultid="107866" />
                    <RANKING order="11" place="11" resultid="107149" />
                    <RANKING order="12" place="12" resultid="110426" />
                    <RANKING order="13" place="-1" resultid="106948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99683" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109058" />
                    <RANKING order="2" place="2" resultid="110479" />
                    <RANKING order="3" place="3" resultid="106862" />
                    <RANKING order="4" place="4" resultid="109067" />
                    <RANKING order="5" place="5" resultid="109398" />
                    <RANKING order="6" place="6" resultid="106997" />
                    <RANKING order="7" place="7" resultid="109513" />
                    <RANKING order="8" place="8" resultid="106844" />
                    <RANKING order="9" place="9" resultid="108918" />
                    <RANKING order="10" place="10" resultid="110407" />
                    <RANKING order="11" place="-1" resultid="108180" />
                    <RANKING order="12" place="-1" resultid="106871" />
                    <RANKING order="13" place="-1" resultid="110085" />
                    <RANKING order="14" place="-1" resultid="110252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99684" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109845" />
                    <RANKING order="2" place="2" resultid="109973" />
                    <RANKING order="3" place="3" resultid="108206" />
                    <RANKING order="4" place="4" resultid="108440" />
                    <RANKING order="5" place="5" resultid="107006" />
                    <RANKING order="6" place="6" resultid="110488" />
                    <RANKING order="7" place="7" resultid="110076" />
                    <RANKING order="8" place="8" resultid="106824" />
                    <RANKING order="9" place="9" resultid="108225" />
                    <RANKING order="10" place="10" resultid="109390" />
                    <RANKING order="11" place="11" resultid="106830" />
                    <RANKING order="12" place="-1" resultid="109362" />
                    <RANKING order="13" place="-1" resultid="106836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99685" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109407" />
                    <RANKING order="2" place="2" resultid="110539" />
                    <RANKING order="3" place="3" resultid="107761" />
                    <RANKING order="4" place="4" resultid="107490" />
                    <RANKING order="5" place="5" resultid="110448" />
                    <RANKING order="6" place="6" resultid="107497" />
                    <RANKING order="7" place="7" resultid="108069" />
                    <RANKING order="8" place="8" resultid="108253" />
                    <RANKING order="9" place="9" resultid="108575" />
                    <RANKING order="10" place="-1" resultid="106819" />
                    <RANKING order="11" place="-1" resultid="107972" />
                    <RANKING order="12" place="-1" resultid="110499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99686" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106405" />
                    <RANKING order="2" place="2" resultid="106705" />
                    <RANKING order="3" place="3" resultid="109377" />
                    <RANKING order="4" place="4" resultid="108030" />
                    <RANKING order="5" place="5" resultid="108530" />
                    <RANKING order="6" place="6" resultid="106806" />
                    <RANKING order="7" place="7" resultid="107788" />
                    <RANKING order="8" place="8" resultid="108008" />
                    <RANKING order="9" place="9" resultid="109468" />
                    <RANKING order="10" place="10" resultid="106716" />
                    <RANKING order="11" place="11" resultid="110147" />
                    <RANKING order="12" place="12" resultid="108360" />
                    <RANKING order="13" place="13" resultid="106813" />
                    <RANKING order="14" place="14" resultid="109995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99687" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107771" />
                    <RANKING order="2" place="2" resultid="110054" />
                    <RANKING order="3" place="3" resultid="109413" />
                    <RANKING order="4" place="4" resultid="110516" />
                    <RANKING order="5" place="5" resultid="107143" />
                    <RANKING order="6" place="6" resultid="107457" />
                    <RANKING order="7" place="7" resultid="108519" />
                    <RANKING order="8" place="8" resultid="108583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99688" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106687" />
                    <RANKING order="2" place="2" resultid="107448" />
                    <RANKING order="3" place="3" resultid="108479" />
                    <RANKING order="4" place="4" resultid="108511" />
                    <RANKING order="5" place="5" resultid="107454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99689" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99690" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99691" agemax="94" agemin="90" name="KAT.N, 90-94 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="108004" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110594" daytime="14:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110595" daytime="14:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110596" daytime="14:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110597" daytime="14:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110598" daytime="14:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110599" daytime="14:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110600" daytime="14:27" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110601" daytime="14:29" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110602" daytime="14:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="110603" daytime="14:32" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="110604" daytime="14:33" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="110605" daytime="14:35" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="110606" daytime="14:36" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="110607" daytime="14:38" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="110608" daytime="14:39" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="110609" daytime="14:41" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="110610" daytime="14:42" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="110611" daytime="14:44" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="110612" daytime="14:45" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="110613" daytime="14:47" number="20" order="20" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98777" daytime="14:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="98779" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107369" />
                    <RANKING order="2" place="2" resultid="107939" />
                    <RANKING order="3" place="3" resultid="108636" />
                    <RANKING order="4" place="4" resultid="108672" />
                    <RANKING order="5" place="5" resultid="110372" />
                    <RANKING order="6" place="6" resultid="110402" />
                    <RANKING order="7" place="7" resultid="107122" />
                    <RANKING order="8" place="-1" resultid="108954" />
                    <RANKING order="9" place="-1" resultid="110440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98780" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106797" />
                    <RANKING order="2" place="2" resultid="106665" />
                    <RANKING order="3" place="3" resultid="108215" />
                    <RANKING order="4" place="4" resultid="107672" />
                    <RANKING order="5" place="5" resultid="110284" />
                    <RANKING order="6" place="6" resultid="107207" />
                    <RANKING order="7" place="7" resultid="107260" />
                    <RANKING order="8" place="8" resultid="107378" />
                    <RANKING order="9" place="-1" resultid="107202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98782" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106586" />
                    <RANKING order="2" place="2" resultid="108621" />
                    <RANKING order="3" place="3" resultid="110295" />
                    <RANKING order="4" place="4" resultid="109048" />
                    <RANKING order="5" place="5" resultid="106433" />
                    <RANKING order="6" place="-1" resultid="107218" />
                    <RANKING order="7" place="-1" resultid="108667" />
                    <RANKING order="8" place="-1" resultid="109872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98783" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108266" />
                    <RANKING order="2" place="2" resultid="107704" />
                    <RANKING order="3" place="3" resultid="107713" />
                    <RANKING order="4" place="4" resultid="109926" />
                    <RANKING order="5" place="5" resultid="108963" />
                    <RANKING order="6" place="6" resultid="106429" />
                    <RANKING order="7" place="7" resultid="106790" />
                    <RANKING order="8" place="8" resultid="110303" />
                    <RANKING order="9" place="9" resultid="110179" />
                    <RANKING order="10" place="10" resultid="106592" />
                    <RANKING order="11" place="11" resultid="110237" />
                    <RANKING order="12" place="-1" resultid="106643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98781" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108083" />
                    <RANKING order="2" place="2" resultid="110128" />
                    <RANKING order="3" place="3" resultid="109837" />
                    <RANKING order="4" place="4" resultid="107464" />
                    <RANKING order="5" place="-1" resultid="107915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98785" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108564" />
                    <RANKING order="2" place="2" resultid="106779" />
                    <RANKING order="3" place="3" resultid="107854" />
                    <RANKING order="4" place="4" resultid="109912" />
                    <RANKING order="5" place="-1" resultid="108431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98784" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108495" />
                    <RANKING order="2" place="2" resultid="108013" />
                    <RANKING order="3" place="3" resultid="107986" />
                    <RANKING order="4" place="4" resultid="108039" />
                    <RANKING order="5" place="5" resultid="106773" />
                    <RANKING order="6" place="6" resultid="109543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98787" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108502" />
                    <RANKING order="2" place="2" resultid="109526" />
                    <RANKING order="3" place="3" resultid="106753" />
                    <RANKING order="4" place="4" resultid="110220" />
                    <RANKING order="5" place="5" resultid="106957" />
                    <RANKING order="6" place="6" resultid="110170" />
                    <RANKING order="7" place="7" resultid="108454" />
                    <RANKING order="8" place="8" resultid="110229" />
                    <RANKING order="9" place="-1" resultid="108394" />
                    <RANKING order="10" place="-1" resultid="108385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98786" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108062" />
                    <RANKING order="2" place="2" resultid="107469" />
                    <RANKING order="3" place="3" resultid="107902" />
                    <RANKING order="4" place="4" resultid="110354" />
                    <RANKING order="5" place="-1" resultid="106746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98789" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110093" />
                    <RANKING order="2" place="2" resultid="109452" />
                    <RANKING order="3" place="3" resultid="106720" />
                    <RANKING order="4" place="4" resultid="108091" />
                    <RANKING order="5" place="5" resultid="108468" />
                    <RANKING order="6" place="6" resultid="106942" />
                    <RANKING order="7" place="7" resultid="109429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98788" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106692" />
                    <RANKING order="2" place="2" resultid="108539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98791" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106741" />
                    <RANKING order="2" place="2" resultid="107812" />
                    <RANKING order="3" place="3" resultid="109130" />
                    <RANKING order="4" place="-1" resultid="107798" />
                    <RANKING order="5" place="-1" resultid="107805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98793" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="98792" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="98795" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110585" daytime="14:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110586" daytime="14:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110587" daytime="14:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110588" daytime="14:07" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110589" daytime="14:09" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110590" daytime="14:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110591" daytime="14:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110592" daytime="14:13" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110593" daytime="14:15" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98830" daytime="15:13" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99707" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107542" />
                    <RANKING order="2" place="2" resultid="109535" />
                    <RANKING order="3" place="3" resultid="110552" />
                    <RANKING order="4" place="4" resultid="109901" />
                    <RANKING order="5" place="5" resultid="110531" />
                    <RANKING order="6" place="6" resultid="110431" />
                    <RANKING order="7" place="7" resultid="108690" />
                    <RANKING order="8" place="8" resultid="110558" />
                    <RANKING order="9" place="-1" resultid="108946" />
                    <RANKING order="10" place="-1" resultid="110508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99708" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107188" />
                    <RANKING order="2" place="2" resultid="107168" />
                    <RANKING order="3" place="3" resultid="106658" />
                    <RANKING order="4" place="4" resultid="109474" />
                    <RANKING order="5" place="5" resultid="110287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99709" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107415" />
                    <RANKING order="2" place="2" resultid="106973" />
                    <RANKING order="3" place="3" resultid="109573" />
                    <RANKING order="4" place="4" resultid="108650" />
                    <RANKING order="5" place="5" resultid="107562" />
                    <RANKING order="6" place="6" resultid="107398" />
                    <RANKING order="7" place="7" resultid="107609" />
                    <RANKING order="8" place="8" resultid="109965" />
                    <RANKING order="9" place="9" resultid="109354" />
                    <RANKING order="10" place="10" resultid="110420" />
                    <RANKING order="11" place="11" resultid="110458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99710" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109552" />
                    <RANKING order="2" place="2" resultid="107664" />
                    <RANKING order="3" place="3" resultid="108049" />
                    <RANKING order="4" place="4" resultid="109606" />
                    <RANKING order="5" place="5" resultid="106966" />
                    <RANKING order="6" place="6" resultid="107590" />
                    <RANKING order="7" place="7" resultid="110245" />
                    <RANKING order="8" place="8" resultid="107581" />
                    <RANKING order="9" place="9" resultid="107949" />
                    <RANKING order="10" place="-1" resultid="108407" />
                    <RANKING order="11" place="-1" resultid="109952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99711" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109864" />
                    <RANKING order="2" place="2" resultid="108417" />
                    <RANKING order="3" place="3" resultid="108399" />
                    <RANKING order="4" place="4" resultid="108971" />
                    <RANKING order="5" place="5" resultid="109337" />
                    <RANKING order="6" place="6" resultid="107742" />
                    <RANKING order="7" place="7" resultid="106700" />
                    <RANKING order="8" place="8" resultid="110154" />
                    <RANKING order="9" place="9" resultid="110394" />
                    <RANKING order="10" place="10" resultid="108659" />
                    <RANKING order="11" place="-1" resultid="108980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99712" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109024" />
                    <RANKING order="2" place="2" resultid="107735" />
                    <RANKING order="3" place="3" resultid="110270" />
                    <RANKING order="4" place="4" resultid="106883" />
                    <RANKING order="5" place="5" resultid="107830" />
                    <RANKING order="6" place="6" resultid="107752" />
                    <RANKING order="7" place="7" resultid="108371" />
                    <RANKING order="8" place="8" resultid="107685" />
                    <RANKING order="9" place="9" resultid="107150" />
                    <RANKING order="10" place="-1" resultid="106949" />
                    <RANKING order="11" place="-1" resultid="110163" />
                    <RANKING order="12" place="-1" resultid="110256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99713" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109399" />
                    <RANKING order="2" place="2" resultid="109059" />
                    <RANKING order="3" place="3" resultid="110480" />
                    <RANKING order="4" place="4" resultid="110263" />
                    <RANKING order="5" place="5" resultid="109567" />
                    <RANKING order="6" place="6" resultid="106610" />
                    <RANKING order="7" place="7" resultid="108181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99714" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107025" />
                    <RANKING order="2" place="2" resultid="108441" />
                    <RANKING order="3" place="3" resultid="109854" />
                    <RANKING order="4" place="4" resultid="110077" />
                    <RANKING order="5" place="5" resultid="109317" />
                    <RANKING order="6" place="-1" resultid="108021" />
                    <RANKING order="7" place="-1" resultid="109363" />
                    <RANKING order="8" place="-1" resultid="108226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99715" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107127" />
                    <RANKING order="2" place="2" resultid="110067" />
                    <RANKING order="3" place="3" resultid="107096" />
                    <RANKING order="4" place="4" resultid="108201" />
                    <RANKING order="5" place="5" resultid="108154" />
                    <RANKING order="6" place="6" resultid="107491" />
                    <RANKING order="7" place="7" resultid="108070" />
                    <RANKING order="8" place="-1" resultid="108233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99716" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109371" />
                    <RANKING order="2" place="2" resultid="106937" />
                    <RANKING order="3" place="3" resultid="106807" />
                    <RANKING order="4" place="4" resultid="108531" />
                    <RANKING order="5" place="5" resultid="108031" />
                    <RANKING order="6" place="6" resultid="108163" />
                    <RANKING order="7" place="7" resultid="110148" />
                    <RANKING order="8" place="8" resultid="110362" />
                    <RANKING order="9" place="9" resultid="107440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99717" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107772" />
                    <RANKING order="2" place="2" resultid="110055" />
                    <RANKING order="3" place="3" resultid="108584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99718" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108480" />
                    <RANKING order="2" place="2" resultid="108172" />
                    <RANKING order="3" place="-1" resultid="109345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99719" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99720" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99721" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110619" daytime="15:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110620" daytime="15:19" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110621" daytime="15:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110622" daytime="15:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110623" daytime="15:33" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110624" daytime="15:37" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110625" daytime="15:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110626" daytime="15:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110627" daytime="15:48" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="110628" daytime="15:51" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98846" daytime="15:55" gender="X" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="98847" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="108716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98848" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107271" />
                    <RANKING order="2" place="-1" resultid="106677" />
                    <RANKING order="3" place="-1" resultid="107261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98849" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107731" />
                    <RANKING order="2" place="2" resultid="109998" />
                    <RANKING order="3" place="3" resultid="107422" />
                    <RANKING order="4" place="4" resultid="106620" />
                    <RANKING order="5" place="5" resultid="107522" />
                    <RANKING order="6" place="6" resultid="108712" />
                    <RANKING order="7" place="7" resultid="106993" />
                    <RANKING order="8" place="8" resultid="107887" />
                    <RANKING order="9" place="-1" resultid="107262" />
                    <RANKING order="10" place="-1" resultid="106492" />
                    <RANKING order="11" place="-1" resultid="108714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98850" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108601" />
                    <RANKING order="2" place="2" resultid="106893" />
                    <RANKING order="3" place="3" resultid="109036" />
                    <RANKING order="4" place="4" resultid="108097" />
                    <RANKING order="5" place="5" resultid="107885" />
                    <RANKING order="6" place="6" resultid="110196" />
                    <RANKING order="7" place="7" resultid="109999" />
                    <RANKING order="8" place="8" resultid="110197" />
                    <RANKING order="9" place="9" resultid="107956" />
                    <RANKING order="10" place="-1" resultid="110254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98851" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108099" />
                    <RANKING order="2" place="2" resultid="106892" />
                    <RANKING order="3" place="3" resultid="110000" />
                    <RANKING order="4" place="4" resultid="108597" />
                    <RANKING order="5" place="5" resultid="109585" />
                    <RANKING order="6" place="-1" resultid="110109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98852" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110584" />
                    <RANKING order="2" place="2" resultid="108101" />
                    <RANKING order="3" place="3" resultid="108491" />
                    <RANKING order="4" place="4" resultid="110001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98853" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106725" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110629" daytime="15:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110630" daytime="15:59" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110631" daytime="16:03" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110632" daytime="16:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98863" daytime="16:09" gender="F" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99722" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99723" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109987" />
                    <RANKING order="2" place="2" resultid="110277" />
                    <RANKING order="3" place="3" resultid="108905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99724" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109921" />
                    <RANKING order="2" place="2" resultid="110296" />
                    <RANKING order="3" place="3" resultid="107386" />
                    <RANKING order="4" place="4" resultid="106434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99725" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99726" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99727" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109823" />
                    <RANKING order="2" place="2" resultid="109913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99728" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99729" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108503" />
                    <RANKING order="2" place="2" resultid="110221" />
                    <RANKING order="3" place="3" resultid="109977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99730" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99731" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99732" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99733" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99734" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99735" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99736" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110633" daytime="16:09" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110634" daytime="16:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="106254" daytime="18:04" gender="F" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="106311" agemax="24" agemin="20" name="KAT.0, 20-24 lat" />
                <AGEGROUP agegroupid="106312" agemax="29" agemin="25" name="KAT.A, 25-29 lat" />
                <AGEGROUP agegroupid="106313" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109873" />
                    <RANKING order="2" place="2" resultid="107032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106314" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106315" agemax="44" agemin="40" name="KAT.D, 40-44 lat" />
                <AGEGROUP agegroupid="106316" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106317" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108196" />
                    <RANKING order="2" place="2" resultid="108923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106318" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107090" />
                    <RANKING order="2" place="2" resultid="110171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106319" agemax="64" agemin="60" name="KAT.H, 60-64 lat" />
                <AGEGROUP agegroupid="106320" agemax="69" agemin="65" name="KAT.I, 65-69 lat" />
                <AGEGROUP agegroupid="106321" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="106322" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106323" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="106324" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="106325" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110640" daytime="18:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98891" daytime="16:43" gender="M" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99737" agemax="24" agemin="20" name="KAT.0, 20-24 lat" />
                <AGEGROUP agegroupid="99738" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107169" />
                    <RANKING order="2" place="2" resultid="109889" />
                    <RANKING order="3" place="3" resultid="110288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99739" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109521" />
                    <RANKING order="2" place="2" resultid="109832" />
                    <RANKING order="3" place="-1" resultid="107254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99740" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110360" />
                    <RANKING order="2" place="2" resultid="107554" />
                    <RANKING order="3" place="3" resultid="107433" />
                    <RANKING order="4" place="4" resultid="110020" />
                    <RANKING order="5" place="5" resultid="107695" />
                    <RANKING order="6" place="6" resultid="106632" />
                    <RANKING order="7" place="-1" resultid="109607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99741" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106573" />
                    <RANKING order="2" place="2" resultid="109463" />
                    <RANKING order="3" place="3" resultid="107049" />
                    <RANKING order="4" place="4" resultid="109338" />
                    <RANKING order="5" place="5" resultid="110496" />
                    <RANKING order="6" place="6" resultid="110155" />
                    <RANKING order="7" place="-1" resultid="108249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99742" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107931" />
                    <RANKING order="2" place="2" resultid="107753" />
                    <RANKING order="3" place="3" resultid="109944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99743" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109514" />
                    <RANKING order="2" place="2" resultid="106863" />
                    <RANKING order="3" place="3" resultid="106845" />
                    <RANKING order="4" place="4" resultid="109501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99744" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109846" />
                    <RANKING order="2" place="2" resultid="108207" />
                    <RANKING order="3" place="3" resultid="109318" />
                    <RANKING order="4" place="4" resultid="109391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99745" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110068" />
                    <RANKING order="2" place="2" resultid="110449" />
                    <RANKING order="3" place="3" resultid="110525" />
                    <RANKING order="4" place="-1" resultid="107762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99746" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110062" />
                    <RANKING order="2" place="2" resultid="106814" />
                    <RANKING order="3" place="3" resultid="108361" />
                    <RANKING order="4" place="4" resultid="109983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99747" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110517" />
                    <RANKING order="2" place="2" resultid="109414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99748" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99749" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99750" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99751" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110635" daytime="16:43" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110636" daytime="16:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110637" daytime="17:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110638" daytime="17:21" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110639" daytime="17:43" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-10-22" daytime="09:00" endtime="13:30" number="2" warmupfrom="08:00" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="99004" daytime="11:55" gender="F" number="18" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99005" agemax="24" agemin="20" name="KAT.0, 20-24 lat" />
                <AGEGROUP agegroupid="99006" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99007" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110298" />
                    <RANKING order="2" place="2" resultid="109875" />
                    <RANKING order="3" place="3" resultid="108624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99008" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108269" />
                    <RANKING order="2" place="-1" resultid="106644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99009" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99010" agemax="49" agemin="45" name="KAT.E, 45-49 lat" />
                <AGEGROUP agegroupid="99011" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108015" />
                    <RANKING order="2" place="2" resultid="109546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99012" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109177" />
                    <RANKING order="2" place="2" resultid="110231" />
                    <RANKING order="3" place="-1" resultid="108505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99013" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108462" />
                    <RANKING order="2" place="2" resultid="107905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99014" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108094" />
                    <RANKING order="2" place="2" resultid="110096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99015" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99016" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99017" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99018" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99019" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110707" daytime="11:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110708" daytime="12:01" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99020" daytime="12:06" gender="M" number="19" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99021" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109537" />
                    <RANKING order="2" place="2" resultid="110434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99022" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106399" />
                    <RANKING order="2" place="2" resultid="107171" />
                    <RANKING order="3" place="3" resultid="110387" />
                    <RANKING order="4" place="4" resultid="110290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99023" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107242" />
                    <RANKING order="2" place="2" resultid="106976" />
                    <RANKING order="3" place="3" resultid="107564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99024" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107235" />
                    <RANKING order="2" place="2" resultid="109555" />
                    <RANKING order="3" place="3" resultid="106968" />
                    <RANKING order="4" place="-1" resultid="108410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99025" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109340" />
                    <RANKING order="2" place="2" resultid="106701" />
                    <RANKING order="3" place="3" resultid="109140" />
                    <RANKING order="4" place="4" resultid="108998" />
                    <RANKING order="5" place="5" resultid="110573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99026" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109171" />
                    <RANKING order="2" place="2" resultid="108930" />
                    <RANKING order="3" place="3" resultid="107755" />
                    <RANKING order="4" place="-1" resultid="108425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99027" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109068" />
                    <RANKING order="2" place="2" resultid="107000" />
                    <RANKING order="3" place="3" resultid="110264" />
                    <RANKING order="4" place="4" resultid="109502" />
                    <RANKING order="5" place="5" resultid="106613" />
                    <RANKING order="6" place="-1" resultid="109435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99028" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109848" />
                    <RANKING order="2" place="2" resultid="109320" />
                    <RANKING order="3" place="3" resultid="110079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99029" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108157" />
                    <RANKING order="2" place="2" resultid="108072" />
                    <RANKING order="3" place="-1" resultid="107098" />
                    <RANKING order="4" place="-1" resultid="108235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99030" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106809" />
                    <RANKING order="2" place="2" resultid="108533" />
                    <RANKING order="3" place="3" resultid="110364" />
                    <RANKING order="4" place="4" resultid="107442" />
                    <RANKING order="5" place="-1" resultid="108033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99031" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99032" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107997" />
                    <RANKING order="2" place="2" resultid="108174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99033" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99034" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99035" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110709" daytime="12:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110710" daytime="12:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110711" daytime="12:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110712" daytime="12:23" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110713" daytime="12:27" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98907" daytime="10:18" gender="F" number="14" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99752" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107372" />
                    <RANKING order="2" place="2" resultid="107941" />
                    <RANKING order="3" place="3" resultid="110374" />
                    <RANKING order="4" place="-1" resultid="110442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99753" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106800" />
                    <RANKING order="2" place="2" resultid="106667" />
                    <RANKING order="3" place="3" resultid="110279" />
                    <RANKING order="4" place="4" resultid="107380" />
                    <RANKING order="5" place="5" resultid="109080" />
                    <RANKING order="6" place="-1" resultid="107203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99754" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109605" />
                    <RANKING order="2" place="2" resultid="106587" />
                    <RANKING order="3" place="3" resultid="110297" />
                    <RANKING order="4" place="4" resultid="109049" />
                    <RANKING order="5" place="5" resultid="106435" />
                    <RANKING order="6" place="-1" resultid="108668" />
                    <RANKING order="7" place="-1" resultid="109874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99755" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108268" />
                    <RANKING order="2" place="2" resultid="107706" />
                    <RANKING order="3" place="3" resultid="107961" />
                    <RANKING order="4" place="4" resultid="108682" />
                    <RANKING order="5" place="5" resultid="108964" />
                    <RANKING order="6" place="6" resultid="106430" />
                    <RANKING order="7" place="7" resultid="110181" />
                    <RANKING order="8" place="8" resultid="110304" />
                    <RANKING order="9" place="9" resultid="106594" />
                    <RANKING order="10" place="10" resultid="110239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99756" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107066" />
                    <RANKING order="2" place="2" resultid="110130" />
                    <RANKING order="3" place="-1" resultid="107917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99757" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108566" />
                    <RANKING order="2" place="2" resultid="106781" />
                    <RANKING order="3" place="3" resultid="109825" />
                    <RANKING order="4" place="4" resultid="109915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99758" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108924" />
                    <RANKING order="2" place="2" resultid="108041" />
                    <RANKING order="3" place="3" resultid="107989" />
                    <RANKING order="4" place="4" resultid="109508" />
                    <RANKING order="5" place="5" resultid="106774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99759" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108504" />
                    <RANKING order="2" place="2" resultid="106754" />
                    <RANKING order="3" place="3" resultid="109978" />
                    <RANKING order="4" place="4" resultid="106960" />
                    <RANKING order="5" place="5" resultid="108456" />
                    <RANKING order="6" place="-1" resultid="108395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99760" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="106749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99761" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109454" />
                    <RANKING order="2" place="2" resultid="109431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99762" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106694" />
                    <RANKING order="2" place="2" resultid="108541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99763" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106742" />
                    <RANKING order="2" place="2" resultid="107814" />
                    <RANKING order="3" place="3" resultid="107807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99764" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99765" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99766" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110671" daytime="10:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110672" daytime="10:23" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110673" daytime="10:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110674" daytime="10:29" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110675" daytime="10:31" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110676" daytime="10:33" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98956" daytime="09:50" gender="M" number="13" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99797" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110532" />
                    <RANKING order="2" place="2" resultid="110554" />
                    <RANKING order="3" place="3" resultid="108948" />
                    <RANKING order="4" place="4" resultid="110559" />
                    <RANKING order="5" place="-1" resultid="110510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99798" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109004" />
                    <RANKING order="2" place="2" resultid="110289" />
                    <RANKING order="3" place="3" resultid="110386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99799" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107510" />
                    <RANKING order="2" place="2" resultid="107256" />
                    <RANKING order="3" place="3" resultid="109966" />
                    <RANKING order="4" place="4" resultid="109522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99800" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109554" />
                    <RANKING order="2" place="2" resultid="109953" />
                    <RANKING order="3" place="3" resultid="108409" />
                    <RANKING order="4" place="4" resultid="106967" />
                    <RANKING order="5" place="5" resultid="107591" />
                    <RANKING order="6" place="6" resultid="107582" />
                    <RANKING order="7" place="7" resultid="107951" />
                    <RANKING order="8" place="-1" resultid="109074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99801" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108418" />
                    <RANKING order="2" place="2" resultid="109339" />
                    <RANKING order="3" place="3" resultid="108560" />
                    <RANKING order="4" place="4" resultid="108981" />
                    <RANKING order="5" place="-1" resultid="110186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99802" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109025" />
                    <RANKING order="2" place="2" resultid="107932" />
                    <RANKING order="3" place="3" resultid="107754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99803" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106864" />
                    <RANKING order="2" place="2" resultid="109568" />
                    <RANKING order="3" place="3" resultid="106872" />
                    <RANKING order="4" place="4" resultid="106846" />
                    <RANKING order="5" place="5" resultid="110086" />
                    <RANKING order="6" place="6" resultid="109434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99804" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107007" />
                    <RANKING order="2" place="2" resultid="110078" />
                    <RANKING order="3" place="3" resultid="109319" />
                    <RANKING order="4" place="-1" resultid="108352" />
                    <RANKING order="5" place="-1" resultid="109856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99805" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107128" />
                    <RANKING order="2" place="2" resultid="108475" />
                    <RANKING order="3" place="3" resultid="108202" />
                    <RANKING order="4" place="-1" resultid="108234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99806" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108009" />
                    <RANKING order="2" place="2" resultid="109814" />
                    <RANKING order="3" place="3" resultid="108165" />
                    <RANKING order="4" place="4" resultid="110149" />
                    <RANKING order="5" place="5" resultid="108362" />
                    <RANKING order="6" place="6" resultid="107441" />
                    <RANKING order="7" place="7" resultid="110363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99807" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107773" />
                    <RANKING order="2" place="2" resultid="107459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99808" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107996" />
                    <RANKING order="2" place="-1" resultid="109346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99809" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99810" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99811" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110665" daytime="09:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110666" daytime="09:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110667" daytime="10:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110668" daytime="10:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110669" daytime="10:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110670" daytime="10:15" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98988" daytime="11:28" gender="M" number="17" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99827" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107113" />
                    <RANKING order="2" place="2" resultid="107543" />
                    <RANKING order="3" place="3" resultid="110533" />
                    <RANKING order="4" place="4" resultid="109903" />
                    <RANKING order="5" place="5" resultid="107106" />
                    <RANKING order="6" place="6" resultid="110416" />
                    <RANKING order="7" place="7" resultid="108692" />
                    <RANKING order="8" place="8" resultid="110560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99828" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107190" />
                    <RANKING order="2" place="2" resultid="106660" />
                    <RANKING order="3" place="3" resultid="107248" />
                    <RANKING order="4" place="4" resultid="107224" />
                    <RANKING order="5" place="5" resultid="109941" />
                    <RANKING order="6" place="6" resultid="108698" />
                    <RANKING order="7" place="7" resultid="110580" />
                    <RANKING order="8" place="-1" resultid="107181" />
                    <RANKING order="9" place="-1" resultid="109476" />
                    <RANKING order="10" place="-1" resultid="110143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99829" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107241" />
                    <RANKING order="2" place="2" resultid="107417" />
                    <RANKING order="3" place="3" resultid="106975" />
                    <RANKING order="4" place="4" resultid="108652" />
                    <RANKING order="5" place="5" resultid="107393" />
                    <RANKING order="6" place="6" resultid="107119" />
                    <RANKING order="7" place="7" resultid="108572" />
                    <RANKING order="8" place="8" resultid="107610" />
                    <RANKING order="9" place="9" resultid="107408" />
                    <RANKING order="10" place="10" resultid="109967" />
                    <RANKING order="11" place="11" resultid="109356" />
                    <RANKING order="12" place="12" resultid="107477" />
                    <RANKING order="13" place="-1" resultid="109575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99830" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107666" />
                    <RANKING order="2" place="2" resultid="108051" />
                    <RANKING order="3" place="3" resultid="109442" />
                    <RANKING order="4" place="4" resultid="107184" />
                    <RANKING order="5" place="5" resultid="109954" />
                    <RANKING order="6" place="6" resultid="107556" />
                    <RANKING order="7" place="7" resultid="109609" />
                    <RANKING order="8" place="8" resultid="109150" />
                    <RANKING order="9" place="9" resultid="107592" />
                    <RANKING order="10" place="10" resultid="106581" />
                    <RANKING order="11" place="11" resultid="106601" />
                    <RANKING order="12" place="12" resultid="107437" />
                    <RANKING order="13" place="13" resultid="107583" />
                    <RANKING order="14" place="14" resultid="107604" />
                    <RANKING order="15" place="-1" resultid="107576" />
                    <RANKING order="16" place="-1" resultid="108058" />
                    <RANKING order="17" place="-1" resultid="109075" />
                    <RANKING order="18" place="-1" resultid="110247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99831" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109866" />
                    <RANKING order="2" place="2" resultid="109033" />
                    <RANKING order="3" place="3" resultid="108419" />
                    <RANKING order="4" place="4" resultid="108973" />
                    <RANKING order="5" place="5" resultid="110122" />
                    <RANKING order="6" place="6" resultid="107967" />
                    <RANKING order="7" place="7" resultid="107745" />
                    <RANKING order="8" place="8" resultid="110156" />
                    <RANKING order="9" place="9" resultid="107050" />
                    <RANKING order="10" place="10" resultid="110396" />
                    <RANKING order="11" place="11" resultid="108661" />
                    <RANKING order="12" place="-1" resultid="110187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99832" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110258" />
                    <RANKING order="2" place="2" resultid="107737" />
                    <RANKING order="3" place="3" resultid="110272" />
                    <RANKING order="4" place="4" resultid="106885" />
                    <RANKING order="5" place="5" resultid="107832" />
                    <RANKING order="6" place="6" resultid="109011" />
                    <RANKING order="7" place="7" resultid="108373" />
                    <RANKING order="8" place="8" resultid="109946" />
                    <RANKING order="9" place="9" resultid="107152" />
                    <RANKING order="10" place="-1" resultid="106951" />
                    <RANKING order="11" place="-1" resultid="110165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99833" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109401" />
                    <RANKING order="2" place="2" resultid="109061" />
                    <RANKING order="3" place="3" resultid="109516" />
                    <RANKING order="4" place="4" resultid="106856" />
                    <RANKING order="5" place="5" resultid="106873" />
                    <RANKING order="6" place="6" resultid="109569" />
                    <RANKING order="7" place="7" resultid="108183" />
                    <RANKING order="8" place="8" resultid="110087" />
                    <RANKING order="9" place="-1" resultid="110484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99834" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107027" />
                    <RANKING order="2" place="2" resultid="107008" />
                    <RANKING order="3" place="3" resultid="108353" />
                    <RANKING order="4" place="4" resultid="109857" />
                    <RANKING order="5" place="5" resultid="108242" />
                    <RANKING order="6" place="-1" resultid="106826" />
                    <RANKING order="7" place="-1" resultid="109365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99835" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109409" />
                    <RANKING order="2" place="2" resultid="107129" />
                    <RANKING order="3" place="3" resultid="107498" />
                    <RANKING order="4" place="4" resultid="107492" />
                    <RANKING order="5" place="5" resultid="110070" />
                    <RANKING order="6" place="6" resultid="110451" />
                    <RANKING order="7" place="-1" resultid="107973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99836" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109373" />
                    <RANKING order="2" place="2" resultid="106706" />
                    <RANKING order="3" place="3" resultid="108032" />
                    <RANKING order="4" place="4" resultid="110150" />
                    <RANKING order="5" place="5" resultid="108166" />
                    <RANKING order="6" place="-1" resultid="108363" />
                    <RANKING order="7" place="-1" resultid="107791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99837" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107774" />
                    <RANKING order="2" place="2" resultid="110519" />
                    <RANKING order="3" place="3" resultid="108586" />
                    <RANKING order="4" place="-1" resultid="107782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99838" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108482" />
                    <RANKING order="2" place="-1" resultid="109347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99839" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99840" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99841" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110696" daytime="11:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110697" daytime="11:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110698" daytime="11:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110699" daytime="11:37" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110700" daytime="11:39" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110701" daytime="11:42" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110702" daytime="11:44" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110703" daytime="11:46" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110704" daytime="11:48" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="110705" daytime="11:50" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="110706" daytime="11:52" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99036" daytime="12:31" gender="F" number="20" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99512" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="99513" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110314" />
                    <RANKING order="2" place="2" resultid="107270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99514" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110002" />
                    <RANKING order="2" place="2" resultid="107882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99515" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106891" />
                    <RANKING order="2" place="2" resultid="108103" />
                    <RANKING order="3" place="3" resultid="110201" />
                    <RANKING order="4" place="4" resultid="110003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99516" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108599" />
                    <RANKING order="2" place="2" resultid="106904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99517" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106729" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99518" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110714" daytime="12:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110715" daytime="12:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98924" daytime="09:12" gender="M" number="11" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99767" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110553" />
                    <RANKING order="2" place="2" resultid="110415" />
                    <RANKING order="3" place="3" resultid="109902" />
                    <RANKING order="4" place="4" resultid="109312" />
                    <RANKING order="5" place="5" resultid="110433" />
                    <RANKING order="6" place="6" resultid="108691" />
                    <RANKING order="7" place="-1" resultid="108947" />
                    <RANKING order="8" place="-1" resultid="110509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99768" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106654" />
                    <RANKING order="2" place="2" resultid="107170" />
                    <RANKING order="3" place="3" resultid="107189" />
                    <RANKING order="4" place="4" resultid="106659" />
                    <RANKING order="5" place="5" resultid="107878" />
                    <RANKING order="6" place="6" resultid="107678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99769" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107416" />
                    <RANKING order="2" place="2" resultid="110468" />
                    <RANKING order="3" place="3" resultid="109574" />
                    <RANKING order="4" place="4" resultid="107399" />
                    <RANKING order="5" place="5" resultid="107118" />
                    <RANKING order="6" place="6" resultid="107563" />
                    <RANKING order="7" place="7" resultid="107255" />
                    <RANKING order="8" place="8" resultid="110421" />
                    <RANKING order="9" place="9" resultid="107503" />
                    <RANKING order="10" place="10" resultid="110459" />
                    <RANKING order="11" place="11" resultid="109355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99770" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107234" />
                    <RANKING order="2" place="2" resultid="107725" />
                    <RANKING order="3" place="3" resultid="109055" />
                    <RANKING order="4" place="4" resultid="109562" />
                    <RANKING order="5" place="5" resultid="108050" />
                    <RANKING order="6" place="6" resultid="108057" />
                    <RANKING order="7" place="7" resultid="109608" />
                    <RANKING order="8" place="8" resultid="106600" />
                    <RANKING order="9" place="9" resultid="109934" />
                    <RANKING order="10" place="10" resultid="107696" />
                    <RANKING order="11" place="11" resultid="107626" />
                    <RANKING order="12" place="12" resultid="107616" />
                    <RANKING order="13" place="13" resultid="107950" />
                    <RANKING order="14" place="-1" resultid="110246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99771" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108400" />
                    <RANKING order="2" place="2" resultid="107966" />
                    <RANKING order="3" place="3" resultid="110121" />
                    <RANKING order="4" place="4" resultid="107548" />
                    <RANKING order="5" place="5" resultid="108990" />
                    <RANKING order="6" place="6" resultid="108559" />
                    <RANKING order="7" place="7" resultid="108554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99772" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107736" />
                    <RANKING order="2" place="2" resultid="106884" />
                    <RANKING order="3" place="3" resultid="107831" />
                    <RANKING order="4" place="4" resultid="110164" />
                    <RANKING order="5" place="5" resultid="109170" />
                    <RANKING order="6" place="6" resultid="109945" />
                    <RANKING order="7" place="7" resultid="108424" />
                    <RANKING order="8" place="8" resultid="109010" />
                    <RANKING order="9" place="9" resultid="107687" />
                    <RANKING order="10" place="10" resultid="107151" />
                    <RANKING order="11" place="11" resultid="107136" />
                    <RANKING order="12" place="-1" resultid="106950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99773" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109400" />
                    <RANKING order="2" place="2" resultid="109060" />
                    <RANKING order="3" place="3" resultid="109515" />
                    <RANKING order="4" place="4" resultid="106852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99774" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107026" />
                    <RANKING order="2" place="2" resultid="109847" />
                    <RANKING order="3" place="3" resultid="108023" />
                    <RANKING order="4" place="4" resultid="108442" />
                    <RANKING order="5" place="5" resultid="106825" />
                    <RANKING order="6" place="6" resultid="109392" />
                    <RANKING order="7" place="-1" resultid="108227" />
                    <RANKING order="8" place="-1" resultid="108241" />
                    <RANKING order="9" place="-1" resultid="110490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99775" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110450" />
                    <RANKING order="2" place="2" resultid="107763" />
                    <RANKING order="3" place="3" resultid="110069" />
                    <RANKING order="4" place="4" resultid="108156" />
                    <RANKING order="5" place="5" resultid="108576" />
                    <RANKING order="6" place="-1" resultid="106820" />
                    <RANKING order="7" place="-1" resultid="108254" />
                    <RANKING order="8" place="-1" resultid="108259" />
                    <RANKING order="9" place="-1" resultid="110501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99776" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109372" />
                    <RANKING order="2" place="2" resultid="109379" />
                    <RANKING order="3" place="3" resultid="106722" />
                    <RANKING order="4" place="4" resultid="110063" />
                    <RANKING order="5" place="5" resultid="106717" />
                    <RANKING order="6" place="6" resultid="109469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99777" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110056" />
                    <RANKING order="2" place="2" resultid="109415" />
                    <RANKING order="3" place="3" resultid="110518" />
                    <RANKING order="4" place="4" resultid="107458" />
                    <RANKING order="5" place="5" resultid="107144" />
                    <RANKING order="6" place="6" resultid="108520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99778" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108481" />
                    <RANKING order="2" place="2" resultid="108173" />
                    <RANKING order="3" place="3" resultid="107449" />
                    <RANKING order="4" place="4" resultid="107070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99779" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108487" />
                    <RANKING order="2" place="2" resultid="107822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99780" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99781" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110651" daytime="09:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110652" daytime="09:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110653" daytime="09:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110654" daytime="09:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110655" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110656" daytime="09:21" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110657" daytime="09:23" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110658" daytime="09:24" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110659" daytime="09:26" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="110660" daytime="09:27" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="106294" daytime="09:00" gender="F" number="10" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="106295" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108638" />
                    <RANKING order="2" place="2" resultid="108674" />
                    <RANKING order="3" place="3" resultid="107371" />
                    <RANKING order="4" place="-1" resultid="110441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106296" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106799" />
                    <RANKING order="2" place="2" resultid="106666" />
                    <RANKING order="3" place="3" resultid="107209" />
                    <RANKING order="4" place="4" resultid="107911" />
                    <RANKING order="5" place="5" resultid="110278" />
                    <RANKING order="6" place="6" resultid="109422" />
                    <RANKING order="7" place="-1" resultid="110285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106297" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107227" />
                    <RANKING order="2" place="-1" resultid="107219" />
                    <RANKING order="3" place="-1" resultid="107837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106298" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109928" />
                    <RANKING order="2" place="2" resultid="110180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106299" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108085" />
                    <RANKING order="2" place="2" resultid="107916" />
                    <RANKING order="3" place="3" resultid="108548" />
                    <RANKING order="4" place="4" resultid="109838" />
                    <RANKING order="5" place="5" resultid="107465" />
                    <RANKING order="6" place="6" resultid="110129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106300" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108565" />
                    <RANKING order="2" place="2" resultid="106780" />
                    <RANKING order="3" place="3" resultid="107861" />
                    <RANKING order="4" place="4" resultid="109914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106301" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108496" />
                    <RANKING order="2" place="2" resultid="108014" />
                    <RANKING order="3" place="3" resultid="107988" />
                    <RANKING order="4" place="4" resultid="108380" />
                    <RANKING order="5" place="5" resultid="109507" />
                    <RANKING order="6" place="-1" resultid="106766" />
                    <RANKING order="7" place="-1" resultid="106759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106302" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108348" />
                    <RANKING order="2" place="2" resultid="110222" />
                    <RANKING order="3" place="3" resultid="108455" />
                    <RANKING order="4" place="4" resultid="106959" />
                    <RANKING order="5" place="-1" resultid="108389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106303" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108063" />
                    <RANKING order="2" place="2" resultid="108461" />
                    <RANKING order="3" place="3" resultid="107904" />
                    <RANKING order="4" place="4" resultid="107470" />
                    <RANKING order="5" place="5" resultid="110355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106304" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109453" />
                    <RANKING order="2" place="2" resultid="110095" />
                    <RANKING order="3" place="3" resultid="107081" />
                    <RANKING order="4" place="4" resultid="106697" />
                    <RANKING order="5" place="5" resultid="108469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106305" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106306" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107014" />
                    <RANKING order="2" place="2" resultid="107799" />
                    <RANKING order="3" place="3" resultid="109131" />
                    <RANKING order="4" place="4" resultid="107813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106307" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="106308" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="106309" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110645" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110646" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110647" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110648" daytime="09:07" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110649" daytime="09:09" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110650" daytime="09:10" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98972" daytime="11:11" gender="F" number="16" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99812" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107942" />
                    <RANKING order="2" place="2" resultid="108639" />
                    <RANKING order="3" place="3" resultid="108675" />
                    <RANKING order="4" place="4" resultid="110404" />
                    <RANKING order="5" place="5" resultid="110375" />
                    <RANKING order="6" place="6" resultid="109896" />
                    <RANKING order="7" place="7" resultid="107123" />
                    <RANKING order="8" place="-1" resultid="108957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99813" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108218" />
                    <RANKING order="2" place="2" resultid="107210" />
                    <RANKING order="3" place="3" resultid="109423" />
                    <RANKING order="4" place="-1" resultid="110567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99814" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107484" />
                    <RANKING order="2" place="2" resultid="108623" />
                    <RANKING order="3" place="3" resultid="107872" />
                    <RANKING order="4" place="4" resultid="107838" />
                    <RANKING order="5" place="5" resultid="107033" />
                    <RANKING order="6" place="-1" resultid="110310" />
                    <RANKING order="7" place="-1" resultid="107220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99815" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107707" />
                    <RANKING order="2" place="2" resultid="107715" />
                    <RANKING order="3" place="3" resultid="108683" />
                    <RANKING order="4" place="4" resultid="109018" />
                    <RANKING order="5" place="5" resultid="109929" />
                    <RANKING order="6" place="6" resultid="108965" />
                    <RANKING order="7" place="7" resultid="106792" />
                    <RANKING order="8" place="8" resultid="106595" />
                    <RANKING order="9" place="-1" resultid="110305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99816" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108086" />
                    <RANKING order="2" place="2" resultid="106983" />
                    <RANKING order="3" place="3" resultid="106426" />
                    <RANKING order="4" place="4" resultid="108549" />
                    <RANKING order="5" place="5" resultid="107466" />
                    <RANKING order="6" place="-1" resultid="110136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99817" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108079" />
                    <RANKING order="2" place="2" resultid="108434" />
                    <RANKING order="3" place="3" resultid="107856" />
                    <RANKING order="4" place="4" resultid="107042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99818" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108497" />
                    <RANKING order="2" place="2" resultid="108526" />
                    <RANKING order="3" place="3" resultid="108042" />
                    <RANKING order="4" place="4" resultid="110104" />
                    <RANKING order="5" place="5" resultid="106767" />
                    <RANKING order="6" place="-1" resultid="106760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99819" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109529" />
                    <RANKING order="2" place="2" resultid="110353" />
                    <RANKING order="3" place="3" resultid="110173" />
                    <RANKING order="4" place="-1" resultid="108390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99820" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108064" />
                    <RANKING order="2" place="2" resultid="107084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99821" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108093" />
                    <RANKING order="2" place="2" resultid="108470" />
                    <RANKING order="3" place="3" resultid="110583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99822" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99823" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107015" />
                    <RANKING order="2" place="2" resultid="109132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99824" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99825" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99826" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110690" daytime="11:11" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110691" daytime="11:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110692" daytime="11:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110693" daytime="11:21" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110694" daytime="11:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110695" daytime="11:26" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="106277" daytime="10:35" gender="M" number="15" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="106278" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107112" />
                    <RANKING order="2" place="2" resultid="109536" />
                    <RANKING order="3" place="3" resultid="107105" />
                    <RANKING order="4" place="4" resultid="109213" />
                    <RANKING order="5" place="5" resultid="106673" />
                    <RANKING order="6" place="6" resultid="107924" />
                    <RANKING order="7" place="7" resultid="108703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106279" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107721" />
                    <RANKING order="2" place="2" resultid="109475" />
                    <RANKING order="3" place="3" resultid="110382" />
                    <RANKING order="4" place="4" resultid="107630" />
                    <RANKING order="5" place="5" resultid="107849" />
                    <RANKING order="6" place="6" resultid="108697" />
                    <RANKING order="7" place="7" resultid="110579" />
                    <RANKING order="8" place="8" resultid="106606" />
                    <RANKING order="9" place="9" resultid="107679" />
                    <RANKING order="10" place="-1" resultid="106649" />
                    <RANKING order="11" place="-1" resultid="107247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106280" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108651" />
                    <RANKING order="2" place="2" resultid="107392" />
                    <RANKING order="3" place="3" resultid="107400" />
                    <RANKING order="4" place="4" resultid="108571" />
                    <RANKING order="5" place="5" resultid="107407" />
                    <RANKING order="6" place="6" resultid="108630" />
                    <RANKING order="7" place="7" resultid="107504" />
                    <RANKING order="8" place="8" resultid="109833" />
                    <RANKING order="9" place="9" resultid="110422" />
                    <RANKING order="10" place="10" resultid="110460" />
                    <RANKING order="11" place="11" resultid="106639" />
                    <RANKING order="12" place="12" resultid="107476" />
                    <RANKING order="13" place="-1" resultid="107620" />
                    <RANKING order="14" place="-1" resultid="108711" />
                    <RANKING order="15" place="-1" resultid="109820" />
                    <RANKING order="16" place="-1" resultid="107022" />
                    <RANKING order="17" place="-1" resultid="109459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106281" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107665" />
                    <RANKING order="2" place="2" resultid="109441" />
                    <RANKING order="3" place="3" resultid="107726" />
                    <RANKING order="4" place="4" resultid="106580" />
                    <RANKING order="5" place="5" resultid="107434" />
                    <RANKING order="6" place="6" resultid="107555" />
                    <RANKING order="7" place="7" resultid="107571" />
                    <RANKING order="8" place="8" resultid="109149" />
                    <RANKING order="9" place="9" resultid="109935" />
                    <RANKING order="10" place="10" resultid="109385" />
                    <RANKING order="11" place="11" resultid="107697" />
                    <RANKING order="12" place="12" resultid="107599" />
                    <RANKING order="13" place="13" resultid="106633" />
                    <RANKING order="14" place="14" resultid="107617" />
                    <RANKING order="15" place="15" resultid="108592" />
                    <RANKING order="16" place="-1" resultid="106890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106282" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109865" />
                    <RANKING order="2" place="2" resultid="109032" />
                    <RANKING order="3" place="3" resultid="108972" />
                    <RANKING order="4" place="4" resultid="108401" />
                    <RANKING order="5" place="5" resultid="107844" />
                    <RANKING order="6" place="6" resultid="107744" />
                    <RANKING order="7" place="7" resultid="109464" />
                    <RANKING order="8" place="8" resultid="108982" />
                    <RANKING order="9" place="9" resultid="109883" />
                    <RANKING order="10" place="10" resultid="108997" />
                    <RANKING order="11" place="11" resultid="110193" />
                    <RANKING order="12" place="12" resultid="108660" />
                    <RANKING order="13" place="13" resultid="109960" />
                    <RANKING order="14" place="-1" resultid="110395" />
                    <RANKING order="15" place="-1" resultid="107252" />
                    <RANKING order="16" place="-1" resultid="108991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106283" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110271" />
                    <RANKING order="2" place="2" resultid="110257" />
                    <RANKING order="3" place="3" resultid="107933" />
                    <RANKING order="4" place="4" resultid="108372" />
                    <RANKING order="5" place="5" resultid="106878" />
                    <RANKING order="6" place="6" resultid="107688" />
                    <RANKING order="7" place="7" resultid="107867" />
                    <RANKING order="8" place="8" resultid="107137" />
                    <RANKING order="9" place="-1" resultid="110427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106284" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109581" />
                    <RANKING order="2" place="2" resultid="110483" />
                    <RANKING order="3" place="3" resultid="107077" />
                    <RANKING order="4" place="4" resultid="106865" />
                    <RANKING order="5" place="5" resultid="106999" />
                    <RANKING order="6" place="6" resultid="106612" />
                    <RANKING order="7" place="7" resultid="109166" />
                    <RANKING order="8" place="8" resultid="108182" />
                    <RANKING order="9" place="9" resultid="108920" />
                    <RANKING order="10" place="10" resultid="110409" />
                    <RANKING order="11" place="-1" resultid="110253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106285" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109974" />
                    <RANKING order="2" place="2" resultid="108443" />
                    <RANKING order="3" place="3" resultid="108024" />
                    <RANKING order="4" place="4" resultid="108208" />
                    <RANKING order="5" place="5" resultid="110491" />
                    <RANKING order="6" place="6" resultid="109393" />
                    <RANKING order="7" place="7" resultid="106832" />
                    <RANKING order="8" place="-1" resultid="108228" />
                    <RANKING order="9" place="-1" resultid="109364" />
                    <RANKING order="10" place="-1" resultid="106838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106286" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109408" />
                    <RANKING order="2" place="2" resultid="110540" />
                    <RANKING order="3" place="3" resultid="107764" />
                    <RANKING order="4" place="4" resultid="110526" />
                    <RANKING order="5" place="5" resultid="108071" />
                    <RANKING order="6" place="6" resultid="108260" />
                    <RANKING order="7" place="7" resultid="108255" />
                    <RANKING order="8" place="8" resultid="108577" />
                    <RANKING order="9" place="-1" resultid="110502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106287" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106406" />
                    <RANKING order="2" place="2" resultid="109380" />
                    <RANKING order="3" place="3" resultid="106938" />
                    <RANKING order="4" place="4" resultid="108532" />
                    <RANKING order="5" place="5" resultid="106808" />
                    <RANKING order="6" place="6" resultid="107790" />
                    <RANKING order="7" place="7" resultid="109470" />
                    <RANKING order="8" place="8" resultid="106815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106288" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110057" />
                    <RANKING order="2" place="2" resultid="109416" />
                    <RANKING order="3" place="3" resultid="108585" />
                    <RANKING order="4" place="-1" resultid="108521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106289" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106688" />
                    <RANKING order="2" place="2" resultid="106349" />
                    <RANKING order="3" place="3" resultid="108513" />
                    <RANKING order="4" place="4" resultid="107071" />
                    <RANKING order="5" place="-1" resultid="107450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106290" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="106291" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="106292" agemax="94" agemin="90" name="KAT.N, 90-94 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="108005" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110677" daytime="10:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110678" daytime="10:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110679" daytime="10:47" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110680" daytime="10:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110681" daytime="10:53" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110682" daytime="10:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110683" daytime="10:57" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110684" daytime="10:59" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110685" daytime="11:01" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="110686" daytime="11:03" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="110687" daytime="11:05" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="110688" daytime="11:07" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="110689" daytime="11:09" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98940" daytime="09:29" gender="F" number="12" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99782" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108956" />
                    <RANKING order="2" place="2" resultid="109895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99783" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107673" />
                    <RANKING order="2" place="2" resultid="108217" />
                    <RANKING order="3" place="3" resultid="108645" />
                    <RANKING order="4" place="4" resultid="109988" />
                    <RANKING order="5" place="5" resultid="107379" />
                    <RANKING order="6" place="-1" resultid="110566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99784" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107483" />
                    <RANKING order="2" place="2" resultid="107871" />
                    <RANKING order="3" place="3" resultid="106988" />
                    <RANKING order="4" place="4" resultid="107387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99785" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106785" />
                    <RANKING order="2" place="2" resultid="107714" />
                    <RANKING order="3" place="3" resultid="109017" />
                    <RANKING order="4" place="4" resultid="106791" />
                    <RANKING order="5" place="5" resultid="110238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99786" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99787" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107855" />
                    <RANKING order="2" place="2" resultid="108433" />
                    <RANKING order="3" place="3" resultid="109824" />
                    <RANKING order="4" place="4" resultid="107041" />
                    <RANKING order="5" place="5" resultid="107862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99788" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109446" />
                    <RANKING order="2" place="2" resultid="110103" />
                    <RANKING order="3" place="3" resultid="108381" />
                    <RANKING order="4" place="4" resultid="109545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99789" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109528" />
                    <RANKING order="2" place="2" resultid="109176" />
                    <RANKING order="3" place="3" resultid="106422" />
                    <RANKING order="4" place="4" resultid="110172" />
                    <RANKING order="5" place="5" resultid="110230" />
                    <RANKING order="6" place="-1" resultid="108386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99790" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109908" />
                    <RANKING order="2" place="2" resultid="110356" />
                    <RANKING order="3" place="-1" resultid="106748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99791" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99792" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99793" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99794" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99795" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99796" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110661" daytime="09:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110662" daytime="09:37" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110663" daytime="09:41" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110664" daytime="09:46" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99059" daytime="12:39" gender="M" number="21" order="13" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99519" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="108722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99520" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107267" />
                    <RANKING order="2" place="2" resultid="106679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99521" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107268" />
                    <RANKING order="2" place="2" resultid="107424" />
                    <RANKING order="3" place="3" resultid="109586" />
                    <RANKING order="4" place="4" resultid="109038" />
                    <RANKING order="5" place="5" resultid="107632" />
                    <RANKING order="6" place="6" resultid="110194" />
                    <RANKING order="7" place="7" resultid="106622" />
                    <RANKING order="8" place="8" resultid="109482" />
                    <RANKING order="9" place="9" resultid="108720" />
                    <RANKING order="10" place="10" resultid="107633" />
                    <RANKING order="11" place="11" resultid="110004" />
                    <RANKING order="12" place="-1" resultid="108603" />
                    <RANKING order="13" place="-1" resultid="107634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99522" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108448" />
                    <RANKING order="2" place="2" resultid="110315" />
                    <RANKING order="3" place="3" resultid="110005" />
                    <RANKING order="4" place="4" resultid="107884" />
                    <RANKING order="5" place="5" resultid="107525" />
                    <RANKING order="6" place="6" resultid="107055" />
                    <RANKING order="7" place="-1" resultid="109039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99523" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108105" />
                    <RANKING order="2" place="2" resultid="106896" />
                    <RANKING order="3" place="3" resultid="109587" />
                    <RANKING order="4" place="4" resultid="110006" />
                    <RANKING order="5" place="5" resultid="110111" />
                    <RANKING order="6" place="6" resultid="107157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99524" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109481" />
                    <RANKING order="2" place="2" resultid="106895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99525" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106726" />
                    <RANKING order="2" place="2" resultid="107521" />
                    <RANKING order="3" place="-1" resultid="108595" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110716" daytime="12:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110717" daytime="12:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110718" daytime="12:47" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110719" daytime="12:50" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-10-22" daytime="16:00" endtime="20:21" number="3" warmupfrom="15:00" warmupuntil="15:50">
          <EVENTS>
            <EVENT eventid="99314" daytime="17:16" gender="F" number="26" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99872" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108640" />
                    <RANKING order="2" place="2" resultid="108676" />
                    <RANKING order="3" place="-1" resultid="110444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99873" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108220" />
                    <RANKING order="2" place="2" resultid="110280" />
                    <RANKING order="3" place="3" resultid="107912" />
                    <RANKING order="4" place="4" resultid="109425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99874" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107229" />
                    <RANKING order="2" place="2" resultid="109876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99875" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108684" />
                    <RANKING order="2" place="2" resultid="109930" />
                    <RANKING order="3" place="3" resultid="110182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99876" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108088" />
                    <RANKING order="2" place="2" resultid="106984" />
                    <RANKING order="3" place="3" resultid="107918" />
                    <RANKING order="4" place="4" resultid="109839" />
                    <RANKING order="5" place="5" resultid="107467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99877" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106782" />
                    <RANKING order="2" place="2" resultid="109916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99878" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108499" />
                    <RANKING order="2" place="2" resultid="107990" />
                    <RANKING order="3" place="3" resultid="108017" />
                    <RANKING order="4" place="4" resultid="108382" />
                    <RANKING order="5" place="5" resultid="109547" />
                    <RANKING order="6" place="-1" resultid="109509" />
                    <RANKING order="7" place="-1" resultid="106761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99879" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107091" />
                    <RANKING order="2" place="2" resultid="108349" />
                    <RANKING order="3" place="3" resultid="110224" />
                    <RANKING order="4" place="4" resultid="108457" />
                    <RANKING order="5" place="-1" resultid="108391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99880" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108464" />
                    <RANKING order="2" place="2" resultid="107907" />
                    <RANKING order="3" place="3" resultid="107472" />
                    <RANKING order="4" place="4" resultid="110358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99881" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109455" />
                    <RANKING order="2" place="2" resultid="108472" />
                    <RANKING order="3" place="3" resultid="110475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99882" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99883" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107017" />
                    <RANKING order="2" place="2" resultid="109134" />
                    <RANKING order="3" place="3" resultid="107801" />
                    <RANKING order="4" place="4" resultid="107815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99884" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99885" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99886" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110752" daytime="17:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110753" daytime="17:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110754" daytime="17:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110755" daytime="17:27" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110756" daytime="17:30" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99282" daytime="19:39" gender="M" number="33" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99947" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109539" />
                    <RANKING order="2" place="2" resultid="109905" />
                    <RANKING order="3" place="3" resultid="110436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99948" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107173" />
                    <RANKING order="2" place="2" resultid="110292" />
                    <RANKING order="3" place="-1" resultid="106401" />
                    <RANKING order="4" place="-1" resultid="109478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99949" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106978" />
                    <RANKING order="2" place="2" resultid="109577" />
                    <RANKING order="3" place="3" resultid="108654" />
                    <RANKING order="4" place="4" resultid="109969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99950" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109557" />
                    <RANKING order="2" place="2" resultid="109956" />
                    <RANKING order="3" place="-1" resultid="106970" />
                    <RANKING order="4" place="-1" resultid="108412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99951" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109868" />
                    <RANKING order="2" place="2" resultid="110158" />
                    <RANKING order="3" place="3" resultid="110575" />
                    <RANKING order="4" place="-1" resultid="107051" />
                    <RANKING order="5" place="-1" resultid="109000" />
                    <RANKING order="6" place="-1" resultid="109341" />
                    <RANKING order="7" place="-1" resultid="110189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99952" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109027" />
                    <RANKING order="2" place="2" resultid="110274" />
                    <RANKING order="3" place="3" resultid="109173" />
                    <RANKING order="4" place="4" resultid="107757" />
                    <RANKING order="5" place="5" resultid="109948" />
                    <RANKING order="6" place="6" resultid="107690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99953" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109063" />
                    <RANKING order="2" place="2" resultid="110266" />
                    <RANKING order="3" place="3" resultid="109167" />
                    <RANKING order="4" place="4" resultid="106848" />
                    <RANKING order="5" place="-1" resultid="106615" />
                    <RANKING order="6" place="-1" resultid="108185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99954" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108445" />
                    <RANKING order="2" place="2" resultid="109859" />
                    <RANKING order="3" place="3" resultid="109322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99955" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110072" />
                    <RANKING order="2" place="2" resultid="107131" />
                    <RANKING order="3" place="3" resultid="108159" />
                    <RANKING order="4" place="4" resultid="110453" />
                    <RANKING order="5" place="5" resultid="108074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99956" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106939" />
                    <RANKING order="2" place="2" resultid="108535" />
                    <RANKING order="3" place="3" resultid="108168" />
                    <RANKING order="4" place="4" resultid="107444" />
                    <RANKING order="5" place="-1" resultid="108365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99957" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="107784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99958" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99959" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99960" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99961" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110788" daytime="19:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110789" daytime="19:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110790" daytime="19:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110791" daytime="20:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110792" daytime="20:12" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99091" daytime="16:21" gender="M" number="23" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99124" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110534" />
                    <RANKING order="2" place="2" resultid="110555" />
                    <RANKING order="3" place="3" resultid="107925" />
                    <RANKING order="4" place="4" resultid="108949" />
                    <RANKING order="5" place="5" resultid="110561" />
                    <RANKING order="6" place="-1" resultid="110511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99125" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107177" />
                    <RANKING order="2" place="2" resultid="109005" />
                    <RANKING order="3" place="3" resultid="110291" />
                    <RANKING order="4" place="4" resultid="110388" />
                    <RANKING order="5" place="5" resultid="107850" />
                    <RANKING order="6" place="6" resultid="107879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99126" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107243" />
                    <RANKING order="2" place="2" resultid="107394" />
                    <RANKING order="3" place="3" resultid="107511" />
                    <RANKING order="4" place="4" resultid="107257" />
                    <RANKING order="5" place="5" resultid="107611" />
                    <RANKING order="6" place="6" resultid="109968" />
                    <RANKING order="7" place="7" resultid="107565" />
                    <RANKING order="8" place="8" resultid="108631" />
                    <RANKING order="9" place="9" resultid="107478" />
                    <RANKING order="10" place="-1" resultid="110858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99127" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109955" />
                    <RANKING order="2" place="2" resultid="109610" />
                    <RANKING order="3" place="3" resultid="108411" />
                    <RANKING order="4" place="4" resultid="107593" />
                    <RANKING order="5" place="5" resultid="109076" />
                    <RANKING order="6" place="6" resultid="107584" />
                    <RANKING order="7" place="7" resultid="108593" />
                    <RANKING order="8" place="8" resultid="107952" />
                    <RANKING order="9" place="-1" resultid="107577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99128" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108420" />
                    <RANKING order="2" place="2" resultid="107968" />
                    <RANKING order="3" place="3" resultid="108984" />
                    <RANKING order="4" place="4" resultid="108561" />
                    <RANKING order="5" place="5" resultid="107746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99129" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109026" />
                    <RANKING order="2" place="2" resultid="107934" />
                    <RANKING order="3" place="3" resultid="109012" />
                    <RANKING order="4" place="4" resultid="108374" />
                    <RANKING order="5" place="5" resultid="107756" />
                    <RANKING order="6" place="6" resultid="107153" />
                    <RANKING order="7" place="7" resultid="110428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99130" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106866" />
                    <RANKING order="2" place="2" resultid="106857" />
                    <RANKING order="3" place="3" resultid="110088" />
                    <RANKING order="4" place="4" resultid="109570" />
                    <RANKING order="5" place="5" resultid="106847" />
                    <RANKING order="6" place="6" resultid="106874" />
                    <RANKING order="7" place="7" resultid="109436" />
                    <RANKING order="8" place="8" resultid="110410" />
                    <RANKING order="9" place="-1" resultid="110265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99131" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107009" />
                    <RANKING order="2" place="2" resultid="108354" />
                    <RANKING order="3" place="3" resultid="110080" />
                    <RANKING order="4" place="4" resultid="110862" />
                    <RANKING order="5" place="5" resultid="106827" />
                    <RANKING order="6" place="6" resultid="108229" />
                    <RANKING order="7" place="-1" resultid="109366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99132" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107130" />
                    <RANKING order="2" place="2" resultid="108476" />
                    <RANKING order="3" place="3" resultid="108203" />
                    <RANKING order="4" place="4" resultid="107499" />
                    <RANKING order="5" place="5" resultid="107765" />
                    <RANKING order="6" place="6" resultid="108261" />
                    <RANKING order="7" place="7" resultid="108256" />
                    <RANKING order="8" place="8" resultid="108578" />
                    <RANKING order="9" place="-1" resultid="106821" />
                    <RANKING order="10" place="-1" resultid="108236" />
                    <RANKING order="11" place="-1" resultid="107974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99133" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108010" />
                    <RANKING order="2" place="2" resultid="109815" />
                    <RANKING order="3" place="3" resultid="110151" />
                    <RANKING order="4" place="4" resultid="108167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99134" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107775" />
                    <RANKING order="2" place="2" resultid="107145" />
                    <RANKING order="3" place="3" resultid="107460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99135" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107998" />
                    <RANKING order="2" place="2" resultid="108483" />
                    <RANKING order="3" place="3" resultid="108514" />
                    <RANKING order="4" place="4" resultid="107072" />
                    <RANKING order="5" place="-1" resultid="109348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99136" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99137" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99138" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110726" daytime="16:21" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110727" daytime="16:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110728" daytime="16:29" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110729" daytime="16:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110730" daytime="16:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110731" daytime="16:37" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110732" daytime="16:39" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110733" daytime="16:42" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110734" daytime="16:44" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99266" daytime="19:12" gender="F" number="32" order="13" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99932" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108677" />
                    <RANKING order="2" place="-1" resultid="109898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99933" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109991" />
                    <RANKING order="2" place="2" resultid="108906" />
                    <RANKING order="3" place="3" resultid="110569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99934" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107486" />
                    <RANKING order="2" place="2" resultid="108626" />
                    <RANKING order="3" place="3" resultid="107388" />
                    <RANKING order="4" place="4" resultid="107874" />
                    <RANKING order="5" place="5" resultid="107840" />
                    <RANKING order="6" place="6" resultid="107035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99935" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108271" />
                    <RANKING order="2" place="2" resultid="106597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99936" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106427" />
                    <RANKING order="2" place="2" resultid="110139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99937" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109827" />
                    <RANKING order="2" place="2" resultid="107044" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99938" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108925" />
                    <RANKING order="2" place="2" resultid="108527" />
                    <RANKING order="3" place="3" resultid="109548" />
                    <RANKING order="4" place="-1" resultid="106762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99939" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107092" />
                    <RANKING order="2" place="2" resultid="110175" />
                    <RANKING order="3" place="3" resultid="110233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99940" agemax="64" agemin="60" name="KAT.H, 60-64 lat" />
                <AGEGROUP agegroupid="99941" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99942" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99943" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99944" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99945" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99946" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110785" daytime="19:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110786" daytime="19:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110787" daytime="19:31" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99154" daytime="16:46" gender="F" number="24" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99842" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107373" />
                    <RANKING order="2" place="2" resultid="110376" />
                    <RANKING order="3" place="3" resultid="109897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99843" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106801" />
                    <RANKING order="2" place="2" resultid="106669" />
                    <RANKING order="3" place="3" resultid="109990" />
                    <RANKING order="4" place="4" resultid="109424" />
                    <RANKING order="5" place="-1" resultid="107204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99844" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106588" />
                    <RANKING order="2" place="2" resultid="110299" />
                    <RANKING order="3" place="3" resultid="106990" />
                    <RANKING order="4" place="4" resultid="108625" />
                    <RANKING order="5" place="5" resultid="110312" />
                    <RANKING order="6" place="6" resultid="106619" />
                    <RANKING order="7" place="7" resultid="107839" />
                    <RANKING order="8" place="8" resultid="107034" />
                    <RANKING order="9" place="-1" resultid="107221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99845" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108270" />
                    <RANKING order="2" place="2" resultid="107708" />
                    <RANKING order="3" place="3" resultid="106787" />
                    <RANKING order="4" place="4" resultid="107717" />
                    <RANKING order="5" place="5" resultid="108966" />
                    <RANKING order="6" place="6" resultid="109020" />
                    <RANKING order="7" place="7" resultid="110306" />
                    <RANKING order="8" place="8" resultid="106794" />
                    <RANKING order="9" place="-1" resultid="106645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99846" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108087" />
                    <RANKING order="2" place="2" resultid="108550" />
                    <RANKING order="3" place="3" resultid="107067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99847" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108080" />
                    <RANKING order="2" place="2" resultid="108567" />
                    <RANKING order="3" place="3" resultid="107858" />
                    <RANKING order="4" place="4" resultid="108436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99848" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108498" />
                    <RANKING order="2" place="2" resultid="108016" />
                    <RANKING order="3" place="3" resultid="110106" />
                    <RANKING order="4" place="4" resultid="106769" />
                    <RANKING order="5" place="5" resultid="106775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99849" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108506" />
                    <RANKING order="2" place="2" resultid="109531" />
                    <RANKING order="3" place="3" resultid="109179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99850" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108065" />
                    <RANKING order="2" place="2" resultid="107906" />
                    <RANKING order="3" place="3" resultid="108463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99851" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110097" />
                    <RANKING order="2" place="2" resultid="108095" />
                    <RANKING order="3" place="3" resultid="106943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99852" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106695" />
                    <RANKING order="2" place="2" resultid="108544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99853" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107016" />
                    <RANKING order="2" place="2" resultid="109133" />
                    <RANKING order="3" place="3" resultid="107809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99854" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99855" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99856" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110735" daytime="16:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110736" daytime="16:49" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110737" daytime="16:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110738" daytime="16:53" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110739" daytime="16:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110740" daytime="16:56" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99234" daytime="18:52" gender="F" number="30" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99526" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="99527" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107269" />
                    <RANKING order="2" place="2" resultid="110317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99528" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110007" />
                    <RANKING order="2" place="2" resultid="107881" />
                    <RANKING order="3" place="-1" resultid="108719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99529" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106898" />
                    <RANKING order="2" place="2" resultid="108104" />
                    <RANKING order="3" place="3" resultid="110200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99530" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108600" />
                    <RANKING order="2" place="2" resultid="106897" />
                    <RANKING order="3" place="3" resultid="110008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99531" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="99532" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110779" daytime="18:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110780" daytime="18:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99186" daytime="17:32" gender="M" number="27" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99887" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109904" />
                    <RANKING order="2" place="2" resultid="110435" />
                    <RANKING order="3" place="3" resultid="108951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99888" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107172" />
                    <RANKING order="2" place="2" resultid="106662" />
                    <RANKING order="3" place="3" resultid="107680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99889" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107419" />
                    <RANKING order="2" place="2" resultid="110469" />
                    <RANKING order="3" place="3" resultid="109576" />
                    <RANKING order="4" place="4" resultid="107566" />
                    <RANKING order="5" place="5" resultid="107402" />
                    <RANKING order="6" place="6" resultid="110859" />
                    <RANKING order="7" place="7" resultid="110461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99890" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107237" />
                    <RANKING order="2" place="2" resultid="107728" />
                    <RANKING order="3" place="3" resultid="109563" />
                    <RANKING order="4" place="4" resultid="108059" />
                    <RANKING order="5" place="5" resultid="108053" />
                    <RANKING order="6" place="6" resultid="107698" />
                    <RANKING order="7" place="7" resultid="106602" />
                    <RANKING order="8" place="8" resultid="107585" />
                    <RANKING order="9" place="9" resultid="107605" />
                    <RANKING order="10" place="10" resultid="107953" />
                    <RANKING order="11" place="-1" resultid="109936" />
                    <RANKING order="12" place="-1" resultid="110249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99891" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108403" />
                    <RANKING order="2" place="2" resultid="110124" />
                    <RANKING order="3" place="3" resultid="110397" />
                    <RANKING order="4" place="4" resultid="110157" />
                    <RANKING order="5" place="-1" resultid="107969" />
                    <RANKING order="6" place="-1" resultid="109884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99892" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107738" />
                    <RANKING order="2" place="2" resultid="110260" />
                    <RANKING order="3" place="3" resultid="106886" />
                    <RANKING order="4" place="4" resultid="110166" />
                    <RANKING order="5" place="5" resultid="109172" />
                    <RANKING order="6" place="6" resultid="108427" />
                    <RANKING order="7" place="7" resultid="107689" />
                    <RANKING order="8" place="-1" resultid="106953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99893" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109402" />
                    <RANKING order="2" place="2" resultid="109517" />
                    <RANKING order="3" place="3" resultid="107001" />
                    <RANKING order="4" place="-1" resultid="106854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99894" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107028" />
                    <RANKING order="2" place="2" resultid="108444" />
                    <RANKING order="3" place="3" resultid="109975" />
                    <RANKING order="4" place="4" resultid="108355" />
                    <RANKING order="5" place="5" resultid="108230" />
                    <RANKING order="6" place="6" resultid="108244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99895" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109410" />
                    <RANKING order="2" place="2" resultid="110071" />
                    <RANKING order="3" place="3" resultid="110452" />
                    <RANKING order="4" place="4" resultid="108158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99896" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109374" />
                    <RANKING order="2" place="2" resultid="109381" />
                    <RANKING order="3" place="3" resultid="106723" />
                    <RANKING order="4" place="4" resultid="110064" />
                    <RANKING order="5" place="5" resultid="110366" />
                    <RANKING order="6" place="-1" resultid="108035" />
                    <RANKING order="7" place="-1" resultid="108364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99897" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110058" />
                    <RANKING order="2" place="2" resultid="109417" />
                    <RANKING order="3" place="3" resultid="108522" />
                    <RANKING order="4" place="-1" resultid="107146" />
                    <RANKING order="5" place="-1" resultid="107461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99898" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107451" />
                    <RANKING order="2" place="2" resultid="107073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99899" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108489" />
                    <RANKING order="2" place="2" resultid="107824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99900" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99901" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110757" daytime="17:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110758" daytime="17:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110759" daytime="17:39" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110760" daytime="17:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110761" daytime="17:44" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110762" daytime="17:46" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110763" daytime="17:49" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99250" daytime="18:59" gender="M" number="31" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99533" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="108723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99534" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107266" />
                    <RANKING order="2" place="2" resultid="106678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99535" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107265" />
                    <RANKING order="2" place="2" resultid="107425" />
                    <RANKING order="3" place="3" resultid="110009" />
                    <RANKING order="4" place="4" resultid="109588" />
                    <RANKING order="5" place="5" resultid="107635" />
                    <RANKING order="6" place="6" resultid="106623" />
                    <RANKING order="7" place="7" resultid="110195" />
                    <RANKING order="8" place="8" resultid="107636" />
                    <RANKING order="9" place="9" resultid="109483" />
                    <RANKING order="10" place="10" resultid="108721" />
                    <RANKING order="11" place="11" resultid="110010" />
                    <RANKING order="12" place="-1" resultid="107637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99536" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109040" />
                    <RANKING order="2" place="2" resultid="110318" />
                    <RANKING order="3" place="3" resultid="107883" />
                    <RANKING order="4" place="4" resultid="109041" />
                    <RANKING order="5" place="5" resultid="107524" />
                    <RANKING order="6" place="6" resultid="107056" />
                    <RANKING order="7" place="7" resultid="110011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99537" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106900" />
                    <RANKING order="2" place="2" resultid="108106" />
                    <RANKING order="3" place="3" resultid="109589" />
                    <RANKING order="4" place="4" resultid="110112" />
                    <RANKING order="5" place="5" resultid="107158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99538" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109480" />
                    <RANKING order="2" place="2" resultid="106899" />
                    <RANKING order="3" place="3" resultid="110012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99539" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106727" />
                    <RANKING order="2" place="2" resultid="108596" />
                    <RANKING order="3" place="3" resultid="107520" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110781" daytime="18:59" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110782" daytime="19:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110783" daytime="19:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110784" daytime="19:09" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99218" daytime="18:14" gender="M" number="29" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99917" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107545" />
                    <RANKING order="2" place="2" resultid="109538" />
                    <RANKING order="3" place="3" resultid="110556" />
                    <RANKING order="4" place="4" resultid="107108" />
                    <RANKING order="5" place="5" resultid="106674" />
                    <RANKING order="6" place="6" resultid="107926" />
                    <RANKING order="7" place="7" resultid="108705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99918" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109890" />
                    <RANKING order="2" place="2" resultid="110383" />
                    <RANKING order="3" place="3" resultid="106400" />
                    <RANKING order="4" place="4" resultid="107851" />
                    <RANKING order="5" place="5" resultid="110861" />
                    <RANKING order="6" place="6" resultid="106607" />
                    <RANKING order="7" place="7" resultid="107681" />
                    <RANKING order="8" place="-1" resultid="106650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99919" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107244" />
                    <RANKING order="2" place="2" resultid="106977" />
                    <RANKING order="3" place="3" resultid="107512" />
                    <RANKING order="4" place="4" resultid="109523" />
                    <RANKING order="5" place="5" resultid="107410" />
                    <RANKING order="6" place="6" resultid="109358" />
                    <RANKING order="7" place="7" resultid="109835" />
                    <RANKING order="8" place="8" resultid="106640" />
                    <RANKING order="9" place="9" resultid="110462" />
                    <RANKING order="10" place="10" resultid="107506" />
                    <RANKING order="11" place="11" resultid="107479" />
                    <RANKING order="12" place="-1" resultid="107622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99920" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109556" />
                    <RANKING order="2" place="2" resultid="107668" />
                    <RANKING order="3" place="3" resultid="107558" />
                    <RANKING order="4" place="4" resultid="109443" />
                    <RANKING order="5" place="5" resultid="109564" />
                    <RANKING order="6" place="6" resultid="110210" />
                    <RANKING order="7" place="7" resultid="109387" />
                    <RANKING order="8" place="8" resultid="109937" />
                    <RANKING order="9" place="9" resultid="107699" />
                    <RANKING order="10" place="10" resultid="106634" />
                    <RANKING order="11" place="-1" resultid="106583" />
                    <RANKING order="12" place="-1" resultid="107594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99921" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108975" />
                    <RANKING order="2" place="2" resultid="107747" />
                    <RANKING order="3" place="3" resultid="106575" />
                    <RANKING order="4" place="4" resultid="109465" />
                    <RANKING order="5" place="5" resultid="108999" />
                    <RANKING order="6" place="6" resultid="110398" />
                    <RANKING order="7" place="7" resultid="109142" />
                    <RANKING order="8" place="8" resultid="109885" />
                    <RANKING order="9" place="9" resultid="108663" />
                    <RANKING order="10" place="10" resultid="109962" />
                    <RANKING order="11" place="11" resultid="108250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99922" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110273" />
                    <RANKING order="2" place="2" resultid="107935" />
                    <RANKING order="3" place="3" resultid="106879" />
                    <RANKING order="4" place="4" resultid="108931" />
                    <RANKING order="5" place="5" resultid="107139" />
                    <RANKING order="6" place="6" resultid="107154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99923" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109069" />
                    <RANKING order="2" place="2" resultid="109403" />
                    <RANKING order="3" place="3" resultid="109582" />
                    <RANKING order="4" place="4" resultid="107078" />
                    <RANKING order="5" place="5" resultid="107002" />
                    <RANKING order="6" place="6" resultid="106867" />
                    <RANKING order="7" place="7" resultid="106858" />
                    <RANKING order="8" place="8" resultid="106614" />
                    <RANKING order="9" place="9" resultid="110089" />
                    <RANKING order="10" place="10" resultid="108919" />
                    <RANKING order="11" place="11" resultid="110411" />
                    <RANKING order="12" place="-1" resultid="110482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99924" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109850" />
                    <RANKING order="2" place="2" resultid="108026" />
                    <RANKING order="3" place="3" resultid="108209" />
                    <RANKING order="4" place="4" resultid="109858" />
                    <RANKING order="5" place="5" resultid="110493" />
                    <RANKING order="6" place="6" resultid="109395" />
                    <RANKING order="7" place="7" resultid="106833" />
                    <RANKING order="8" place="-1" resultid="109367" />
                    <RANKING order="9" place="-1" resultid="106840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99925" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106412" />
                    <RANKING order="2" place="2" resultid="107766" />
                    <RANKING order="3" place="3" resultid="107099" />
                    <RANKING order="4" place="4" resultid="107494" />
                    <RANKING order="5" place="5" resultid="110527" />
                    <RANKING order="6" place="6" resultid="108073" />
                    <RANKING order="7" place="7" resultid="108579" />
                    <RANKING order="8" place="-1" resultid="110503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99926" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109382" />
                    <RANKING order="2" place="2" resultid="108534" />
                    <RANKING order="3" place="3" resultid="107793" />
                    <RANKING order="4" place="4" resultid="106816" />
                    <RANKING order="5" place="5" resultid="107443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99927" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109418" />
                    <RANKING order="2" place="2" resultid="110521" />
                    <RANKING order="3" place="3" resultid="108588" />
                    <RANKING order="4" place="-1" resultid="107783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99928" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106689" />
                    <RANKING order="2" place="2" resultid="106350" />
                    <RANKING order="3" place="3" resultid="108484" />
                    <RANKING order="4" place="4" resultid="108515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99929" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99930" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99931" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110769" daytime="18:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110770" daytime="18:19" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110771" daytime="18:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110772" daytime="18:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110773" daytime="18:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110774" daytime="18:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110775" daytime="18:39" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110776" daytime="18:42" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110777" daytime="18:46" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="110778" daytime="18:49" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99170" daytime="16:58" gender="M" number="25" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99857" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107114" />
                    <RANKING order="2" place="2" resultid="109214" />
                    <RANKING order="3" place="3" resultid="107544" />
                    <RANKING order="4" place="4" resultid="110535" />
                    <RANKING order="5" place="5" resultid="107107" />
                    <RANKING order="6" place="6" resultid="110417" />
                    <RANKING order="7" place="7" resultid="108704" />
                    <RANKING order="8" place="8" resultid="108693" />
                    <RANKING order="9" place="9" resultid="110562" />
                    <RANKING order="10" place="-1" resultid="109314" />
                    <RANKING order="11" place="-1" resultid="110512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99858" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106655" />
                    <RANKING order="2" place="2" resultid="107191" />
                    <RANKING order="3" place="3" resultid="109477" />
                    <RANKING order="4" place="4" resultid="106441" />
                    <RANKING order="5" place="5" resultid="110144" />
                    <RANKING order="6" place="6" resultid="107722" />
                    <RANKING order="7" place="7" resultid="107249" />
                    <RANKING order="8" place="8" resultid="106661" />
                    <RANKING order="9" place="9" resultid="107631" />
                    <RANKING order="10" place="10" resultid="110389" />
                    <RANKING order="11" place="11" resultid="110581" />
                    <RANKING order="12" place="12" resultid="108699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99859" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107200" />
                    <RANKING order="2" place="2" resultid="107418" />
                    <RANKING order="3" place="3" resultid="107401" />
                    <RANKING order="4" place="4" resultid="107258" />
                    <RANKING order="5" place="5" resultid="108653" />
                    <RANKING order="6" place="6" resultid="108573" />
                    <RANKING order="7" place="7" resultid="107612" />
                    <RANKING order="8" place="8" resultid="107409" />
                    <RANKING order="9" place="9" resultid="110863" />
                    <RANKING order="10" place="10" resultid="108632" />
                    <RANKING order="11" place="11" resultid="109357" />
                    <RANKING order="12" place="12" resultid="107505" />
                    <RANKING order="13" place="13" resultid="109834" />
                    <RANKING order="14" place="-1" resultid="107621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99860" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107236" />
                    <RANKING order="2" place="2" resultid="107727" />
                    <RANKING order="3" place="3" resultid="107667" />
                    <RANKING order="4" place="4" resultid="108052" />
                    <RANKING order="5" place="4" resultid="109611" />
                    <RANKING order="6" place="6" resultid="107557" />
                    <RANKING order="7" place="7" resultid="107572" />
                    <RANKING order="8" place="8" resultid="107185" />
                    <RANKING order="9" place="9" resultid="106582" />
                    <RANKING order="10" place="10" resultid="106969" />
                    <RANKING order="11" place="11" resultid="107600" />
                    <RANKING order="12" place="12" resultid="107627" />
                    <RANKING order="13" place="13" resultid="109077" />
                    <RANKING order="14" place="-1" resultid="109151" />
                    <RANKING order="15" place="-1" resultid="109386" />
                    <RANKING order="16" place="-1" resultid="110248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99861" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109034" />
                    <RANKING order="2" place="2" resultid="106574" />
                    <RANKING order="3" place="3" resultid="109867" />
                    <RANKING order="4" place="4" resultid="110123" />
                    <RANKING order="5" place="5" resultid="108974" />
                    <RANKING order="6" place="6" resultid="108402" />
                    <RANKING order="7" place="7" resultid="107549" />
                    <RANKING order="8" place="8" resultid="108555" />
                    <RANKING order="9" place="9" resultid="108992" />
                    <RANKING order="10" place="10" resultid="107845" />
                    <RANKING order="11" place="11" resultid="106702" />
                    <RANKING order="12" place="12" resultid="108662" />
                    <RANKING order="13" place="13" resultid="110574" />
                    <RANKING order="14" place="14" resultid="109141" />
                    <RANKING order="15" place="15" resultid="109961" />
                    <RANKING order="16" place="-1" resultid="108985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99862" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110259" />
                    <RANKING order="2" place="2" resultid="107833" />
                    <RANKING order="3" place="3" resultid="108375" />
                    <RANKING order="4" place="4" resultid="109013" />
                    <RANKING order="5" place="5" resultid="109947" />
                    <RANKING order="6" place="6" resultid="107868" />
                    <RANKING order="7" place="7" resultid="107138" />
                    <RANKING order="8" place="-1" resultid="108426" />
                    <RANKING order="9" place="-1" resultid="106952" />
                    <RANKING order="10" place="-1" resultid="108928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99863" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110481" />
                    <RANKING order="2" place="2" resultid="109062" />
                    <RANKING order="3" place="3" resultid="108184" />
                    <RANKING order="4" place="4" resultid="109503" />
                    <RANKING order="5" place="5" resultid="106853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99864" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109849" />
                    <RANKING order="2" place="2" resultid="108025" />
                    <RANKING order="3" place="3" resultid="110081" />
                    <RANKING order="4" place="4" resultid="110492" />
                    <RANKING order="5" place="5" resultid="109394" />
                    <RANKING order="6" place="6" resultid="108243" />
                    <RANKING order="7" place="-1" resultid="106839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99865" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110541" />
                    <RANKING order="2" place="2" resultid="107493" />
                    <RANKING order="3" place="3" resultid="108262" />
                    <RANKING order="4" place="-1" resultid="107975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99866" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106407" />
                    <RANKING order="2" place="2" resultid="106707" />
                    <RANKING order="3" place="3" resultid="108034" />
                    <RANKING order="4" place="4" resultid="106810" />
                    <RANKING order="5" place="5" resultid="109471" />
                    <RANKING order="6" place="6" resultid="106718" />
                    <RANKING order="7" place="7" resultid="110365" />
                    <RANKING order="8" place="-1" resultid="107792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99867" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107776" />
                    <RANKING order="2" place="2" resultid="110520" />
                    <RANKING order="3" place="3" resultid="108587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99868" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107999" />
                    <RANKING order="2" place="2" resultid="108175" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99869" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99870" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99871" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110741" daytime="16:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110742" daytime="17:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110743" daytime="17:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110744" daytime="17:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110745" daytime="17:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110746" daytime="17:07" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110747" daytime="17:08" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110748" daytime="17:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110749" daytime="17:11" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="110750" daytime="17:13" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="110751" daytime="17:14" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99089" daytime="16:00" gender="F" number="22" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99109" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107943" />
                    <RANKING order="2" place="2" resultid="110403" />
                    <RANKING order="3" place="3" resultid="108958" />
                    <RANKING order="4" place="-1" resultid="110443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99110" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106668" />
                    <RANKING order="2" place="2" resultid="107674" />
                    <RANKING order="3" place="3" resultid="108219" />
                    <RANKING order="4" place="4" resultid="108646" />
                    <RANKING order="5" place="5" resultid="110568" />
                    <RANKING order="6" place="6" resultid="107381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99111" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107485" />
                    <RANKING order="2" place="2" resultid="110311" />
                    <RANKING order="3" place="3" resultid="107873" />
                    <RANKING order="4" place="4" resultid="109922" />
                    <RANKING order="5" place="5" resultid="106989" />
                    <RANKING order="6" place="6" resultid="109050" />
                    <RANKING order="7" place="-1" resultid="108669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99112" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106786" />
                    <RANKING order="2" place="2" resultid="107716" />
                    <RANKING order="3" place="3" resultid="109019" />
                    <RANKING order="4" place="4" resultid="106793" />
                    <RANKING order="5" place="5" resultid="110240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99113" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106711" />
                    <RANKING order="2" place="2" resultid="110131" />
                    <RANKING order="3" place="3" resultid="110138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99114" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107857" />
                    <RANKING order="2" place="2" resultid="108435" />
                    <RANKING order="3" place="3" resultid="107863" />
                    <RANKING order="4" place="4" resultid="107043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99115" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109447" />
                    <RANKING order="2" place="2" resultid="110105" />
                    <RANKING order="3" place="3" resultid="108043" />
                    <RANKING order="4" place="4" resultid="106768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99116" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109530" />
                    <RANKING order="2" place="2" resultid="109178" />
                    <RANKING order="3" place="3" resultid="106961" />
                    <RANKING order="4" place="4" resultid="106423" />
                    <RANKING order="5" place="5" resultid="109979" />
                    <RANKING order="6" place="6" resultid="110174" />
                    <RANKING order="7" place="7" resultid="110232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99117" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107085" />
                    <RANKING order="2" place="2" resultid="107471" />
                    <RANKING order="3" place="3" resultid="109909" />
                    <RANKING order="4" place="4" resultid="110357" />
                    <RANKING order="5" place="-1" resultid="106750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99118" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108471" />
                    <RANKING order="2" place="2" resultid="110474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99119" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99120" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106743" />
                    <RANKING order="2" place="2" resultid="107808" />
                    <RANKING order="3" place="3" resultid="107800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99121" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99122" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99123" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110720" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110721" daytime="16:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110722" daytime="16:11" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110723" daytime="16:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110724" daytime="16:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110725" daytime="16:19" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99202" daytime="17:51" gender="F" number="28" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99902" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107944" />
                    <RANKING order="2" place="2" resultid="107374" />
                    <RANKING order="3" place="3" resultid="108641" />
                    <RANKING order="4" place="4" resultid="110377" />
                    <RANKING order="5" place="5" resultid="108959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99903" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110281" />
                    <RANKING order="2" place="2" resultid="107382" />
                    <RANKING order="3" place="3" resultid="109081" />
                    <RANKING order="4" place="-1" resultid="106802" />
                    <RANKING order="5" place="-1" resultid="107205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99904" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107230" />
                    <RANKING order="2" place="2" resultid="109923" />
                    <RANKING order="3" place="3" resultid="106589" />
                    <RANKING order="4" place="4" resultid="110300" />
                    <RANKING order="5" place="5" resultid="109877" />
                    <RANKING order="6" place="6" resultid="109051" />
                    <RANKING order="7" place="7" resultid="106436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99905" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107962" />
                    <RANKING order="2" place="2" resultid="107709" />
                    <RANKING order="3" place="3" resultid="108685" />
                    <RANKING order="4" place="4" resultid="108967" />
                    <RANKING order="5" place="5" resultid="110307" />
                    <RANKING order="6" place="6" resultid="110241" />
                    <RANKING order="7" place="-1" resultid="106596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99906" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106712" />
                    <RANKING order="2" place="2" resultid="110132" />
                    <RANKING order="3" place="3" resultid="107919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99907" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109826" />
                    <RANKING order="2" place="2" resultid="109917" />
                    <RANKING order="3" place="-1" resultid="108568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99908" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108197" />
                    <RANKING order="2" place="2" resultid="107991" />
                    <RANKING order="3" place="3" resultid="109448" />
                    <RANKING order="4" place="4" resultid="108044" />
                    <RANKING order="5" place="5" resultid="109510" />
                    <RANKING order="6" place="6" resultid="106776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99909" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108507" />
                    <RANKING order="2" place="2" resultid="110225" />
                    <RANKING order="3" place="3" resultid="109980" />
                    <RANKING order="4" place="4" resultid="108458" />
                    <RANKING order="5" place="-1" resultid="106755" />
                    <RANKING order="6" place="-1" resultid="106962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99910" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99911" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99912" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99913" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99914" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99915" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99916" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110764" daytime="17:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110765" daytime="17:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110766" daytime="18:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110767" daytime="18:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110768" daytime="18:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-10-23" daytime="09:00" endtime="13:13" number="4" warmupfrom="08:00" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="99361" daytime="09:12" gender="M" number="35" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99977" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107115" />
                    <RANKING order="2" place="2" resultid="109215" />
                    <RANKING order="3" place="3" resultid="109540" />
                    <RANKING order="4" place="4" resultid="110536" />
                    <RANKING order="5" place="5" resultid="109906" />
                    <RANKING order="6" place="6" resultid="108706" />
                    <RANKING order="7" place="-1" resultid="110513" />
                    <RANKING order="8" place="-1" resultid="110563" />
                    <RANKING order="9" place="-1" resultid="110857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99978" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106656" />
                    <RANKING order="2" place="2" resultid="109891" />
                    <RANKING order="3" place="3" resultid="109479" />
                    <RANKING order="4" place="4" resultid="110390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99979" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107420" />
                    <RANKING order="2" place="2" resultid="106979" />
                    <RANKING order="3" place="3" resultid="109578" />
                    <RANKING order="4" place="4" resultid="107403" />
                    <RANKING order="5" place="5" resultid="109970" />
                    <RANKING order="6" place="6" resultid="107411" />
                    <RANKING order="7" place="-1" resultid="107623" />
                    <RANKING order="8" place="-1" resultid="108633" />
                    <RANKING order="9" place="-1" resultid="109359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99980" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107238" />
                    <RANKING order="2" place="2" resultid="107729" />
                    <RANKING order="3" place="3" resultid="107669" />
                    <RANKING order="4" place="4" resultid="109558" />
                    <RANKING order="5" place="5" resultid="108054" />
                    <RANKING order="6" place="6" resultid="107573" />
                    <RANKING order="7" place="7" resultid="107559" />
                    <RANKING order="8" place="8" resultid="106971" />
                    <RANKING order="9" place="-1" resultid="109444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99981" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109869" />
                    <RANKING order="2" place="2" resultid="108976" />
                    <RANKING order="3" place="3" resultid="110125" />
                    <RANKING order="4" place="4" resultid="106703" />
                    <RANKING order="5" place="5" resultid="107748" />
                    <RANKING order="6" place="6" resultid="109143" />
                    <RANKING order="7" place="7" resultid="110576" />
                    <RANKING order="8" place="-1" resultid="106576" />
                    <RANKING order="9" place="-1" resultid="108986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99982" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110261" />
                    <RANKING order="2" place="2" resultid="109028" />
                    <RANKING order="3" place="3" resultid="108929" />
                    <RANKING order="4" place="4" resultid="107834" />
                    <RANKING order="5" place="-1" resultid="106954" />
                    <RANKING order="6" place="-1" resultid="107140" />
                    <RANKING order="7" place="-1" resultid="107758" />
                    <RANKING order="8" place="-1" resultid="108376" />
                    <RANKING order="9" place="-1" resultid="108428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99983" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109070" />
                    <RANKING order="2" place="2" resultid="109404" />
                    <RANKING order="3" place="3" resultid="110485" />
                    <RANKING order="4" place="4" resultid="109064" />
                    <RANKING order="5" place="5" resultid="110267" />
                    <RANKING order="6" place="6" resultid="107003" />
                    <RANKING order="7" place="7" resultid="108186" />
                    <RANKING order="8" place="8" resultid="106868" />
                    <RANKING order="9" place="9" resultid="110090" />
                    <RANKING order="10" place="10" resultid="106616" />
                    <RANKING order="11" place="11" resultid="109437" />
                    <RANKING order="12" place="-1" resultid="109583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99984" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109851" />
                    <RANKING order="2" place="2" resultid="108027" />
                    <RANKING order="3" place="3" resultid="109323" />
                    <RANKING order="4" place="4" resultid="109860" />
                    <RANKING order="5" place="5" resultid="110082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99985" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108160" />
                    <RANKING order="2" place="2" resultid="107100" />
                    <RANKING order="3" place="3" resultid="107132" />
                    <RANKING order="4" place="4" resultid="108263" />
                    <RANKING order="5" place="5" resultid="108075" />
                    <RANKING order="6" place="-1" resultid="108237" />
                    <RANKING order="7" place="-1" resultid="107976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99986" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106408" />
                    <RANKING order="2" place="2" resultid="106811" />
                    <RANKING order="3" place="3" resultid="108036" />
                    <RANKING order="4" place="4" resultid="108536" />
                    <RANKING order="5" place="5" resultid="108169" />
                    <RANKING order="6" place="6" resultid="110367" />
                    <RANKING order="7" place="7" resultid="107445" />
                    <RANKING order="8" place="-1" resultid="107794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99987" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107777" />
                    <RANKING order="2" place="2" resultid="110522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99988" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108000" />
                    <RANKING order="2" place="2" resultid="106690" />
                    <RANKING order="3" place="3" resultid="108177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99989" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99990" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99991" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110797" daytime="09:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110798" daytime="09:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110799" daytime="09:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110800" daytime="09:21" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110801" daytime="09:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110802" daytime="09:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110803" daytime="09:28" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110804" daytime="09:30" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110805" daytime="09:33" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99393" daytime="09:56" gender="M" number="37" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100007" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107546" />
                    <RANKING order="2" place="2" resultid="110437" />
                    <RANKING order="3" place="3" resultid="107927" />
                    <RANKING order="4" place="4" resultid="108952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100008" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107174" />
                    <RANKING order="2" place="2" resultid="106663" />
                    <RANKING order="3" place="3" resultid="110293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100009" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107421" />
                    <RANKING order="2" place="2" resultid="110470" />
                    <RANKING order="3" place="3" resultid="109579" />
                    <RANKING order="4" place="4" resultid="107567" />
                    <RANKING order="5" place="5" resultid="110423" />
                    <RANKING order="6" place="6" resultid="110463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100010" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107239" />
                    <RANKING order="2" place="2" resultid="107730" />
                    <RANKING order="3" place="3" resultid="109565" />
                    <RANKING order="4" place="4" resultid="108060" />
                    <RANKING order="5" place="5" resultid="107700" />
                    <RANKING order="6" place="6" resultid="106603" />
                    <RANKING order="7" place="7" resultid="108413" />
                    <RANKING order="8" place="8" resultid="107954" />
                    <RANKING order="9" place="-1" resultid="107586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100011" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108404" />
                    <RANKING order="2" place="2" resultid="110159" />
                    <RANKING order="3" place="3" resultid="110399" />
                    <RANKING order="4" place="4" resultid="107550" />
                    <RANKING order="5" place="-1" resultid="109342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100012" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107739" />
                    <RANKING order="2" place="2" resultid="106887" />
                    <RANKING order="3" place="3" resultid="110167" />
                    <RANKING order="4" place="4" resultid="109174" />
                    <RANKING order="5" place="5" resultid="107691" />
                    <RANKING order="6" place="-1" resultid="106955" />
                    <RANKING order="7" place="-1" resultid="107155" />
                    <RANKING order="8" place="-1" resultid="108429" />
                    <RANKING order="9" place="-1" resultid="109949" />
                    <RANKING order="10" place="-1" resultid="110262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100013" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109405" />
                    <RANKING order="2" place="2" resultid="109518" />
                    <RANKING order="3" place="3" resultid="109504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100014" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107029" />
                    <RANKING order="2" place="2" resultid="108446" />
                    <RANKING order="3" place="3" resultid="108231" />
                    <RANKING order="4" place="4" resultid="108245" />
                    <RANKING order="5" place="-1" resultid="108028" />
                    <RANKING order="6" place="-1" resultid="108356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100015" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109411" />
                    <RANKING order="2" place="2" resultid="110073" />
                    <RANKING order="3" place="3" resultid="108161" />
                    <RANKING order="4" place="4" resultid="110454" />
                    <RANKING order="5" place="5" resultid="108580" />
                    <RANKING order="6" place="-1" resultid="110504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100016" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109375" />
                    <RANKING order="2" place="2" resultid="106724" />
                    <RANKING order="3" place="3" resultid="110065" />
                    <RANKING order="4" place="4" resultid="107446" />
                    <RANKING order="5" place="-1" resultid="108366" />
                    <RANKING order="6" place="-1" resultid="109816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100017" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110059" />
                    <RANKING order="2" place="2" resultid="109419" />
                    <RANKING order="3" place="3" resultid="108523" />
                    <RANKING order="4" place="-1" resultid="108589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100018" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108178" />
                    <RANKING order="2" place="2" resultid="107074" />
                    <RANKING order="3" place="3" resultid="107452" />
                    <RANKING order="4" place="-1" resultid="109350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100019" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100020" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100021" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110810" daytime="09:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110811" daytime="10:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110812" daytime="10:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110813" daytime="10:13" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110814" daytime="10:17" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110815" daytime="10:21" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110816" daytime="10:24" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99425" daytime="10:41" gender="M" number="39" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100037" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110537" />
                    <RANKING order="2" place="2" resultid="108953" />
                    <RANKING order="3" place="3" resultid="110564" />
                    <RANKING order="4" place="4" resultid="108694" />
                    <RANKING order="5" place="-1" resultid="109313" />
                    <RANKING order="6" place="-1" resultid="110514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100038" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107178" />
                    <RANKING order="2" place="2" resultid="109006" />
                    <RANKING order="3" place="3" resultid="110294" />
                    <RANKING order="4" place="4" resultid="107880" />
                    <RANKING order="5" place="5" resultid="110391" />
                    <RANKING order="6" place="6" resultid="107852" />
                    <RANKING order="7" place="7" resultid="108700" />
                    <RANKING order="8" place="-1" resultid="106608" />
                    <RANKING order="9" place="-1" resultid="107197" />
                    <RANKING order="10" place="-1" resultid="110145" />
                    <RANKING order="11" place="-1" resultid="110582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100039" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107395" />
                    <RANKING order="2" place="2" resultid="107120" />
                    <RANKING order="3" place="3" resultid="107513" />
                    <RANKING order="4" place="4" resultid="107568" />
                    <RANKING order="5" place="5" resultid="107613" />
                    <RANKING order="6" place="6" resultid="107404" />
                    <RANKING order="7" place="7" resultid="109971" />
                    <RANKING order="8" place="8" resultid="108655" />
                    <RANKING order="9" place="9" resultid="107412" />
                    <RANKING order="10" place="10" resultid="110424" />
                    <RANKING order="11" place="11" resultid="109843" />
                    <RANKING order="12" place="-1" resultid="108634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100040" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109957" />
                    <RANKING order="2" place="2" resultid="108055" />
                    <RANKING order="3" place="3" resultid="107670" />
                    <RANKING order="4" place="4" resultid="109612" />
                    <RANKING order="5" place="5" resultid="107601" />
                    <RANKING order="6" place="6" resultid="109078" />
                    <RANKING order="7" place="7" resultid="107438" />
                    <RANKING order="8" place="8" resultid="107595" />
                    <RANKING order="9" place="9" resultid="108594" />
                    <RANKING order="10" place="10" resultid="107955" />
                    <RANKING order="11" place="-1" resultid="106584" />
                    <RANKING order="12" place="-1" resultid="107578" />
                    <RANKING order="13" place="-1" resultid="107587" />
                    <RANKING order="14" place="-1" resultid="107606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100041" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108421" />
                    <RANKING order="2" place="2" resultid="108977" />
                    <RANKING order="3" place="3" resultid="107846" />
                    <RANKING order="4" place="4" resultid="109035" />
                    <RANKING order="5" place="5" resultid="108987" />
                    <RANKING order="6" place="6" resultid="110126" />
                    <RANKING order="7" place="7" resultid="108993" />
                    <RANKING order="8" place="8" resultid="108556" />
                    <RANKING order="9" place="9" resultid="108664" />
                    <RANKING order="10" place="-1" resultid="107970" />
                    <RANKING order="11" place="-1" resultid="108405" />
                    <RANKING order="12" place="-1" resultid="108562" />
                    <RANKING order="13" place="-1" resultid="110190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100042" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107936" />
                    <RANKING order="2" place="2" resultid="109029" />
                    <RANKING order="3" place="3" resultid="109014" />
                    <RANKING order="4" place="4" resultid="110168" />
                    <RANKING order="5" place="5" resultid="110429" />
                    <RANKING order="6" place="-1" resultid="106880" />
                    <RANKING order="7" place="-1" resultid="107156" />
                    <RANKING order="8" place="-1" resultid="108377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100043" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106869" />
                    <RANKING order="2" place="2" resultid="109065" />
                    <RANKING order="3" place="3" resultid="110091" />
                    <RANKING order="4" place="4" resultid="106859" />
                    <RANKING order="5" place="5" resultid="110486" />
                    <RANKING order="6" place="6" resultid="109571" />
                    <RANKING order="7" place="7" resultid="106849" />
                    <RANKING order="8" place="8" resultid="106875" />
                    <RANKING order="9" place="9" resultid="110268" />
                    <RANKING order="10" place="10" resultid="109438" />
                    <RANKING order="11" place="11" resultid="110412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100044" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107010" />
                    <RANKING order="2" place="2" resultid="109324" />
                    <RANKING order="3" place="3" resultid="106828" />
                    <RANKING order="4" place="4" resultid="108357" />
                    <RANKING order="5" place="5" resultid="110083" />
                    <RANKING order="6" place="-1" resultid="108246" />
                    <RANKING order="7" place="-1" resultid="109368" />
                    <RANKING order="8" place="-1" resultid="106841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100045" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107133" />
                    <RANKING order="2" place="2" resultid="108204" />
                    <RANKING order="3" place="3" resultid="108477" />
                    <RANKING order="4" place="4" resultid="107500" />
                    <RANKING order="5" place="5" resultid="107767" />
                    <RANKING order="6" place="6" resultid="108257" />
                    <RANKING order="7" place="7" resultid="108581" />
                    <RANKING order="8" place="-1" resultid="106822" />
                    <RANKING order="9" place="-1" resultid="108238" />
                    <RANKING order="10" place="-1" resultid="107977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100046" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108011" />
                    <RANKING order="2" place="2" resultid="110152" />
                    <RANKING order="3" place="3" resultid="109817" />
                    <RANKING order="4" place="4" resultid="109984" />
                    <RANKING order="5" place="5" resultid="110368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100047" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107778" />
                    <RANKING order="2" place="2" resultid="110060" />
                    <RANKING order="3" place="3" resultid="107462" />
                    <RANKING order="4" place="4" resultid="107147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100048" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108001" />
                    <RANKING order="2" place="2" resultid="108485" />
                    <RANKING order="3" place="3" resultid="108516" />
                    <RANKING order="4" place="4" resultid="107075" />
                    <RANKING order="5" place="5" resultid="107455" />
                    <RANKING order="6" place="-1" resultid="109351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100049" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100050" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100051" agemax="94" agemin="90" name="KAT.N, 90-94 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="108006" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110824" daytime="10:41" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110825" daytime="10:43" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110826" daytime="10:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110827" daytime="10:47" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110828" daytime="10:49" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110829" daytime="10:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110830" daytime="10:52" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110831" daytime="10:54" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110832" daytime="10:55" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="110833" daytime="10:57" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="110834" daytime="10:59" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99473" daytime="11:50" gender="M" number="42" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100067" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109541" />
                    <RANKING order="2" place="2" resultid="107109" />
                    <RANKING order="3" place="3" resultid="110438" />
                    <RANKING order="4" place="4" resultid="106675" />
                    <RANKING order="5" place="-1" resultid="107928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100068" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109892" />
                    <RANKING order="2" place="2" resultid="106402" />
                    <RANKING order="3" place="3" resultid="110384" />
                    <RANKING order="4" place="4" resultid="107682" />
                    <RANKING order="5" place="-1" resultid="106651" />
                    <RANKING order="6" place="-1" resultid="109007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100069" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107514" />
                    <RANKING order="2" place="2" resultid="106980" />
                    <RANKING order="3" place="3" resultid="109524" />
                    <RANKING order="4" place="4" resultid="108656" />
                    <RANKING order="5" place="5" resultid="109360" />
                    <RANKING order="6" place="6" resultid="106641" />
                    <RANKING order="7" place="7" resultid="110464" />
                    <RANKING order="8" place="8" resultid="107507" />
                    <RANKING order="9" place="9" resultid="107480" />
                    <RANKING order="10" place="-1" resultid="109461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100070" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109559" />
                    <RANKING order="2" place="2" resultid="107560" />
                    <RANKING order="3" place="3" resultid="109388" />
                    <RANKING order="4" place="4" resultid="109938" />
                    <RANKING order="5" place="5" resultid="107701" />
                    <RANKING order="6" place="6" resultid="106635" />
                    <RANKING order="7" place="-1" resultid="107596" />
                    <RANKING order="8" place="-1" resultid="108414" />
                    <RANKING order="9" place="-1" resultid="110250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100071" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109870" />
                    <RANKING order="2" place="2" resultid="107749" />
                    <RANKING order="3" place="3" resultid="106577" />
                    <RANKING order="4" place="4" resultid="109466" />
                    <RANKING order="5" place="5" resultid="109001" />
                    <RANKING order="6" place="6" resultid="109144" />
                    <RANKING order="7" place="7" resultid="110400" />
                    <RANKING order="8" place="8" resultid="110497" />
                    <RANKING order="9" place="9" resultid="110160" />
                    <RANKING order="10" place="10" resultid="108665" />
                    <RANKING order="11" place="11" resultid="109963" />
                    <RANKING order="12" place="12" resultid="108251" />
                    <RANKING order="13" place="-1" resultid="109343" />
                    <RANKING order="14" place="-1" resultid="109886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100072" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110275" />
                    <RANKING order="2" place="2" resultid="106881" />
                    <RANKING order="3" place="3" resultid="109950" />
                    <RANKING order="4" place="4" resultid="107692" />
                    <RANKING order="5" place="-1" resultid="107141" />
                    <RANKING order="6" place="-1" resultid="107937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100073" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109584" />
                    <RANKING order="2" place="2" resultid="107079" />
                    <RANKING order="3" place="3" resultid="107004" />
                    <RANKING order="4" place="4" resultid="109168" />
                    <RANKING order="5" place="5" resultid="109519" />
                    <RANKING order="6" place="6" resultid="106860" />
                    <RANKING order="7" place="7" resultid="106850" />
                    <RANKING order="8" place="8" resultid="106617" />
                    <RANKING order="9" place="9" resultid="108921" />
                    <RANKING order="10" place="10" resultid="110413" />
                    <RANKING order="11" place="-1" resultid="108187" />
                    <RANKING order="12" place="-1" resultid="109071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100074" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109852" />
                    <RANKING order="2" place="2" resultid="108210" />
                    <RANKING order="3" place="3" resultid="109861" />
                    <RANKING order="4" place="4" resultid="109396" />
                    <RANKING order="5" place="-1" resultid="106834" />
                    <RANKING order="6" place="-1" resultid="108447" />
                    <RANKING order="7" place="-1" resultid="109369" />
                    <RANKING order="8" place="-1" resultid="110494" />
                    <RANKING order="9" place="-1" resultid="106842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100075" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106413" />
                    <RANKING order="2" place="2" resultid="107101" />
                    <RANKING order="3" place="3" resultid="110074" />
                    <RANKING order="4" place="4" resultid="107495" />
                    <RANKING order="5" place="5" resultid="110455" />
                    <RANKING order="6" place="6" resultid="110528" />
                    <RANKING order="7" place="7" resultid="108076" />
                    <RANKING order="8" place="-1" resultid="107768" />
                    <RANKING order="9" place="-1" resultid="110505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100076" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109383" />
                    <RANKING order="2" place="2" resultid="106940" />
                    <RANKING order="3" place="3" resultid="108537" />
                    <RANKING order="4" place="4" resultid="107795" />
                    <RANKING order="5" place="5" resultid="106817" />
                    <RANKING order="6" place="6" resultid="109997" />
                    <RANKING order="7" place="-1" resultid="108037" />
                    <RANKING order="8" place="-1" resultid="108170" />
                    <RANKING order="9" place="-1" resultid="108367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100077" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110523" />
                    <RANKING order="2" place="2" resultid="109420" />
                    <RANKING order="3" place="-1" resultid="107785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100078" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106351" />
                    <RANKING order="2" place="2" resultid="108517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100079" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100080" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100081" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110843" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110844" daytime="11:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110845" daytime="12:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110846" daytime="12:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110847" daytime="12:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110848" daytime="12:21" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110849" daytime="12:28" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="110850" daytime="12:36" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="110851" daytime="12:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="110852" daytime="12:53" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99344" daytime="09:00" gender="F" number="34" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99962" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107945" />
                    <RANKING order="2" place="2" resultid="108678" />
                    <RANKING order="3" place="3" resultid="109899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99963" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109992" />
                    <RANKING order="2" place="2" resultid="108221" />
                    <RANKING order="3" place="3" resultid="108907" />
                    <RANKING order="4" place="-1" resultid="106803" />
                    <RANKING order="5" place="-1" resultid="109426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99964" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110301" />
                    <RANKING order="2" place="2" resultid="108627" />
                    <RANKING order="3" place="3" resultid="106590" />
                    <RANKING order="4" place="4" resultid="109878" />
                    <RANKING order="5" place="5" resultid="106991" />
                    <RANKING order="6" place="6" resultid="107036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99965" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108272" />
                    <RANKING order="2" place="2" resultid="107710" />
                    <RANKING order="3" place="3" resultid="108686" />
                    <RANKING order="4" place="4" resultid="108968" />
                    <RANKING order="5" place="-1" resultid="106646" />
                    <RANKING order="6" place="-1" resultid="109021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99966" agemax="44" agemin="40" name="KAT.D, 40-44 lat" />
                <AGEGROUP agegroupid="99967" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108081" />
                    <RANKING order="2" place="2" resultid="108437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99968" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108528" />
                    <RANKING order="2" place="2" resultid="110107" />
                    <RANKING order="3" place="3" resultid="108018" />
                    <RANKING order="4" place="4" resultid="106770" />
                    <RANKING order="5" place="5" resultid="109549" />
                    <RANKING order="6" place="-1" resultid="106763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99969" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109180" />
                    <RANKING order="2" place="2" resultid="108508" />
                    <RANKING order="3" place="3" resultid="110234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99970" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107908" />
                    <RANKING order="2" place="2" resultid="108465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99971" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99972" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99973" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99974" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99975" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99976" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110793" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110794" daytime="09:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110795" daytime="09:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110796" daytime="09:09" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99457" daytime="11:16" gender="F" number="41" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100052" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107376" />
                    <RANKING order="2" place="2" resultid="108642" />
                    <RANKING order="3" place="3" resultid="110379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100053" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109993" />
                    <RANKING order="2" place="2" resultid="110283" />
                    <RANKING order="3" place="3" resultid="108908" />
                    <RANKING order="4" place="4" resultid="109082" />
                    <RANKING order="5" place="-1" resultid="110571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100054" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107232" />
                    <RANKING order="2" place="2" resultid="107488" />
                    <RANKING order="3" place="3" resultid="107389" />
                    <RANKING order="4" place="4" resultid="109879" />
                    <RANKING order="5" place="5" resultid="109924" />
                    <RANKING order="6" place="6" resultid="110302" />
                    <RANKING order="7" place="7" resultid="106437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100055" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107963" />
                    <RANKING order="2" place="2" resultid="110309" />
                    <RANKING order="3" place="3" resultid="106598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100056" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106714" />
                    <RANKING order="2" place="2" resultid="110466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100057" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109829" />
                    <RANKING order="2" place="2" resultid="107046" />
                    <RANKING order="3" place="3" resultid="109919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100058" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108199" />
                    <RANKING order="2" place="2" resultid="108926" />
                    <RANKING order="3" place="3" resultid="109450" />
                    <RANKING order="4" place="4" resultid="107993" />
                    <RANKING order="5" place="5" resultid="109511" />
                    <RANKING order="6" place="-1" resultid="108046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100059" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108509" />
                    <RANKING order="2" place="2" resultid="107094" />
                    <RANKING order="3" place="3" resultid="110177" />
                    <RANKING order="4" place="4" resultid="109981" />
                    <RANKING order="5" place="5" resultid="108459" />
                    <RANKING order="6" place="-1" resultid="106756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100060" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100061" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110100" />
                    <RANKING order="2" place="2" resultid="109432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100062" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="100063" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107019" />
                    <RANKING order="2" place="2" resultid="107818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100064" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="100065" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100066" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110839" daytime="11:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110840" daytime="11:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110841" daytime="11:29" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110842" daytime="11:37" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99377" daytime="09:35" gender="F" number="36" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99992" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108960" />
                    <RANKING order="2" place="-1" resultid="110445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99993" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="110282" />
                    <RANKING order="2" place="2" resultid="107913" />
                    <RANKING order="3" place="3" resultid="107383" />
                    <RANKING order="4" place="-1" resultid="109427" />
                    <RANKING order="5" place="-1" resultid="110570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99994" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107231" />
                    <RANKING order="2" place="2" resultid="107841" />
                    <RANKING order="3" place="3" resultid="107037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99995" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108687" />
                    <RANKING order="2" place="2" resultid="109931" />
                    <RANKING order="3" place="3" resultid="110183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99996" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108089" />
                    <RANKING order="2" place="2" resultid="106985" />
                    <RANKING order="3" place="3" resultid="108551" />
                    <RANKING order="4" place="4" resultid="107920" />
                    <RANKING order="5" place="5" resultid="109840" />
                    <RANKING order="6" place="6" resultid="107068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99997" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106783" />
                    <RANKING order="2" place="2" resultid="109828" />
                    <RANKING order="3" place="3" resultid="109918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99998" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108198" />
                    <RANKING order="2" place="2" resultid="107992" />
                    <RANKING order="3" place="3" resultid="108383" />
                    <RANKING order="4" place="4" resultid="109550" />
                    <RANKING order="5" place="-1" resultid="108019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99999" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107093" />
                    <RANKING order="2" place="2" resultid="108350" />
                    <RANKING order="3" place="3" resultid="110176" />
                    <RANKING order="4" place="4" resultid="110226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100000" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107909" />
                    <RANKING order="2" place="2" resultid="108466" />
                    <RANKING order="3" place="3" resultid="110359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100001" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109456" />
                    <RANKING order="2" place="2" resultid="110476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100002" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="100003" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107018" />
                    <RANKING order="2" place="2" resultid="109135" />
                    <RANKING order="3" place="3" resultid="107802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100004" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="100005" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100006" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110806" daytime="09:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110807" daytime="09:43" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110808" daytime="09:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110809" daytime="09:52" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99441" daytime="11:00" gender="X" number="40" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99540" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99541" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107264" />
                    <RANKING order="2" place="-1" resultid="106676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99542" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107732" />
                    <RANKING order="2" place="2" resultid="110316" />
                    <RANKING order="3" place="3" resultid="110013" />
                    <RANKING order="4" place="4" resultid="107423" />
                    <RANKING order="5" place="5" resultid="108713" />
                    <RANKING order="6" place="6" resultid="106994" />
                    <RANKING order="7" place="7" resultid="109037" />
                    <RANKING order="8" place="8" resultid="107523" />
                    <RANKING order="9" place="9" resultid="106621" />
                    <RANKING order="10" place="10" resultid="110199" />
                    <RANKING order="11" place="-1" resultid="106493" />
                    <RANKING order="12" place="-1" resultid="107263" />
                    <RANKING order="13" place="-1" resultid="107888" />
                    <RANKING order="14" place="-1" resultid="108715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99543" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108098" />
                    <RANKING order="2" place="2" resultid="107886" />
                    <RANKING order="3" place="3" resultid="109590" />
                    <RANKING order="4" place="4" resultid="110014" />
                    <RANKING order="5" place="5" resultid="110198" />
                    <RANKING order="6" place="6" resultid="107957" />
                    <RANKING order="7" place="-1" resultid="106903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99544" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108602" />
                    <RANKING order="2" place="2" resultid="110015" />
                    <RANKING order="3" place="3" resultid="108100" />
                    <RANKING order="4" place="4" resultid="106902" />
                    <RANKING order="5" place="-1" resultid="108598" />
                    <RANKING order="6" place="-1" resultid="110110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99545" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106901" />
                    <RANKING order="2" place="2" resultid="108102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99546" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106728" />
                    <RANKING order="2" place="2" resultid="108492" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110835" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110836" daytime="11:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110837" daytime="11:09" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110838" daytime="11:13" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99409" daytime="10:28" gender="F" number="38" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100022" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107946" />
                    <RANKING order="2" place="2" resultid="110405" />
                    <RANKING order="3" place="3" resultid="108961" />
                    <RANKING order="4" place="4" resultid="107375" />
                    <RANKING order="5" place="5" resultid="107124" />
                    <RANKING order="6" place="6" resultid="110378" />
                    <RANKING order="7" place="-1" resultid="110446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100023" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106670" />
                    <RANKING order="2" place="2" resultid="107675" />
                    <RANKING order="3" place="3" resultid="108222" />
                    <RANKING order="4" place="4" resultid="110286" />
                    <RANKING order="5" place="5" resultid="108647" />
                    <RANKING order="6" place="6" resultid="107384" />
                    <RANKING order="7" place="-1" resultid="106804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100024" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107487" />
                    <RANKING order="2" place="2" resultid="106992" />
                    <RANKING order="3" place="3" resultid="110865" />
                    <RANKING order="4" place="4" resultid="109052" />
                    <RANKING order="5" place="-1" resultid="108670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100025" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106788" />
                    <RANKING order="2" place="2" resultid="108273" />
                    <RANKING order="3" place="3" resultid="107718" />
                    <RANKING order="4" place="4" resultid="107711" />
                    <RANKING order="5" place="5" resultid="109022" />
                    <RANKING order="6" place="6" resultid="110308" />
                    <RANKING order="7" place="7" resultid="110242" />
                    <RANKING order="8" place="-1" resultid="106795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100026" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106713" />
                    <RANKING order="2" place="2" resultid="110133" />
                    <RANKING order="3" place="3" resultid="107921" />
                    <RANKING order="4" place="4" resultid="106428" />
                    <RANKING order="5" place="5" resultid="110140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100027" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107859" />
                    <RANKING order="2" place="2" resultid="108438" />
                    <RANKING order="3" place="3" resultid="107864" />
                    <RANKING order="4" place="4" resultid="107045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100028" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108500" />
                    <RANKING order="2" place="2" resultid="108045" />
                    <RANKING order="3" place="3" resultid="109449" />
                    <RANKING order="4" place="4" resultid="110108" />
                    <RANKING order="5" place="5" resultid="106771" />
                    <RANKING order="6" place="6" resultid="106777" />
                    <RANKING order="7" place="-1" resultid="106764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100029" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="109532" />
                    <RANKING order="2" place="2" resultid="109181" />
                    <RANKING order="3" place="3" resultid="106963" />
                    <RANKING order="4" place="4" resultid="106424" />
                    <RANKING order="5" place="5" resultid="110227" />
                    <RANKING order="6" place="6" resultid="110235" />
                    <RANKING order="7" place="-1" resultid="108387" />
                    <RANKING order="8" place="-1" resultid="108392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100030" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="107086" />
                    <RANKING order="2" place="2" resultid="108067" />
                    <RANKING order="3" place="3" resultid="109910" />
                    <RANKING order="4" place="4" resultid="107473" />
                    <RANKING order="5" place="-1" resultid="106751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100031" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106698" />
                    <RANKING order="2" place="2" resultid="108473" />
                    <RANKING order="3" place="3" resultid="107082" />
                    <RANKING order="4" place="4" resultid="110477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100032" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100033" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="106744" />
                    <RANKING order="2" place="2" resultid="107810" />
                    <RANKING order="3" place="3" resultid="107803" />
                    <RANKING order="4" place="-1" resultid="107817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100034" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="108194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100035" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100036" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="110817" daytime="10:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="110818" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="110819" daytime="10:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="110820" daytime="10:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="110821" daytime="10:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="110822" daytime="10:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="110823" daytime="10:40" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="RUS" clubid="106414" name="105 ELEMENT DUBNA">
          <ATHLETES>
            <ATHLETE birthdate="1959-01-01" firstname="IRINA" gender="F" lastname="MIGULINA" nation="RUS" athleteid="106415">
              <RESULTS>
                <RESULT eventid="98940" points="225" swimtime="00:03:40.95" resultid="106422" heatid="110662" lane="0" entrytime="00:03:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.46" />
                    <SPLIT distance="50" swimtime="00:00:49.14" />
                    <SPLIT distance="75" swimtime="00:01:16.59" />
                    <SPLIT distance="100" swimtime="00:01:45.52" />
                    <SPLIT distance="125" swimtime="00:02:13.90" />
                    <SPLIT distance="150" swimtime="00:02:43.64" />
                    <SPLIT distance="175" swimtime="00:03:12.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="230" reactiontime="+102" swimtime="00:01:41.72" resultid="106423" heatid="110722" lane="1" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.97" />
                    <SPLIT distance="50" swimtime="00:00:47.84" />
                    <SPLIT distance="75" swimtime="00:01:14.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="251" reactiontime="+95" swimtime="00:00:45.61" resultid="106424" heatid="110819" lane="5" entrytime="00:00:46.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-09-09" firstname="VARVARA" gender="F" lastname="KLIDZHAN" nation="RUS" athleteid="106417">
              <RESULTS>
                <RESULT eventid="98777" points="362" reactiontime="+87" swimtime="00:00:32.58" resultid="106429" heatid="110591" lane="8" entrytime="00:00:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="354" reactiontime="+84" swimtime="00:01:11.94" resultid="106430" heatid="110675" lane="2" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.17" />
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="75" swimtime="00:00:51.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-09-09" firstname="SVETLANA" gender="F" lastname="SMIRNOVA" nation="RUS" athleteid="106416">
              <RESULTS>
                <RESULT eventid="98814" points="267" reactiontime="+79" swimtime="00:03:09.04" resultid="106425" heatid="110616" lane="7" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.63" />
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                    <SPLIT distance="75" swimtime="00:01:08.61" />
                    <SPLIT distance="100" swimtime="00:01:33.46" />
                    <SPLIT distance="125" swimtime="00:01:59.56" />
                    <SPLIT distance="150" swimtime="00:02:25.77" />
                    <SPLIT distance="175" swimtime="00:02:48.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="245" reactiontime="+106" swimtime="00:01:30.51" resultid="106426" heatid="110692" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.95" />
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="75" swimtime="00:01:09.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="245" reactiontime="+87" swimtime="00:06:54.14" resultid="106427" heatid="110786" lane="3" entrytime="00:06:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.39" />
                    <SPLIT distance="50" swimtime="00:00:45.63" />
                    <SPLIT distance="75" swimtime="00:01:12.11" />
                    <SPLIT distance="100" swimtime="00:01:40.27" />
                    <SPLIT distance="125" swimtime="00:02:07.95" />
                    <SPLIT distance="150" swimtime="00:02:34.59" />
                    <SPLIT distance="175" swimtime="00:03:01.12" />
                    <SPLIT distance="200" swimtime="00:03:28.18" />
                    <SPLIT distance="225" swimtime="00:03:55.97" />
                    <SPLIT distance="250" swimtime="00:04:23.89" />
                    <SPLIT distance="275" swimtime="00:04:51.85" />
                    <SPLIT distance="300" swimtime="00:05:20.11" />
                    <SPLIT distance="325" swimtime="00:05:44.25" />
                    <SPLIT distance="350" swimtime="00:06:08.94" />
                    <SPLIT distance="375" swimtime="00:06:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="226" swimtime="00:00:47.22" resultid="106428" heatid="110819" lane="6" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-09-09" firstname="VALENTINA" gender="F" lastname="GORODULINA" nation="RUS" athleteid="106418">
              <RESULTS>
                <RESULT eventid="98777" points="231" reactiontime="+86" swimtime="00:00:37.87" resultid="106433" heatid="110589" lane="6" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="238" reactiontime="+107" swimtime="00:12:52.73" resultid="106434" heatid="110634" lane="3" entrytime="00:13:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.35" />
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="75" swimtime="00:01:02.25" />
                    <SPLIT distance="100" swimtime="00:01:25.25" />
                    <SPLIT distance="125" swimtime="00:01:49.16" />
                    <SPLIT distance="150" swimtime="00:02:12.90" />
                    <SPLIT distance="175" swimtime="00:02:37.60" />
                    <SPLIT distance="200" swimtime="00:03:01.68" />
                    <SPLIT distance="225" swimtime="00:03:26.58" />
                    <SPLIT distance="250" swimtime="00:03:50.78" />
                    <SPLIT distance="275" swimtime="00:04:15.61" />
                    <SPLIT distance="300" swimtime="00:04:40.31" />
                    <SPLIT distance="325" swimtime="00:05:05.17" />
                    <SPLIT distance="350" swimtime="00:05:29.52" />
                    <SPLIT distance="375" swimtime="00:05:54.65" />
                    <SPLIT distance="400" swimtime="00:06:18.92" />
                    <SPLIT distance="425" swimtime="00:06:44.03" />
                    <SPLIT distance="450" swimtime="00:07:08.09" />
                    <SPLIT distance="475" swimtime="00:07:32.73" />
                    <SPLIT distance="500" swimtime="00:07:56.84" />
                    <SPLIT distance="525" swimtime="00:08:21.75" />
                    <SPLIT distance="550" swimtime="00:08:46.34" />
                    <SPLIT distance="575" swimtime="00:09:10.94" />
                    <SPLIT distance="600" swimtime="00:09:35.72" />
                    <SPLIT distance="625" swimtime="00:09:59.98" />
                    <SPLIT distance="650" swimtime="00:11:14.35" />
                    <SPLIT distance="675" swimtime="00:10:50.08" />
                    <SPLIT distance="700" swimtime="00:12:04.17" />
                    <SPLIT distance="725" swimtime="00:11:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="234" swimtime="00:01:22.53" resultid="106435" heatid="110674" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="75" swimtime="00:01:01.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="253" swimtime="00:02:55.06" resultid="106436" heatid="110765" lane="4" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.05" />
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                    <SPLIT distance="75" swimtime="00:01:01.35" />
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="125" swimtime="00:01:47.13" />
                    <SPLIT distance="150" swimtime="00:02:10.09" />
                    <SPLIT distance="175" swimtime="00:02:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="241" swimtime="00:06:16.55" resultid="106437" heatid="110841" lane="0" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                    <SPLIT distance="75" swimtime="00:01:02.71" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="125" swimtime="00:01:49.76" />
                    <SPLIT distance="150" swimtime="00:02:13.67" />
                    <SPLIT distance="175" swimtime="00:02:37.57" />
                    <SPLIT distance="200" swimtime="00:03:02.42" />
                    <SPLIT distance="225" swimtime="00:03:26.70" />
                    <SPLIT distance="250" swimtime="00:03:51.08" />
                    <SPLIT distance="275" swimtime="00:04:15.65" />
                    <SPLIT distance="300" swimtime="00:04:39.57" />
                    <SPLIT distance="325" swimtime="00:05:03.65" />
                    <SPLIT distance="350" swimtime="00:05:27.82" />
                    <SPLIT distance="375" swimtime="00:05:52.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="109627" name="AQUASFERA Masters Olsztyn">
          <CONTACT email="annamariaaneczka@gmail.com" name="Goździejewska" />
          <ATHLETES>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="109925">
              <RESULTS>
                <RESULT eventid="98777" points="393" reactiontime="+92" swimtime="00:00:31.71" resultid="109926" heatid="110591" lane="3" entrytime="00:00:31.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="321" reactiontime="+75" swimtime="00:02:57.97" resultid="109927" heatid="110617" lane="7" entrytime="00:02:57.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.82" />
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="75" swimtime="00:01:00.19" />
                    <SPLIT distance="100" swimtime="00:01:22.48" />
                    <SPLIT distance="125" swimtime="00:01:50.34" />
                    <SPLIT distance="150" swimtime="00:02:17.75" />
                    <SPLIT distance="175" swimtime="00:02:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="339" reactiontime="+80" swimtime="00:00:36.79" resultid="109928" heatid="110649" lane="7" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="349" swimtime="00:01:20.43" resultid="109929" heatid="110694" lane="0" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.52" />
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="75" swimtime="00:01:01.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="303" reactiontime="+80" swimtime="00:01:21.93" resultid="109930" heatid="110755" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.10" />
                    <SPLIT distance="50" swimtime="00:00:39.63" />
                    <SPLIT distance="75" swimtime="00:01:01.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="295" reactiontime="+77" swimtime="00:02:58.92" resultid="109931" heatid="110809" lane="9" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.63" />
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="75" swimtime="00:01:03.35" />
                    <SPLIT distance="100" swimtime="00:01:26.40" />
                    <SPLIT distance="125" swimtime="00:01:50.01" />
                    <SPLIT distance="150" swimtime="00:02:13.62" />
                    <SPLIT distance="175" swimtime="00:02:36.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-16" firstname="Krzysztof" gender="M" lastname="Sopyła" nation="POL" athleteid="109818">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="109819" heatid="110600" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="109820" heatid="110680" lane="2" entrytime="00:01:22.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="Zaleska" nation="POL" athleteid="109985">
              <RESULTS>
                <RESULT eventid="98814" points="427" reactiontime="+65" swimtime="00:02:41.81" resultid="109986" heatid="110615" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.39" />
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="75" swimtime="00:00:55.07" />
                    <SPLIT distance="100" swimtime="00:01:15.65" />
                    <SPLIT distance="125" swimtime="00:01:39.58" />
                    <SPLIT distance="150" swimtime="00:02:03.24" />
                    <SPLIT distance="175" swimtime="00:02:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="413" swimtime="00:10:43.17" resultid="109987" heatid="110633" lane="6" entrytime="00:11:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.28" />
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="75" swimtime="00:00:55.41" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="125" swimtime="00:01:35.31" />
                    <SPLIT distance="150" swimtime="00:01:55.63" />
                    <SPLIT distance="175" swimtime="00:02:15.91" />
                    <SPLIT distance="200" swimtime="00:02:36.13" />
                    <SPLIT distance="225" swimtime="00:02:56.39" />
                    <SPLIT distance="250" swimtime="00:03:16.79" />
                    <SPLIT distance="275" swimtime="00:03:36.99" />
                    <SPLIT distance="300" swimtime="00:03:57.48" />
                    <SPLIT distance="325" swimtime="00:04:17.86" />
                    <SPLIT distance="350" swimtime="00:04:38.49" />
                    <SPLIT distance="375" swimtime="00:04:59.08" />
                    <SPLIT distance="400" swimtime="00:05:20.01" />
                    <SPLIT distance="425" swimtime="00:05:40.39" />
                    <SPLIT distance="450" swimtime="00:06:01.02" />
                    <SPLIT distance="475" swimtime="00:06:21.74" />
                    <SPLIT distance="500" swimtime="00:06:42.78" />
                    <SPLIT distance="525" swimtime="00:07:02.95" />
                    <SPLIT distance="550" swimtime="00:07:23.37" />
                    <SPLIT distance="575" swimtime="00:07:43.42" />
                    <SPLIT distance="600" swimtime="00:08:04.34" />
                    <SPLIT distance="625" swimtime="00:08:24.60" />
                    <SPLIT distance="650" swimtime="00:08:45.33" />
                    <SPLIT distance="675" swimtime="00:09:05.81" />
                    <SPLIT distance="700" swimtime="00:09:26.45" />
                    <SPLIT distance="725" swimtime="00:09:45.30" />
                    <SPLIT distance="750" swimtime="00:10:04.93" />
                    <SPLIT distance="775" swimtime="00:10:24.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="311" reactiontime="+80" swimtime="00:03:18.50" resultid="109988" heatid="110663" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.92" />
                    <SPLIT distance="50" swimtime="00:00:45.09" />
                    <SPLIT distance="75" swimtime="00:01:10.08" />
                    <SPLIT distance="100" swimtime="00:01:35.50" />
                    <SPLIT distance="125" swimtime="00:02:00.75" />
                    <SPLIT distance="150" swimtime="00:02:26.89" />
                    <SPLIT distance="175" swimtime="00:02:52.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="435" reactiontime="+68" swimtime="00:02:37.80" resultid="109989" heatid="110708" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.97" />
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="75" swimtime="00:00:54.77" />
                    <SPLIT distance="100" swimtime="00:01:14.76" />
                    <SPLIT distance="125" swimtime="00:01:35.11" />
                    <SPLIT distance="150" swimtime="00:01:55.86" />
                    <SPLIT distance="175" swimtime="00:02:16.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="416" reactiontime="+70" swimtime="00:00:32.64" resultid="109990" heatid="110739" lane="7" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="424" reactiontime="+71" swimtime="00:05:45.22" resultid="109991" heatid="110787" lane="7" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.27" />
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="75" swimtime="00:00:55.77" />
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="125" swimtime="00:01:40.29" />
                    <SPLIT distance="150" swimtime="00:02:02.90" />
                    <SPLIT distance="175" swimtime="00:02:25.85" />
                    <SPLIT distance="200" swimtime="00:02:48.33" />
                    <SPLIT distance="225" swimtime="00:03:13.50" />
                    <SPLIT distance="250" swimtime="00:03:38.28" />
                    <SPLIT distance="275" swimtime="00:04:03.22" />
                    <SPLIT distance="300" swimtime="00:04:28.09" />
                    <SPLIT distance="325" swimtime="00:04:48.28" />
                    <SPLIT distance="350" swimtime="00:05:07.87" />
                    <SPLIT distance="375" swimtime="00:05:27.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="424" reactiontime="+80" swimtime="00:01:12.65" resultid="109992" heatid="110796" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.98" />
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="75" swimtime="00:00:53.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="412" reactiontime="+99" swimtime="00:05:15.05" resultid="109993" heatid="110840" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.49" />
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="75" swimtime="00:00:56.74" />
                    <SPLIT distance="100" swimtime="00:01:16.63" />
                    <SPLIT distance="125" swimtime="00:01:36.66" />
                    <SPLIT distance="150" swimtime="00:01:56.61" />
                    <SPLIT distance="175" swimtime="00:02:16.90" />
                    <SPLIT distance="200" swimtime="00:02:37.23" />
                    <SPLIT distance="225" swimtime="00:02:57.40" />
                    <SPLIT distance="250" swimtime="00:03:17.51" />
                    <SPLIT distance="275" swimtime="00:03:37.78" />
                    <SPLIT distance="300" swimtime="00:03:58.13" />
                    <SPLIT distance="325" swimtime="00:04:17.97" />
                    <SPLIT distance="350" swimtime="00:04:38.20" />
                    <SPLIT distance="375" swimtime="00:04:57.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-25" firstname="Adam" gender="M" lastname="Matusiak vel Matuszewski" nation="POL" athleteid="109958">
              <RESULTS>
                <RESULT eventid="98798" points="191" reactiontime="+75" swimtime="00:00:35.12" resultid="109959" heatid="110595" lane="8">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="181" reactiontime="+75" swimtime="00:01:19.34" resultid="109960" heatid="110678" lane="8">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.40" />
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="75" swimtime="00:00:59.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="131" swimtime="00:00:42.87" resultid="109961" heatid="110741" lane="6">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="171" reactiontime="+89" swimtime="00:02:58.82" resultid="109962" heatid="110769" lane="7">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.49" />
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                    <SPLIT distance="75" swimtime="00:01:03.42" />
                    <SPLIT distance="100" swimtime="00:01:26.97" />
                    <SPLIT distance="125" swimtime="00:01:51.37" />
                    <SPLIT distance="150" swimtime="00:02:14.96" />
                    <SPLIT distance="175" swimtime="00:02:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="160" reactiontime="+99" swimtime="00:06:30.18" resultid="109963" heatid="110852" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.43" />
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                    <SPLIT distance="75" swimtime="00:01:09.47" />
                    <SPLIT distance="100" swimtime="00:01:34.62" />
                    <SPLIT distance="125" swimtime="00:02:00.60" />
                    <SPLIT distance="150" swimtime="00:02:25.96" />
                    <SPLIT distance="175" swimtime="00:02:51.29" />
                    <SPLIT distance="200" swimtime="00:03:16.27" />
                    <SPLIT distance="225" swimtime="00:03:41.57" />
                    <SPLIT distance="250" swimtime="00:04:06.47" />
                    <SPLIT distance="275" swimtime="00:04:31.30" />
                    <SPLIT distance="300" swimtime="00:04:56.58" />
                    <SPLIT distance="325" swimtime="00:05:21.31" />
                    <SPLIT distance="350" swimtime="00:05:46.13" />
                    <SPLIT distance="375" swimtime="00:06:09.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-08-31" firstname="Iwona" gender="F" lastname="Bardzicka" nation="POL" athleteid="109907">
              <RESULTS>
                <RESULT eventid="98940" points="106" swimtime="00:04:43.79" resultid="109908" heatid="110661" lane="2" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.24" />
                    <SPLIT distance="50" swimtime="00:01:05.26" />
                    <SPLIT distance="75" swimtime="00:01:40.83" />
                    <SPLIT distance="100" swimtime="00:02:16.61" />
                    <SPLIT distance="125" swimtime="00:02:53.90" />
                    <SPLIT distance="150" swimtime="00:03:31.07" />
                    <SPLIT distance="175" swimtime="00:04:07.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="111" swimtime="00:02:09.69" resultid="109909" heatid="110721" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.66" />
                    <SPLIT distance="50" swimtime="00:01:03.28" />
                    <SPLIT distance="75" swimtime="00:01:36.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="121" swimtime="00:00:58.22" resultid="109910" heatid="110818" lane="8" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-16" firstname="Paweł" gender="M" lastname="Szczuka" nation="POL" athleteid="109900">
              <RESULTS>
                <RESULT eventid="98830" points="448" reactiontime="+80" swimtime="00:02:23.22" resultid="109901" heatid="110627" lane="3" entrytime="00:02:28.28">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="75" swimtime="00:00:48.63" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="125" swimtime="00:01:27.00" />
                    <SPLIT distance="150" swimtime="00:01:48.09" />
                    <SPLIT distance="175" swimtime="00:02:05.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="375" reactiontime="+85" swimtime="00:00:30.81" resultid="109902" heatid="110651" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="480" reactiontime="+73" swimtime="00:01:04.68" resultid="109903" heatid="110705" lane="8" entrytime="00:01:06.66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.06" />
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                    <SPLIT distance="75" swimtime="00:00:48.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="378" reactiontime="+88" swimtime="00:01:07.64" resultid="109904" heatid="110757" lane="7">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.69" />
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="75" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="450" swimtime="00:05:07.15" resultid="109905" heatid="110792" lane="0" entrytime="00:05:26.28">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.98" />
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="75" swimtime="00:00:48.62" />
                    <SPLIT distance="100" swimtime="00:01:07.16" />
                    <SPLIT distance="125" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:01:47.26" />
                    <SPLIT distance="175" swimtime="00:02:07.49" />
                    <SPLIT distance="200" swimtime="00:02:27.42" />
                    <SPLIT distance="225" swimtime="00:02:48.93" />
                    <SPLIT distance="250" swimtime="00:03:11.05" />
                    <SPLIT distance="275" swimtime="00:03:33.04" />
                    <SPLIT distance="300" swimtime="00:03:56.13" />
                    <SPLIT distance="325" swimtime="00:04:14.08" />
                    <SPLIT distance="350" swimtime="00:04:31.76" />
                    <SPLIT distance="375" swimtime="00:04:49.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="442" reactiontime="+64" swimtime="00:01:03.56" resultid="109906" heatid="110797" lane="4">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                    <SPLIT distance="75" swimtime="00:00:45.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-14" firstname="Wojciech" gender="M" lastname="Kłujszo" nation="POL" athleteid="109841">
              <RESULTS>
                <RESULT eventid="98798" points="288" reactiontime="+63" swimtime="00:00:30.67" resultid="109842" heatid="110594" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="257" reactiontime="+88" swimtime="00:00:39.67" resultid="109843" heatid="110824" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-02-28" firstname="Dawid" gender="M" lastname="Zieja" nation="POL" athleteid="109887">
              <RESULTS>
                <RESULT eventid="98798" points="535" reactiontime="+89" swimtime="00:00:24.95" resultid="109888" heatid="110613" lane="2" entrytime="00:00:23.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="404" reactiontime="+74" swimtime="00:09:59.46" resultid="109889" heatid="110635" lane="6" entrytime="00:09:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="75" swimtime="00:00:50.11" />
                    <SPLIT distance="100" swimtime="00:01:08.61" />
                    <SPLIT distance="125" swimtime="00:01:27.19" />
                    <SPLIT distance="150" swimtime="00:01:45.93" />
                    <SPLIT distance="175" swimtime="00:02:04.91" />
                    <SPLIT distance="200" swimtime="00:02:23.83" />
                    <SPLIT distance="225" swimtime="00:02:42.68" />
                    <SPLIT distance="250" swimtime="00:03:01.57" />
                    <SPLIT distance="275" swimtime="00:03:20.33" />
                    <SPLIT distance="300" swimtime="00:03:39.45" />
                    <SPLIT distance="325" swimtime="00:03:58.21" />
                    <SPLIT distance="350" swimtime="00:04:17.28" />
                    <SPLIT distance="375" swimtime="00:04:36.06" />
                    <SPLIT distance="400" swimtime="00:04:55.04" />
                    <SPLIT distance="425" swimtime="00:05:13.64" />
                    <SPLIT distance="450" swimtime="00:05:32.54" />
                    <SPLIT distance="475" swimtime="00:05:51.60" />
                    <SPLIT distance="500" swimtime="00:06:10.95" />
                    <SPLIT distance="525" swimtime="00:06:29.93" />
                    <SPLIT distance="550" swimtime="00:06:49.32" />
                    <SPLIT distance="575" swimtime="00:07:09.03" />
                    <SPLIT distance="600" swimtime="00:07:28.09" />
                    <SPLIT distance="625" swimtime="00:07:47.42" />
                    <SPLIT distance="650" swimtime="00:08:06.76" />
                    <SPLIT distance="675" swimtime="00:08:26.47" />
                    <SPLIT distance="700" swimtime="00:08:45.83" />
                    <SPLIT distance="725" swimtime="00:09:04.68" />
                    <SPLIT distance="750" swimtime="00:09:24.07" />
                    <SPLIT distance="775" swimtime="00:09:42.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="577" reactiontime="+74" swimtime="00:01:59.34" resultid="109890" heatid="110778" lane="5" entrytime="00:01:56.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.64" />
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                    <SPLIT distance="75" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:00:57.48" />
                    <SPLIT distance="125" swimtime="00:01:13.02" />
                    <SPLIT distance="150" swimtime="00:01:28.67" />
                    <SPLIT distance="175" swimtime="00:01:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="561" reactiontime="+64" swimtime="00:00:58.71" resultid="109891" heatid="110805" lane="7" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.67" />
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="75" swimtime="00:00:42.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="468" swimtime="00:04:33.19" resultid="109892" heatid="110843" lane="9" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.88" />
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="75" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:03.97" />
                    <SPLIT distance="125" swimtime="00:01:20.97" />
                    <SPLIT distance="150" swimtime="00:01:38.64" />
                    <SPLIT distance="175" swimtime="00:01:56.08" />
                    <SPLIT distance="200" swimtime="00:02:13.87" />
                    <SPLIT distance="225" swimtime="00:02:31.36" />
                    <SPLIT distance="250" swimtime="00:02:49.03" />
                    <SPLIT distance="275" swimtime="00:03:06.48" />
                    <SPLIT distance="300" swimtime="00:03:24.01" />
                    <SPLIT distance="325" swimtime="00:03:41.40" />
                    <SPLIT distance="350" swimtime="00:03:59.03" />
                    <SPLIT distance="375" swimtime="00:04:16.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-09" firstname="Marek" gender="M" lastname="Koźlikowski" nation="POL" athleteid="109853">
              <RESULTS>
                <RESULT eventid="98830" points="237" reactiontime="+90" swimtime="00:02:56.95" resultid="109854" heatid="110622" lane="8" entrytime="00:03:08.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.39" />
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="75" swimtime="00:01:02.12" />
                    <SPLIT distance="100" swimtime="00:01:27.81" />
                    <SPLIT distance="125" swimtime="00:01:51.53" />
                    <SPLIT distance="150" swimtime="00:02:16.46" />
                    <SPLIT distance="175" swimtime="00:02:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="219" reactiontime="+102" swimtime="00:23:26.79" resultid="109855" heatid="110643" lane="4" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.54" />
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                    <SPLIT distance="75" swimtime="00:01:05.18" />
                    <SPLIT distance="100" swimtime="00:01:28.89" />
                    <SPLIT distance="125" swimtime="00:01:52.82" />
                    <SPLIT distance="150" swimtime="00:02:16.29" />
                    <SPLIT distance="175" swimtime="00:02:40.31" />
                    <SPLIT distance="200" swimtime="00:03:03.77" />
                    <SPLIT distance="225" swimtime="00:03:27.77" />
                    <SPLIT distance="250" swimtime="00:03:51.89" />
                    <SPLIT distance="275" swimtime="00:04:16.44" />
                    <SPLIT distance="300" swimtime="00:04:40.22" />
                    <SPLIT distance="325" swimtime="00:05:04.38" />
                    <SPLIT distance="350" swimtime="00:05:28.52" />
                    <SPLIT distance="375" swimtime="00:05:53.06" />
                    <SPLIT distance="400" swimtime="00:06:16.80" />
                    <SPLIT distance="425" swimtime="00:06:40.82" />
                    <SPLIT distance="450" swimtime="00:07:04.86" />
                    <SPLIT distance="475" swimtime="00:07:29.42" />
                    <SPLIT distance="500" swimtime="00:07:53.37" />
                    <SPLIT distance="525" swimtime="00:08:17.15" />
                    <SPLIT distance="550" swimtime="00:08:41.23" />
                    <SPLIT distance="575" swimtime="00:09:05.18" />
                    <SPLIT distance="600" swimtime="00:09:29.21" />
                    <SPLIT distance="625" swimtime="00:09:53.46" />
                    <SPLIT distance="650" swimtime="00:10:17.25" />
                    <SPLIT distance="675" swimtime="00:10:40.92" />
                    <SPLIT distance="700" swimtime="00:11:04.55" />
                    <SPLIT distance="725" swimtime="00:11:27.87" />
                    <SPLIT distance="750" swimtime="00:11:51.21" />
                    <SPLIT distance="775" swimtime="00:12:14.65" />
                    <SPLIT distance="800" swimtime="00:12:37.79" />
                    <SPLIT distance="825" swimtime="00:13:01.44" />
                    <SPLIT distance="850" swimtime="00:13:24.79" />
                    <SPLIT distance="875" swimtime="00:13:48.47" />
                    <SPLIT distance="900" swimtime="00:14:11.54" />
                    <SPLIT distance="925" swimtime="00:14:34.87" />
                    <SPLIT distance="950" swimtime="00:14:58.31" />
                    <SPLIT distance="975" swimtime="00:15:21.47" />
                    <SPLIT distance="1000" swimtime="00:15:44.75" />
                    <SPLIT distance="1025" swimtime="00:16:08.12" />
                    <SPLIT distance="1050" swimtime="00:16:31.67" />
                    <SPLIT distance="1075" swimtime="00:16:54.89" />
                    <SPLIT distance="1100" swimtime="00:17:18.27" />
                    <SPLIT distance="1125" swimtime="00:17:41.74" />
                    <SPLIT distance="1150" swimtime="00:18:05.07" />
                    <SPLIT distance="1175" swimtime="00:18:28.82" />
                    <SPLIT distance="1200" swimtime="00:18:52.07" />
                    <SPLIT distance="1225" swimtime="00:19:15.65" />
                    <SPLIT distance="1250" swimtime="00:19:38.51" />
                    <SPLIT distance="1275" swimtime="00:20:01.84" />
                    <SPLIT distance="1300" swimtime="00:20:24.87" />
                    <SPLIT distance="1325" swimtime="00:20:48.25" />
                    <SPLIT distance="1350" swimtime="00:21:11.59" />
                    <SPLIT distance="1375" swimtime="00:21:34.22" />
                    <SPLIT distance="1400" swimtime="00:21:56.89" />
                    <SPLIT distance="1425" swimtime="00:22:19.63" />
                    <SPLIT distance="1450" swimtime="00:22:42.54" />
                    <SPLIT distance="1475" swimtime="00:23:05.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="109856" heatid="110667" lane="0" entrytime="00:03:22.53" />
                <RESULT eventid="98988" points="242" reactiontime="+78" swimtime="00:01:21.26" resultid="109857" heatid="110698" lane="7" entrytime="00:01:25.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.43" />
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="75" swimtime="00:01:02.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="240" reactiontime="+89" swimtime="00:02:39.88" resultid="109858" heatid="110771" lane="8" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.52" />
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="75" swimtime="00:00:57.67" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="125" swimtime="00:01:39.78" />
                    <SPLIT distance="150" swimtime="00:02:00.44" />
                    <SPLIT distance="175" swimtime="00:02:21.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="208" reactiontime="+107" swimtime="00:06:37.41" resultid="109859" heatid="110789" lane="1" entrytime="00:06:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.02" />
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="75" swimtime="00:01:07.50" />
                    <SPLIT distance="100" swimtime="00:01:34.51" />
                    <SPLIT distance="125" swimtime="00:02:03.01" />
                    <SPLIT distance="150" swimtime="00:02:31.05" />
                    <SPLIT distance="175" swimtime="00:02:58.03" />
                    <SPLIT distance="200" swimtime="00:03:25.36" />
                    <SPLIT distance="225" swimtime="00:03:51.53" />
                    <SPLIT distance="250" swimtime="00:04:18.08" />
                    <SPLIT distance="275" swimtime="00:04:44.10" />
                    <SPLIT distance="300" swimtime="00:05:10.76" />
                    <SPLIT distance="325" swimtime="00:05:33.16" />
                    <SPLIT distance="350" swimtime="00:05:55.52" />
                    <SPLIT distance="375" swimtime="00:06:16.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="180" reactiontime="+87" swimtime="00:01:25.69" resultid="109860" heatid="110800" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.80" />
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="75" swimtime="00:01:01.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="231" swimtime="00:05:45.79" resultid="109861" heatid="110848" lane="0" entrytime="00:05:59.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.09" />
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="75" swimtime="00:00:58.31" />
                    <SPLIT distance="100" swimtime="00:01:19.52" />
                    <SPLIT distance="125" swimtime="00:01:41.22" />
                    <SPLIT distance="150" swimtime="00:02:03.51" />
                    <SPLIT distance="175" swimtime="00:02:26.04" />
                    <SPLIT distance="200" swimtime="00:02:48.15" />
                    <SPLIT distance="225" swimtime="00:03:10.86" />
                    <SPLIT distance="250" swimtime="00:03:33.12" />
                    <SPLIT distance="275" swimtime="00:03:55.81" />
                    <SPLIT distance="300" swimtime="00:04:18.31" />
                    <SPLIT distance="325" swimtime="00:04:40.67" />
                    <SPLIT distance="350" swimtime="00:05:03.02" />
                    <SPLIT distance="375" swimtime="00:05:25.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-03-29" firstname="Jarosław" gender="M" lastname="Szczepanik" nation="POL" athleteid="109939">
              <RESULTS>
                <RESULT eventid="98798" points="321" reactiontime="+93" swimtime="00:00:29.57" resultid="109940" heatid="110594" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="291" reactiontime="+55" swimtime="00:01:16.44" resultid="109941" heatid="110696" lane="2">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.06" />
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="75" swimtime="00:00:56.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-25" firstname="Piotr" gender="M" lastname="Markowicz" nation="POL" athleteid="109942">
              <RESULTS>
                <RESULT eventid="98798" points="321" reactiontime="+88" swimtime="00:00:29.56" resultid="109943" heatid="110603" lane="3" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="326" reactiontime="+107" swimtime="00:10:43.84" resultid="109944" heatid="110636" lane="0" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.45" />
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="75" swimtime="00:00:55.81" />
                    <SPLIT distance="100" swimtime="00:01:15.47" />
                    <SPLIT distance="125" swimtime="00:01:35.67" />
                    <SPLIT distance="150" swimtime="00:01:55.82" />
                    <SPLIT distance="175" swimtime="00:02:16.30" />
                    <SPLIT distance="200" swimtime="00:02:37.11" />
                    <SPLIT distance="225" swimtime="00:02:57.87" />
                    <SPLIT distance="250" swimtime="00:03:18.52" />
                    <SPLIT distance="275" swimtime="00:03:38.91" />
                    <SPLIT distance="300" swimtime="00:03:59.60" />
                    <SPLIT distance="325" swimtime="00:04:20.03" />
                    <SPLIT distance="350" swimtime="00:04:40.39" />
                    <SPLIT distance="375" swimtime="00:05:00.37" />
                    <SPLIT distance="400" swimtime="00:05:20.41" />
                    <SPLIT distance="425" swimtime="00:05:40.63" />
                    <SPLIT distance="450" swimtime="00:06:00.66" />
                    <SPLIT distance="475" swimtime="00:06:21.15" />
                    <SPLIT distance="500" swimtime="00:06:41.59" />
                    <SPLIT distance="525" swimtime="00:07:01.56" />
                    <SPLIT distance="550" swimtime="00:07:21.73" />
                    <SPLIT distance="575" swimtime="00:07:42.02" />
                    <SPLIT distance="600" swimtime="00:08:02.31" />
                    <SPLIT distance="625" swimtime="00:08:22.31" />
                    <SPLIT distance="650" swimtime="00:08:42.78" />
                    <SPLIT distance="675" swimtime="00:09:03.13" />
                    <SPLIT distance="700" swimtime="00:09:23.72" />
                    <SPLIT distance="725" swimtime="00:09:43.83" />
                    <SPLIT distance="750" swimtime="00:10:04.54" />
                    <SPLIT distance="775" swimtime="00:10:24.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="252" reactiontime="+90" swimtime="00:00:35.14" resultid="109945" heatid="110656" lane="0" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="305" reactiontime="+91" swimtime="00:01:15.19" resultid="109946" heatid="110701" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.36" />
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="75" swimtime="00:00:56.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="306" swimtime="00:00:32.34" resultid="109947" heatid="110744" lane="6" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="256" reactiontime="+85" swimtime="00:06:10.66" resultid="109948" heatid="110790" lane="7" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.62" />
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="75" swimtime="00:00:57.81" />
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                    <SPLIT distance="125" swimtime="00:01:43.68" />
                    <SPLIT distance="150" swimtime="00:02:06.86" />
                    <SPLIT distance="175" swimtime="00:02:30.58" />
                    <SPLIT distance="200" swimtime="00:02:54.09" />
                    <SPLIT distance="225" swimtime="00:03:21.70" />
                    <SPLIT distance="250" swimtime="00:03:49.04" />
                    <SPLIT distance="275" swimtime="00:04:16.51" />
                    <SPLIT distance="300" swimtime="00:04:44.36" />
                    <SPLIT distance="325" swimtime="00:05:07.03" />
                    <SPLIT distance="350" swimtime="00:05:29.19" />
                    <SPLIT distance="375" swimtime="00:05:50.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="109949" heatid="110813" lane="3" entrytime="00:02:55.00" />
                <RESULT eventid="99473" points="317" reactiontime="+84" swimtime="00:05:11.11" resultid="109950" heatid="110846" lane="7" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.29" />
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="75" swimtime="00:00:54.61" />
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                    <SPLIT distance="125" swimtime="00:01:32.93" />
                    <SPLIT distance="150" swimtime="00:01:52.16" />
                    <SPLIT distance="175" swimtime="00:02:11.57" />
                    <SPLIT distance="200" swimtime="00:02:31.42" />
                    <SPLIT distance="225" swimtime="00:02:51.36" />
                    <SPLIT distance="250" swimtime="00:03:11.11" />
                    <SPLIT distance="275" swimtime="00:03:31.20" />
                    <SPLIT distance="300" swimtime="00:03:51.41" />
                    <SPLIT distance="325" swimtime="00:04:11.91" />
                    <SPLIT distance="350" swimtime="00:04:31.84" />
                    <SPLIT distance="375" swimtime="00:04:51.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="109844">
              <RESULTS>
                <RESULT eventid="98798" points="328" reactiontime="+92" swimtime="00:00:29.37" resultid="109845" heatid="110607" lane="0" entrytime="00:00:28.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="349" reactiontime="+72" swimtime="00:10:29.77" resultid="109846" heatid="110635" lane="7" entrytime="00:10:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.67" />
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="75" swimtime="00:00:54.30" />
                    <SPLIT distance="100" swimtime="00:01:13.58" />
                    <SPLIT distance="125" swimtime="00:01:32.71" />
                    <SPLIT distance="150" swimtime="00:01:52.42" />
                    <SPLIT distance="175" swimtime="00:02:11.66" />
                    <SPLIT distance="200" swimtime="00:02:31.40" />
                    <SPLIT distance="225" swimtime="00:02:50.91" />
                    <SPLIT distance="250" swimtime="00:03:10.61" />
                    <SPLIT distance="275" swimtime="00:03:30.31" />
                    <SPLIT distance="300" swimtime="00:03:50.02" />
                    <SPLIT distance="325" swimtime="00:04:09.72" />
                    <SPLIT distance="350" swimtime="00:04:29.90" />
                    <SPLIT distance="375" swimtime="00:04:49.68" />
                    <SPLIT distance="400" swimtime="00:05:09.71" />
                    <SPLIT distance="425" swimtime="00:05:29.38" />
                    <SPLIT distance="450" swimtime="00:05:49.52" />
                    <SPLIT distance="475" swimtime="00:06:09.44" />
                    <SPLIT distance="500" swimtime="00:06:29.42" />
                    <SPLIT distance="525" swimtime="00:06:49.37" />
                    <SPLIT distance="550" swimtime="00:07:09.68" />
                    <SPLIT distance="575" swimtime="00:07:29.38" />
                    <SPLIT distance="600" swimtime="00:07:49.51" />
                    <SPLIT distance="625" swimtime="00:08:09.51" />
                    <SPLIT distance="650" swimtime="00:08:29.87" />
                    <SPLIT distance="675" swimtime="00:08:49.97" />
                    <SPLIT distance="700" swimtime="00:09:10.17" />
                    <SPLIT distance="725" swimtime="00:09:30.31" />
                    <SPLIT distance="750" swimtime="00:09:50.51" />
                    <SPLIT distance="775" swimtime="00:10:10.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="289" reactiontime="+86" swimtime="00:00:33.59" resultid="109847" heatid="110657" lane="5" entrytime="00:00:33.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="254" reactiontime="+86" swimtime="00:02:51.20" resultid="109848" heatid="110713" lane="8" entrytime="00:02:38.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.91" />
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="75" swimtime="00:00:56.68" />
                    <SPLIT distance="100" swimtime="00:01:17.75" />
                    <SPLIT distance="125" swimtime="00:01:39.43" />
                    <SPLIT distance="150" swimtime="00:02:01.57" />
                    <SPLIT distance="175" swimtime="00:02:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="347" reactiontime="+92" swimtime="00:00:31.02" resultid="109849" heatid="110746" lane="1" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="335" swimtime="00:02:23.04" resultid="109850" heatid="110776" lane="0" entrytime="00:02:18.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.23" />
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="75" swimtime="00:00:53.28" />
                    <SPLIT distance="100" swimtime="00:01:11.56" />
                    <SPLIT distance="125" swimtime="00:01:29.64" />
                    <SPLIT distance="150" swimtime="00:01:47.81" />
                    <SPLIT distance="175" swimtime="00:02:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="329" swimtime="00:01:10.15" resultid="109851" heatid="110803" lane="6" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.94" />
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="75" swimtime="00:00:50.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="339" reactiontime="+89" swimtime="00:05:04.22" resultid="109852" heatid="110844" lane="1" entrytime="00:04:49.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.66" />
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="75" swimtime="00:00:54.14" />
                    <SPLIT distance="100" swimtime="00:01:13.35" />
                    <SPLIT distance="125" swimtime="00:01:32.49" />
                    <SPLIT distance="150" swimtime="00:01:51.47" />
                    <SPLIT distance="175" swimtime="00:02:10.85" />
                    <SPLIT distance="200" swimtime="00:02:30.12" />
                    <SPLIT distance="225" swimtime="00:02:49.27" />
                    <SPLIT distance="250" swimtime="00:03:08.67" />
                    <SPLIT distance="275" swimtime="00:03:28.06" />
                    <SPLIT distance="300" swimtime="00:03:47.48" />
                    <SPLIT distance="325" swimtime="00:04:06.84" />
                    <SPLIT distance="350" swimtime="00:04:26.27" />
                    <SPLIT distance="375" swimtime="00:04:45.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-13" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="109951">
              <RESULTS>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="109952" heatid="110623" lane="5" entrytime="00:02:50.00" />
                <RESULT eventid="98956" points="455" reactiontime="+77" swimtime="00:02:36.57" resultid="109953" heatid="110669" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="75" swimtime="00:00:54.78" />
                    <SPLIT distance="100" swimtime="00:01:14.70" />
                    <SPLIT distance="125" swimtime="00:01:34.92" />
                    <SPLIT distance="150" swimtime="00:01:55.33" />
                    <SPLIT distance="175" swimtime="00:02:15.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="418" reactiontime="+64" swimtime="00:01:07.71" resultid="109954" heatid="110704" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="75" swimtime="00:00:51.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="487" reactiontime="+67" swimtime="00:01:10.66" resultid="109955" heatid="110733" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.41" />
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="75" swimtime="00:00:52.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="362" reactiontime="+76" swimtime="00:05:30.17" resultid="109956" heatid="110791" lane="8" entrytime="00:05:55.06">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="75" swimtime="00:00:57.60" />
                    <SPLIT distance="100" swimtime="00:01:19.75" />
                    <SPLIT distance="125" swimtime="00:01:41.61" />
                    <SPLIT distance="150" swimtime="00:02:02.86" />
                    <SPLIT distance="175" swimtime="00:02:23.90" />
                    <SPLIT distance="200" swimtime="00:02:44.17" />
                    <SPLIT distance="225" swimtime="00:03:05.95" />
                    <SPLIT distance="250" swimtime="00:03:27.45" />
                    <SPLIT distance="275" swimtime="00:03:49.03" />
                    <SPLIT distance="300" swimtime="00:04:10.95" />
                    <SPLIT distance="325" swimtime="00:04:31.78" />
                    <SPLIT distance="350" swimtime="00:04:51.46" />
                    <SPLIT distance="375" swimtime="00:05:12.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="491" reactiontime="+79" swimtime="00:00:32.00" resultid="109957" heatid="110833" lane="3" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-01" firstname="Małgorzata" gender="F" lastname="Polito" nation="POL" athleteid="109920">
              <RESULTS>
                <RESULT eventid="98863" points="299" reactiontime="+93" swimtime="00:11:56.59" resultid="109921" heatid="110633" lane="1" entrytime="00:11:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.20" />
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="75" swimtime="00:01:00.04" />
                    <SPLIT distance="100" swimtime="00:01:21.79" />
                    <SPLIT distance="125" swimtime="00:01:43.70" />
                    <SPLIT distance="150" swimtime="00:02:06.18" />
                    <SPLIT distance="175" swimtime="00:02:28.68" />
                    <SPLIT distance="200" swimtime="00:02:51.24" />
                    <SPLIT distance="225" swimtime="00:03:13.98" />
                    <SPLIT distance="250" swimtime="00:03:36.78" />
                    <SPLIT distance="275" swimtime="00:03:59.52" />
                    <SPLIT distance="300" swimtime="00:04:22.33" />
                    <SPLIT distance="325" swimtime="00:04:45.15" />
                    <SPLIT distance="350" swimtime="00:05:07.72" />
                    <SPLIT distance="375" swimtime="00:05:30.49" />
                    <SPLIT distance="400" swimtime="00:05:53.35" />
                    <SPLIT distance="425" swimtime="00:06:16.26" />
                    <SPLIT distance="450" swimtime="00:06:38.97" />
                    <SPLIT distance="475" swimtime="00:07:01.63" />
                    <SPLIT distance="500" swimtime="00:07:24.36" />
                    <SPLIT distance="525" swimtime="00:07:47.08" />
                    <SPLIT distance="550" swimtime="00:08:09.89" />
                    <SPLIT distance="575" swimtime="00:08:32.54" />
                    <SPLIT distance="600" swimtime="00:08:55.55" />
                    <SPLIT distance="625" swimtime="00:09:18.56" />
                    <SPLIT distance="650" swimtime="00:09:41.49" />
                    <SPLIT distance="675" swimtime="00:10:04.27" />
                    <SPLIT distance="700" swimtime="00:10:27.17" />
                    <SPLIT distance="725" swimtime="00:10:50.28" />
                    <SPLIT distance="750" swimtime="00:11:12.89" />
                    <SPLIT distance="775" swimtime="00:11:35.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="321" swimtime="00:01:31.07" resultid="109922" heatid="110724" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.30" />
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                    <SPLIT distance="75" swimtime="00:01:07.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="327" reactiontime="+88" swimtime="00:02:40.79" resultid="109923" heatid="110766" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.29" />
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="75" swimtime="00:00:57.74" />
                    <SPLIT distance="100" swimtime="00:01:18.40" />
                    <SPLIT distance="125" swimtime="00:01:39.20" />
                    <SPLIT distance="150" swimtime="00:02:00.42" />
                    <SPLIT distance="175" swimtime="00:02:21.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="301" swimtime="00:05:49.80" resultid="109924" heatid="110840" lane="6" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.75" />
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="75" swimtime="00:01:02.20" />
                    <SPLIT distance="100" swimtime="00:01:24.44" />
                    <SPLIT distance="125" swimtime="00:01:46.49" />
                    <SPLIT distance="150" swimtime="00:02:08.81" />
                    <SPLIT distance="175" swimtime="00:02:31.00" />
                    <SPLIT distance="200" swimtime="00:02:53.47" />
                    <SPLIT distance="225" swimtime="00:03:15.91" />
                    <SPLIT distance="250" swimtime="00:03:38.30" />
                    <SPLIT distance="275" swimtime="00:04:00.65" />
                    <SPLIT distance="300" swimtime="00:04:22.77" />
                    <SPLIT distance="325" swimtime="00:04:45.05" />
                    <SPLIT distance="350" swimtime="00:05:07.24" />
                    <SPLIT distance="375" swimtime="00:05:29.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-24" firstname="Przemysław" gender="M" lastname="Bielski" nation="POL" athleteid="109880">
              <RESULTS>
                <RESULT eventid="98798" points="315" reactiontime="+95" swimtime="00:00:29.75" resultid="109881" heatid="110603" lane="1" entrytime="00:00:30.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" status="DNS" swimtime="00:00:00.00" resultid="109882" heatid="110642" lane="8" entrytime="00:23:00.00" />
                <RESULT eventid="106277" points="320" reactiontime="+96" swimtime="00:01:05.70" resultid="109883" heatid="110683" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.38" />
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="75" swimtime="00:00:48.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="109884" heatid="110760" lane="8" entrytime="00:01:25.00" />
                <RESULT eventid="99218" points="269" reactiontime="+86" swimtime="00:02:33.86" resultid="109885" heatid="110773" lane="2" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.26" />
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="75" swimtime="00:00:52.05" />
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="125" swimtime="00:01:30.45" />
                    <SPLIT distance="150" swimtime="00:01:50.84" />
                    <SPLIT distance="175" swimtime="00:02:12.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="109886" heatid="110847" lane="2" entrytime="00:05:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-26" firstname="Joanna" gender="F" lastname="Drzewicka" nation="POL" athleteid="109836">
              <RESULTS>
                <RESULT eventid="98777" points="240" swimtime="00:00:37.38" resultid="109837" heatid="110585" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="243" reactiontime="+83" swimtime="00:00:41.09" resultid="109838" heatid="110645" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="224" reactiontime="+88" swimtime="00:01:30.55" resultid="109839" heatid="110752" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.80" />
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="75" swimtime="00:01:07.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="206" reactiontime="+84" swimtime="00:03:21.81" resultid="109840" heatid="110806" lane="0">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.11" />
                    <SPLIT distance="50" swimtime="00:00:46.98" />
                    <SPLIT distance="75" swimtime="00:01:11.65" />
                    <SPLIT distance="100" swimtime="00:01:38.03" />
                    <SPLIT distance="125" swimtime="00:02:59.50" />
                    <SPLIT distance="150" swimtime="00:02:33.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-26" firstname="Grzegorz" gender="M" lastname="Kalinowski" nation="POL" athleteid="109972">
              <RESULTS>
                <RESULT eventid="98798" points="311" reactiontime="+98" swimtime="00:00:29.88" resultid="109973" heatid="110602" lane="0" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="317" reactiontime="+87" swimtime="00:01:05.90" resultid="109974" heatid="110682" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.66" />
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="75" swimtime="00:00:47.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="222" reactiontime="+99" swimtime="00:01:20.72" resultid="109975" heatid="110759" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.57" />
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="75" swimtime="00:01:00.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-02-09" firstname="Aleksandra" gender="F" lastname="Milewska" nation="POL" athleteid="109893">
              <RESULTS>
                <RESULT eventid="98863" points="333" reactiontime="+90" swimtime="00:11:30.99" resultid="109894" heatid="110633" lane="2" entrytime="00:11:22.22">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.67" />
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="75" swimtime="00:00:57.06" />
                    <SPLIT distance="100" swimtime="00:01:17.36" />
                    <SPLIT distance="125" swimtime="00:01:37.93" />
                    <SPLIT distance="150" swimtime="00:01:58.76" />
                    <SPLIT distance="175" swimtime="00:02:19.93" />
                    <SPLIT distance="200" swimtime="00:02:40.92" />
                    <SPLIT distance="225" swimtime="00:03:02.77" />
                    <SPLIT distance="250" swimtime="00:03:24.28" />
                    <SPLIT distance="275" swimtime="00:03:46.15" />
                    <SPLIT distance="300" swimtime="00:04:07.57" />
                    <SPLIT distance="325" swimtime="00:04:29.14" />
                    <SPLIT distance="350" swimtime="00:04:50.76" />
                    <SPLIT distance="375" swimtime="00:05:12.72" />
                    <SPLIT distance="400" swimtime="00:05:34.97" />
                    <SPLIT distance="425" swimtime="00:05:57.09" />
                    <SPLIT distance="450" swimtime="00:06:19.14" />
                    <SPLIT distance="475" swimtime="00:06:41.35" />
                    <SPLIT distance="500" swimtime="00:07:03.31" />
                    <SPLIT distance="525" swimtime="00:07:25.21" />
                    <SPLIT distance="550" swimtime="00:07:48.06" />
                    <SPLIT distance="575" swimtime="00:08:10.55" />
                    <SPLIT distance="600" swimtime="00:08:32.99" />
                    <SPLIT distance="625" swimtime="00:08:56.08" />
                    <SPLIT distance="650" swimtime="00:09:18.61" />
                    <SPLIT distance="675" swimtime="00:09:41.83" />
                    <SPLIT distance="700" swimtime="00:10:04.43" />
                    <SPLIT distance="725" swimtime="00:10:26.59" />
                    <SPLIT distance="750" swimtime="00:10:48.65" />
                    <SPLIT distance="775" swimtime="00:11:10.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="294" swimtime="00:03:22.34" resultid="109895" heatid="110661" lane="0">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.11" />
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                    <SPLIT distance="75" swimtime="00:01:10.77" />
                    <SPLIT distance="100" swimtime="00:01:36.65" />
                    <SPLIT distance="125" swimtime="00:02:02.56" />
                    <SPLIT distance="150" swimtime="00:02:29.19" />
                    <SPLIT distance="175" swimtime="00:02:55.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="365" reactiontime="+84" swimtime="00:01:19.27" resultid="109896" heatid="110694" lane="3" entrytime="00:01:18.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.84" />
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                    <SPLIT distance="75" swimtime="00:01:00.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="371" reactiontime="+73" swimtime="00:00:33.92" resultid="109897" heatid="110739" lane="3" entrytime="00:00:33.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" status="DNS" swimtime="00:00:00.00" resultid="109898" heatid="110787" lane="1" entrytime="00:06:24.20" />
                <RESULT eventid="99344" points="332" swimtime="00:01:18.82" resultid="109899" heatid="110796" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.19" />
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="75" swimtime="00:00:56.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Zdzisław" gender="M" lastname="Choroszewski" nation="POL" athleteid="109994">
              <RESULTS>
                <RESULT eventid="98798" points="83" swimtime="00:00:46.33" resultid="109995" heatid="110596" lane="9" entrytime="00:00:46.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="73" swimtime="00:33:42.02" resultid="109996" heatid="110643" lane="9" entrytime="00:33:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.36" />
                    <SPLIT distance="50" swimtime="00:00:57.57" />
                    <SPLIT distance="75" swimtime="00:01:29.18" />
                    <SPLIT distance="100" swimtime="00:02:03.49" />
                    <SPLIT distance="125" swimtime="00:02:37.13" />
                    <SPLIT distance="150" swimtime="00:03:09.96" />
                    <SPLIT distance="175" swimtime="00:03:44.67" />
                    <SPLIT distance="200" swimtime="00:04:18.40" />
                    <SPLIT distance="225" swimtime="00:04:53.32" />
                    <SPLIT distance="250" swimtime="00:05:27.11" />
                    <SPLIT distance="275" swimtime="00:06:02.20" />
                    <SPLIT distance="300" swimtime="00:06:36.00" />
                    <SPLIT distance="325" swimtime="00:07:11.54" />
                    <SPLIT distance="350" swimtime="00:07:45.86" />
                    <SPLIT distance="375" swimtime="00:08:22.31" />
                    <SPLIT distance="400" swimtime="00:08:56.24" />
                    <SPLIT distance="425" swimtime="00:09:29.59" />
                    <SPLIT distance="450" swimtime="00:10:04.93" />
                    <SPLIT distance="475" swimtime="00:10:40.20" />
                    <SPLIT distance="500" swimtime="00:11:14.01" />
                    <SPLIT distance="525" swimtime="00:11:49.48" />
                    <SPLIT distance="550" swimtime="00:12:22.48" />
                    <SPLIT distance="575" swimtime="00:12:57.25" />
                    <SPLIT distance="600" swimtime="00:13:31.44" />
                    <SPLIT distance="625" swimtime="00:14:05.83" />
                    <SPLIT distance="650" swimtime="00:14:38.55" />
                    <SPLIT distance="675" swimtime="00:15:13.36" />
                    <SPLIT distance="700" swimtime="00:15:46.75" />
                    <SPLIT distance="725" swimtime="00:16:21.63" />
                    <SPLIT distance="750" swimtime="00:16:55.83" />
                    <SPLIT distance="775" swimtime="00:17:31.32" />
                    <SPLIT distance="800" swimtime="00:18:04.15" />
                    <SPLIT distance="825" swimtime="00:18:38.54" />
                    <SPLIT distance="850" swimtime="00:19:12.85" />
                    <SPLIT distance="875" swimtime="00:19:47.41" />
                    <SPLIT distance="900" swimtime="00:20:20.97" />
                    <SPLIT distance="925" swimtime="00:20:55.87" />
                    <SPLIT distance="950" swimtime="00:21:28.77" />
                    <SPLIT distance="975" swimtime="00:22:03.31" />
                    <SPLIT distance="1000" swimtime="00:22:36.82" />
                    <SPLIT distance="1025" swimtime="00:23:11.35" />
                    <SPLIT distance="1050" swimtime="00:23:44.77" />
                    <SPLIT distance="1075" swimtime="00:24:18.68" />
                    <SPLIT distance="1100" swimtime="00:24:51.17" />
                    <SPLIT distance="1125" swimtime="00:25:24.34" />
                    <SPLIT distance="1150" swimtime="00:25:58.31" />
                    <SPLIT distance="1175" swimtime="00:26:32.00" />
                    <SPLIT distance="1200" swimtime="00:27:05.47" />
                    <SPLIT distance="1225" swimtime="00:27:40.21" />
                    <SPLIT distance="1250" swimtime="00:28:12.59" />
                    <SPLIT distance="1275" swimtime="00:28:47.06" />
                    <SPLIT distance="1300" swimtime="00:29:19.74" />
                    <SPLIT distance="1325" swimtime="00:29:53.69" />
                    <SPLIT distance="1350" swimtime="00:30:25.68" />
                    <SPLIT distance="1375" swimtime="00:30:58.97" />
                    <SPLIT distance="1400" swimtime="00:31:31.75" />
                    <SPLIT distance="1425" swimtime="00:32:05.08" />
                    <SPLIT distance="1450" swimtime="00:32:38.39" />
                    <SPLIT distance="1475" swimtime="00:33:12.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="70" reactiontime="+100" swimtime="00:08:32.73" resultid="109997" heatid="110852" lane="4" entrytime="00:08:49.79">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.35" />
                    <SPLIT distance="50" swimtime="00:00:53.77" />
                    <SPLIT distance="75" swimtime="00:01:24.58" />
                    <SPLIT distance="100" swimtime="00:01:56.72" />
                    <SPLIT distance="125" swimtime="00:02:30.13" />
                    <SPLIT distance="150" swimtime="00:03:03.19" />
                    <SPLIT distance="175" swimtime="00:03:37.45" />
                    <SPLIT distance="200" swimtime="00:04:10.97" />
                    <SPLIT distance="225" swimtime="00:04:44.83" />
                    <SPLIT distance="250" swimtime="00:05:18.44" />
                    <SPLIT distance="275" swimtime="00:05:51.82" />
                    <SPLIT distance="300" swimtime="00:06:25.92" />
                    <SPLIT distance="325" swimtime="00:06:59.34" />
                    <SPLIT distance="350" swimtime="00:07:32.03" />
                    <SPLIT distance="375" swimtime="00:08:04.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-26" firstname="Aleksandra" gender="F" lastname="Przybysz" nation="POL" athleteid="109871">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="109872" heatid="110589" lane="5" entrytime="00:00:34.76" />
                <RESULT eventid="106254" points="280" reactiontime="+94" swimtime="00:23:25.40" resultid="109873" heatid="110640" lane="6" entrytime="00:23:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.11" />
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="75" swimtime="00:01:03.06" />
                    <SPLIT distance="100" swimtime="00:01:25.21" />
                    <SPLIT distance="125" swimtime="00:01:47.55" />
                    <SPLIT distance="150" swimtime="00:02:10.56" />
                    <SPLIT distance="175" swimtime="00:02:33.42" />
                    <SPLIT distance="200" swimtime="00:02:56.74" />
                    <SPLIT distance="225" swimtime="00:03:19.83" />
                    <SPLIT distance="250" swimtime="00:03:43.09" />
                    <SPLIT distance="275" swimtime="00:04:06.26" />
                    <SPLIT distance="300" swimtime="00:04:29.62" />
                    <SPLIT distance="325" swimtime="00:04:52.78" />
                    <SPLIT distance="350" swimtime="00:05:16.08" />
                    <SPLIT distance="375" swimtime="00:05:39.24" />
                    <SPLIT distance="400" swimtime="00:06:02.79" />
                    <SPLIT distance="425" swimtime="00:06:25.95" />
                    <SPLIT distance="450" swimtime="00:06:49.34" />
                    <SPLIT distance="475" swimtime="00:07:12.41" />
                    <SPLIT distance="500" swimtime="00:07:36.28" />
                    <SPLIT distance="525" swimtime="00:07:59.36" />
                    <SPLIT distance="550" swimtime="00:08:23.02" />
                    <SPLIT distance="575" swimtime="00:08:46.35" />
                    <SPLIT distance="600" swimtime="00:09:09.71" />
                    <SPLIT distance="625" swimtime="00:09:33.51" />
                    <SPLIT distance="650" swimtime="00:09:57.83" />
                    <SPLIT distance="675" swimtime="00:10:20.78" />
                    <SPLIT distance="700" swimtime="00:10:44.79" />
                    <SPLIT distance="725" swimtime="00:11:08.52" />
                    <SPLIT distance="750" swimtime="00:11:32.20" />
                    <SPLIT distance="775" swimtime="00:11:55.64" />
                    <SPLIT distance="800" swimtime="00:12:19.48" />
                    <SPLIT distance="825" swimtime="00:12:43.12" />
                    <SPLIT distance="850" swimtime="00:13:07.38" />
                    <SPLIT distance="875" swimtime="00:13:31.33" />
                    <SPLIT distance="900" swimtime="00:13:55.30" />
                    <SPLIT distance="925" swimtime="00:14:18.60" />
                    <SPLIT distance="950" swimtime="00:14:42.71" />
                    <SPLIT distance="975" swimtime="00:15:06.16" />
                    <SPLIT distance="1000" swimtime="00:15:30.47" />
                    <SPLIT distance="1025" swimtime="00:15:54.95" />
                    <SPLIT distance="1050" swimtime="00:16:19.11" />
                    <SPLIT distance="1075" swimtime="00:16:42.69" />
                    <SPLIT distance="1100" swimtime="00:17:06.98" />
                    <SPLIT distance="1125" swimtime="00:17:30.50" />
                    <SPLIT distance="1150" swimtime="00:17:54.30" />
                    <SPLIT distance="1175" swimtime="00:18:18.02" />
                    <SPLIT distance="1200" swimtime="00:18:42.26" />
                    <SPLIT distance="1225" swimtime="00:19:06.41" />
                    <SPLIT distance="1250" swimtime="00:19:30.12" />
                    <SPLIT distance="1275" swimtime="00:19:54.34" />
                    <SPLIT distance="1300" swimtime="00:20:18.43" />
                    <SPLIT distance="1325" swimtime="00:20:41.82" />
                    <SPLIT distance="1350" swimtime="00:21:06.00" />
                    <SPLIT distance="1375" swimtime="00:21:29.47" />
                    <SPLIT distance="1400" swimtime="00:21:53.62" />
                    <SPLIT distance="1425" swimtime="00:22:17.16" />
                    <SPLIT distance="1450" swimtime="00:22:41.17" />
                    <SPLIT distance="1475" swimtime="00:23:03.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="109874" heatid="110674" lane="3" entrytime="00:01:14.38" />
                <RESULT eventid="99004" points="236" reactiontime="+91" swimtime="00:03:13.38" resultid="109875" heatid="110708" lane="3" entrytime="00:03:09.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.68" />
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="75" swimtime="00:01:07.25" />
                    <SPLIT distance="100" swimtime="00:01:32.13" />
                    <SPLIT distance="125" swimtime="00:01:57.38" />
                    <SPLIT distance="150" swimtime="00:02:22.82" />
                    <SPLIT distance="175" swimtime="00:02:47.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="251" reactiontime="+84" swimtime="00:01:27.14" resultid="109876" heatid="110754" lane="7" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.04" />
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="75" swimtime="00:01:05.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="307" reactiontime="+85" swimtime="00:02:44.06" resultid="109877" heatid="110767" lane="7" entrytime="00:02:41.43">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.49" />
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="75" swimtime="00:00:58.64" />
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                    <SPLIT distance="125" swimtime="00:01:40.87" />
                    <SPLIT distance="150" swimtime="00:02:02.46" />
                    <SPLIT distance="175" swimtime="00:02:23.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="254" swimtime="00:01:26.21" resultid="109878" heatid="110795" lane="2" entrytime="00:01:25.05">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.02" />
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                    <SPLIT distance="75" swimtime="00:01:03.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="303" reactiontime="+91" swimtime="00:05:49.01" resultid="109879" heatid="110840" lane="5" entrytime="00:05:43.83">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.16" />
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="75" swimtime="00:01:02.02" />
                    <SPLIT distance="100" swimtime="00:01:23.70" />
                    <SPLIT distance="125" swimtime="00:01:45.47" />
                    <SPLIT distance="150" swimtime="00:02:07.32" />
                    <SPLIT distance="175" swimtime="00:02:29.64" />
                    <SPLIT distance="200" swimtime="00:02:51.59" />
                    <SPLIT distance="225" swimtime="00:03:14.10" />
                    <SPLIT distance="250" swimtime="00:03:36.76" />
                    <SPLIT distance="275" swimtime="00:03:59.15" />
                    <SPLIT distance="300" swimtime="00:04:21.33" />
                    <SPLIT distance="325" swimtime="00:04:43.81" />
                    <SPLIT distance="350" swimtime="00:05:06.29" />
                    <SPLIT distance="375" swimtime="00:05:28.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="109821">
              <RESULTS>
                <RESULT eventid="98814" points="229" reactiontime="+91" swimtime="00:03:18.99" resultid="109822" heatid="110615" lane="5" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.33" />
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                    <SPLIT distance="75" swimtime="00:01:11.43" />
                    <SPLIT distance="100" swimtime="00:01:36.65" />
                    <SPLIT distance="125" swimtime="00:02:04.82" />
                    <SPLIT distance="150" swimtime="00:02:32.33" />
                    <SPLIT distance="175" swimtime="00:02:56.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="295" reactiontime="+85" swimtime="00:11:59.55" resultid="109823" heatid="110633" lane="8" entrytime="00:11:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.87" />
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="75" swimtime="00:01:00.76" />
                    <SPLIT distance="100" swimtime="00:01:22.66" />
                    <SPLIT distance="125" swimtime="00:01:44.47" />
                    <SPLIT distance="150" swimtime="00:02:06.66" />
                    <SPLIT distance="175" swimtime="00:02:29.07" />
                    <SPLIT distance="200" swimtime="00:02:51.81" />
                    <SPLIT distance="225" swimtime="00:03:14.53" />
                    <SPLIT distance="250" swimtime="00:03:37.32" />
                    <SPLIT distance="275" swimtime="00:04:00.12" />
                    <SPLIT distance="300" swimtime="00:04:23.13" />
                    <SPLIT distance="325" swimtime="00:04:45.85" />
                    <SPLIT distance="350" swimtime="00:05:08.68" />
                    <SPLIT distance="375" swimtime="00:05:31.48" />
                    <SPLIT distance="400" swimtime="00:05:54.40" />
                    <SPLIT distance="425" swimtime="00:06:17.12" />
                    <SPLIT distance="450" swimtime="00:06:40.03" />
                    <SPLIT distance="475" swimtime="00:07:02.82" />
                    <SPLIT distance="500" swimtime="00:07:25.73" />
                    <SPLIT distance="525" swimtime="00:07:48.36" />
                    <SPLIT distance="550" swimtime="00:08:11.27" />
                    <SPLIT distance="575" swimtime="00:08:34.54" />
                    <SPLIT distance="600" swimtime="00:08:57.26" />
                    <SPLIT distance="625" swimtime="00:09:20.08" />
                    <SPLIT distance="650" swimtime="00:09:43.40" />
                    <SPLIT distance="675" swimtime="00:10:06.47" />
                    <SPLIT distance="700" swimtime="00:10:28.86" />
                    <SPLIT distance="725" swimtime="00:10:51.65" />
                    <SPLIT distance="750" swimtime="00:11:14.46" />
                    <SPLIT distance="775" swimtime="00:11:36.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="250" reactiontime="+87" swimtime="00:03:33.59" resultid="109824" heatid="110662" lane="5" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.78" />
                    <SPLIT distance="50" swimtime="00:00:49.02" />
                    <SPLIT distance="75" swimtime="00:01:16.06" />
                    <SPLIT distance="100" swimtime="00:01:43.36" />
                    <SPLIT distance="125" swimtime="00:02:10.90" />
                    <SPLIT distance="150" swimtime="00:02:38.22" />
                    <SPLIT distance="175" swimtime="00:03:05.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="313" reactiontime="+85" swimtime="00:01:14.93" resultid="109825" heatid="110674" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.12" />
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="75" swimtime="00:00:55.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="314" reactiontime="+85" swimtime="00:02:42.89" resultid="109826" heatid="110764" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.20" />
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="75" swimtime="00:00:58.69" />
                    <SPLIT distance="100" swimtime="00:01:19.63" />
                    <SPLIT distance="125" swimtime="00:01:40.98" />
                    <SPLIT distance="150" swimtime="00:02:02.06" />
                    <SPLIT distance="175" swimtime="00:02:22.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="251" reactiontime="+97" swimtime="00:06:51.30" resultid="109827" heatid="110786" lane="2" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.26" />
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                    <SPLIT distance="75" swimtime="00:01:14.57" />
                    <SPLIT distance="100" swimtime="00:01:42.34" />
                    <SPLIT distance="125" swimtime="00:02:09.38" />
                    <SPLIT distance="150" swimtime="00:02:35.07" />
                    <SPLIT distance="175" swimtime="00:03:00.73" />
                    <SPLIT distance="200" swimtime="00:03:27.32" />
                    <SPLIT distance="225" swimtime="00:03:55.40" />
                    <SPLIT distance="250" swimtime="00:04:23.76" />
                    <SPLIT distance="275" swimtime="00:04:52.10" />
                    <SPLIT distance="300" swimtime="00:05:20.88" />
                    <SPLIT distance="325" swimtime="00:05:44.63" />
                    <SPLIT distance="350" swimtime="00:06:07.27" />
                    <SPLIT distance="375" swimtime="00:06:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="201" reactiontime="+89" swimtime="00:03:23.39" resultid="109828" heatid="110807" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.12" />
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                    <SPLIT distance="75" swimtime="00:01:12.45" />
                    <SPLIT distance="100" swimtime="00:01:38.34" />
                    <SPLIT distance="125" swimtime="00:02:04.15" />
                    <SPLIT distance="150" swimtime="00:02:31.06" />
                    <SPLIT distance="175" swimtime="00:02:58.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="306" reactiontime="+93" swimtime="00:05:47.72" resultid="109829" heatid="110840" lane="3" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.75" />
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                    <SPLIT distance="75" swimtime="00:01:01.36" />
                    <SPLIT distance="100" swimtime="00:01:23.00" />
                    <SPLIT distance="125" swimtime="00:01:45.29" />
                    <SPLIT distance="150" swimtime="00:02:07.61" />
                    <SPLIT distance="175" swimtime="00:02:30.10" />
                    <SPLIT distance="200" swimtime="00:02:52.63" />
                    <SPLIT distance="225" swimtime="00:03:15.10" />
                    <SPLIT distance="250" swimtime="00:03:37.38" />
                    <SPLIT distance="275" swimtime="00:03:59.59" />
                    <SPLIT distance="300" swimtime="00:04:21.50" />
                    <SPLIT distance="325" swimtime="00:04:43.45" />
                    <SPLIT distance="350" swimtime="00:05:05.15" />
                    <SPLIT distance="375" swimtime="00:05:26.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-03-18" firstname="Danuta" gender="F" lastname="Wegen" nation="POL" athleteid="109911">
              <RESULTS>
                <RESULT eventid="98777" points="127" swimtime="00:00:46.13" resultid="109912" heatid="110587" lane="9" entrytime="00:00:47.22">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="96" swimtime="00:17:23.75" resultid="109913" heatid="110634" lane="6" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.76" />
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                    <SPLIT distance="75" swimtime="00:01:20.35" />
                    <SPLIT distance="100" swimtime="00:01:53.07" />
                    <SPLIT distance="125" swimtime="00:02:23.97" />
                    <SPLIT distance="150" swimtime="00:02:57.94" />
                    <SPLIT distance="175" swimtime="00:03:30.85" />
                    <SPLIT distance="200" swimtime="00:04:05.11" />
                    <SPLIT distance="225" swimtime="00:04:36.24" />
                    <SPLIT distance="250" swimtime="00:05:10.47" />
                    <SPLIT distance="275" swimtime="00:05:43.68" />
                    <SPLIT distance="300" swimtime="00:06:16.70" />
                    <SPLIT distance="325" swimtime="00:06:49.39" />
                    <SPLIT distance="350" swimtime="00:07:23.62" />
                    <SPLIT distance="375" swimtime="00:07:57.49" />
                    <SPLIT distance="400" swimtime="00:08:31.30" />
                    <SPLIT distance="425" swimtime="00:09:05.06" />
                    <SPLIT distance="450" swimtime="00:09:39.51" />
                    <SPLIT distance="475" swimtime="00:10:11.48" />
                    <SPLIT distance="500" swimtime="00:10:45.11" />
                    <SPLIT distance="525" swimtime="00:11:18.14" />
                    <SPLIT distance="550" swimtime="00:11:51.84" />
                    <SPLIT distance="575" swimtime="00:12:25.17" />
                    <SPLIT distance="600" swimtime="00:12:58.90" />
                    <SPLIT distance="625" swimtime="00:13:31.05" />
                    <SPLIT distance="650" swimtime="00:14:05.93" />
                    <SPLIT distance="675" swimtime="00:14:38.25" />
                    <SPLIT distance="700" swimtime="00:15:13.06" />
                    <SPLIT distance="725" swimtime="00:15:44.94" />
                    <SPLIT distance="750" swimtime="00:16:18.23" />
                    <SPLIT distance="775" swimtime="00:16:51.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="118" reactiontime="+74" swimtime="00:00:52.19" resultid="109914" heatid="110646" lane="5" entrytime="00:00:55.14">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="107" swimtime="00:01:46.98" resultid="109915" heatid="110672" lane="9" entrytime="00:02:14.06">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.21" />
                    <SPLIT distance="50" swimtime="00:00:50.20" />
                    <SPLIT distance="75" swimtime="00:01:18.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="101" reactiontime="+84" swimtime="00:01:58.13" resultid="109916" heatid="110754" lane="9" entrytime="00:01:59.49">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.62" />
                    <SPLIT distance="50" swimtime="00:00:55.49" />
                    <SPLIT distance="75" swimtime="00:01:26.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="95" reactiontime="+94" swimtime="00:04:02.59" resultid="109917" heatid="110764" lane="5" entrytime="00:03:34.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.49" />
                    <SPLIT distance="50" swimtime="00:00:51.57" />
                    <SPLIT distance="75" swimtime="00:01:22.25" />
                    <SPLIT distance="100" swimtime="00:01:54.55" />
                    <SPLIT distance="125" swimtime="00:02:26.79" />
                    <SPLIT distance="150" swimtime="00:02:59.62" />
                    <SPLIT distance="175" swimtime="00:03:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="111" reactiontime="+90" swimtime="00:04:07.49" resultid="109918" heatid="110806" lane="5" entrytime="00:04:27.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.54" />
                    <SPLIT distance="50" swimtime="00:00:58.39" />
                    <SPLIT distance="75" swimtime="00:01:30.12" />
                    <SPLIT distance="100" swimtime="00:02:01.47" />
                    <SPLIT distance="125" swimtime="00:02:35.32" />
                    <SPLIT distance="150" swimtime="00:03:07.24" />
                    <SPLIT distance="175" swimtime="00:03:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="104" reactiontime="+85" swimtime="00:08:17.33" resultid="109919" heatid="110842" lane="7" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.97" />
                    <SPLIT distance="50" swimtime="00:00:52.66" />
                    <SPLIT distance="75" swimtime="00:01:23.00" />
                    <SPLIT distance="100" swimtime="00:01:55.22" />
                    <SPLIT distance="125" swimtime="00:02:28.35" />
                    <SPLIT distance="150" swimtime="00:03:00.37" />
                    <SPLIT distance="175" swimtime="00:03:32.80" />
                    <SPLIT distance="200" swimtime="00:04:04.40" />
                    <SPLIT distance="225" swimtime="00:04:36.65" />
                    <SPLIT distance="250" swimtime="00:05:09.56" />
                    <SPLIT distance="275" swimtime="00:05:42.08" />
                    <SPLIT distance="300" swimtime="00:06:13.45" />
                    <SPLIT distance="325" swimtime="00:06:44.98" />
                    <SPLIT distance="350" swimtime="00:07:17.24" />
                    <SPLIT distance="375" swimtime="00:07:48.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Piotr" gender="M" lastname="Konopacki" nation="POL" athleteid="109932">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="109933" heatid="110599" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="98924" points="278" reactiontime="+70" swimtime="00:00:34.04" resultid="109934" heatid="110658" lane="8" entrytime="00:00:32.94">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="389" reactiontime="+86" swimtime="00:01:01.52" resultid="109935" heatid="110685" lane="1" entrytime="00:01:02.94">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.83" />
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="75" swimtime="00:00:45.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="109936" heatid="110761" lane="6" entrytime="00:01:14.68" />
                <RESULT eventid="99218" points="366" reactiontime="+77" swimtime="00:02:18.88" resultid="109937" heatid="110773" lane="3" entrytime="00:02:30.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.52" />
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="75" swimtime="00:00:48.87" />
                    <SPLIT distance="100" swimtime="00:01:07.01" />
                    <SPLIT distance="125" swimtime="00:01:24.55" />
                    <SPLIT distance="150" swimtime="00:01:42.55" />
                    <SPLIT distance="175" swimtime="00:02:01.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="344" swimtime="00:05:02.79" resultid="109938" heatid="110852" lane="6">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.03" />
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="75" swimtime="00:00:51.36" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="125" swimtime="00:01:29.31" />
                    <SPLIT distance="150" swimtime="00:01:48.39" />
                    <SPLIT distance="175" swimtime="00:02:07.25" />
                    <SPLIT distance="200" swimtime="00:02:26.78" />
                    <SPLIT distance="225" swimtime="00:02:46.32" />
                    <SPLIT distance="250" swimtime="00:03:06.16" />
                    <SPLIT distance="275" swimtime="00:03:26.22" />
                    <SPLIT distance="300" swimtime="00:03:46.26" />
                    <SPLIT distance="325" swimtime="00:04:06.23" />
                    <SPLIT distance="350" swimtime="00:04:26.15" />
                    <SPLIT distance="375" swimtime="00:04:45.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="335" reactiontime="+73" swimtime="00:10:38.19" resultid="110020" heatid="110635" lane="8" entrytime="00:10:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.67" />
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="75" swimtime="00:00:53.72" />
                    <SPLIT distance="100" swimtime="00:01:13.61" />
                    <SPLIT distance="125" swimtime="00:01:33.47" />
                    <SPLIT distance="150" swimtime="00:01:53.85" />
                    <SPLIT distance="175" swimtime="00:02:14.08" />
                    <SPLIT distance="200" swimtime="00:02:34.19" />
                    <SPLIT distance="225" swimtime="00:02:54.56" />
                    <SPLIT distance="250" swimtime="00:03:15.08" />
                    <SPLIT distance="275" swimtime="00:03:35.39" />
                    <SPLIT distance="300" swimtime="00:03:55.62" />
                    <SPLIT distance="325" swimtime="00:04:15.89" />
                    <SPLIT distance="350" swimtime="00:04:36.19" />
                    <SPLIT distance="375" swimtime="00:04:56.41" />
                    <SPLIT distance="400" swimtime="00:05:16.85" />
                    <SPLIT distance="425" swimtime="00:05:37.02" />
                    <SPLIT distance="450" swimtime="00:05:57.39" />
                    <SPLIT distance="475" swimtime="00:06:17.67" />
                    <SPLIT distance="500" swimtime="00:06:38.17" />
                    <SPLIT distance="525" swimtime="00:06:58.56" />
                    <SPLIT distance="550" swimtime="00:07:18.84" />
                    <SPLIT distance="575" swimtime="00:07:39.29" />
                    <SPLIT distance="600" swimtime="00:07:59.55" />
                    <SPLIT distance="625" swimtime="00:08:19.87" />
                    <SPLIT distance="650" swimtime="00:08:40.24" />
                    <SPLIT distance="675" swimtime="00:09:00.49" />
                    <SPLIT distance="700" swimtime="00:09:20.65" />
                    <SPLIT distance="725" swimtime="00:09:40.79" />
                    <SPLIT distance="750" swimtime="00:10:00.79" />
                    <SPLIT distance="775" swimtime="00:10:20.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-12-31" firstname="Marek" gender="M" lastname="Hasso-Agopsowicz" nation="POL" athleteid="109982">
              <RESULTS>
                <RESULT eventid="98891" points="75" reactiontime="+117" swimtime="00:17:30.99" resultid="109983" heatid="110637" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.82" />
                    <SPLIT distance="50" swimtime="00:00:53.73" />
                    <SPLIT distance="75" swimtime="00:01:24.80" />
                    <SPLIT distance="100" swimtime="00:01:56.34" />
                    <SPLIT distance="125" swimtime="00:02:29.46" />
                    <SPLIT distance="150" swimtime="00:03:01.68" />
                    <SPLIT distance="175" swimtime="00:03:34.18" />
                    <SPLIT distance="200" swimtime="00:04:06.34" />
                    <SPLIT distance="225" swimtime="00:04:38.89" />
                    <SPLIT distance="250" swimtime="00:05:12.37" />
                    <SPLIT distance="275" swimtime="00:05:46.76" />
                    <SPLIT distance="300" swimtime="00:06:20.85" />
                    <SPLIT distance="325" swimtime="00:06:54.34" />
                    <SPLIT distance="350" swimtime="00:07:28.52" />
                    <SPLIT distance="375" swimtime="00:08:00.97" />
                    <SPLIT distance="400" swimtime="00:08:34.39" />
                    <SPLIT distance="425" swimtime="00:09:08.34" />
                    <SPLIT distance="450" swimtime="00:09:42.33" />
                    <SPLIT distance="475" swimtime="00:10:16.30" />
                    <SPLIT distance="500" swimtime="00:10:50.27" />
                    <SPLIT distance="525" swimtime="00:11:23.82" />
                    <SPLIT distance="550" swimtime="00:11:57.22" />
                    <SPLIT distance="575" swimtime="00:12:29.67" />
                    <SPLIT distance="600" swimtime="00:12:28.77" />
                    <SPLIT distance="625" swimtime="00:13:36.64" />
                    <SPLIT distance="650" swimtime="00:13:03.77" />
                    <SPLIT distance="675" swimtime="00:14:44.38" />
                    <SPLIT distance="700" swimtime="00:14:10.65" />
                    <SPLIT distance="725" swimtime="00:15:52.12" />
                    <SPLIT distance="750" swimtime="00:15:17.82" />
                    <SPLIT distance="775" swimtime="00:16:59.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="86" reactiontime="+108" swimtime="00:00:57.14" resultid="109984" heatid="110824" lane="2">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="109862">
              <RESULTS>
                <RESULT eventid="98798" points="499" reactiontime="+66" swimtime="00:00:25.53" resultid="109863" heatid="110608" lane="6" entrytime="00:00:27.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="450" reactiontime="+62" swimtime="00:02:22.97" resultid="109864" heatid="110627" lane="5" entrytime="00:02:26.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="75" swimtime="00:00:50.15" />
                    <SPLIT distance="100" swimtime="00:01:09.01" />
                    <SPLIT distance="125" swimtime="00:01:29.21" />
                    <SPLIT distance="150" swimtime="00:01:49.94" />
                    <SPLIT distance="175" swimtime="00:02:07.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="537" swimtime="00:00:55.26" resultid="109865" heatid="110681" lane="9" entrytime="00:01:16.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.79" />
                    <SPLIT distance="50" swimtime="00:00:26.63" />
                    <SPLIT distance="75" swimtime="00:00:40.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="476" reactiontime="+79" swimtime="00:01:04.88" resultid="109866" heatid="110705" lane="1" entrytime="00:01:05.95">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.37" />
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="75" swimtime="00:00:49.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="464" reactiontime="+83" swimtime="00:00:28.15" resultid="109867" heatid="110749" lane="2" entrytime="00:00:28.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="422" reactiontime="+72" swimtime="00:05:13.78" resultid="109868" heatid="110792" lane="8" entrytime="00:05:23.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.33" />
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="75" swimtime="00:00:50.06" />
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                    <SPLIT distance="125" swimtime="00:01:30.94" />
                    <SPLIT distance="150" swimtime="00:01:52.23" />
                    <SPLIT distance="175" swimtime="00:02:13.10" />
                    <SPLIT distance="200" swimtime="00:02:34.01" />
                    <SPLIT distance="225" swimtime="00:02:56.49" />
                    <SPLIT distance="250" swimtime="00:03:18.83" />
                    <SPLIT distance="275" swimtime="00:03:41.13" />
                    <SPLIT distance="300" swimtime="00:04:03.63" />
                    <SPLIT distance="325" swimtime="00:04:22.19" />
                    <SPLIT distance="350" swimtime="00:04:39.47" />
                    <SPLIT distance="375" swimtime="00:04:56.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="473" reactiontime="+62" swimtime="00:01:02.15" resultid="109869" heatid="110804" lane="5" entrytime="00:01:03.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="75" swimtime="00:00:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="486" reactiontime="+84" swimtime="00:04:29.81" resultid="109870" heatid="110843" lane="2" entrytime="00:04:29.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.81" />
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="75" swimtime="00:00:48.26" />
                    <SPLIT distance="100" swimtime="00:01:05.16" />
                    <SPLIT distance="125" swimtime="00:01:22.09" />
                    <SPLIT distance="150" swimtime="00:01:39.32" />
                    <SPLIT distance="175" swimtime="00:01:56.52" />
                    <SPLIT distance="200" swimtime="00:02:13.97" />
                    <SPLIT distance="225" swimtime="00:02:30.71" />
                    <SPLIT distance="250" swimtime="00:02:47.74" />
                    <SPLIT distance="275" swimtime="00:03:05.01" />
                    <SPLIT distance="300" swimtime="00:03:22.13" />
                    <SPLIT distance="325" swimtime="00:03:39.36" />
                    <SPLIT distance="350" swimtime="00:03:56.76" />
                    <SPLIT distance="375" swimtime="00:04:13.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-29" firstname="Jakub" gender="M" lastname="Stępień" nation="POL" athleteid="109830">
              <RESULTS>
                <RESULT eventid="98798" points="349" reactiontime="+89" swimtime="00:00:28.76" resultid="109831" heatid="110604" lane="1" entrytime="00:00:29.95">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="239" swimtime="00:11:54.14" resultid="109832" heatid="110638" lane="9">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.87" />
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="75" swimtime="00:01:00.24" />
                    <SPLIT distance="100" swimtime="00:01:21.63" />
                    <SPLIT distance="125" swimtime="00:01:43.95" />
                    <SPLIT distance="150" swimtime="00:02:05.73" />
                    <SPLIT distance="175" swimtime="00:02:28.03" />
                    <SPLIT distance="200" swimtime="00:02:50.64" />
                    <SPLIT distance="225" swimtime="00:03:13.01" />
                    <SPLIT distance="250" swimtime="00:03:35.91" />
                    <SPLIT distance="275" swimtime="00:03:58.18" />
                    <SPLIT distance="300" swimtime="00:04:21.06" />
                    <SPLIT distance="325" swimtime="00:04:44.63" />
                    <SPLIT distance="350" swimtime="00:05:07.28" />
                    <SPLIT distance="375" swimtime="00:05:30.79" />
                    <SPLIT distance="400" swimtime="00:05:53.67" />
                    <SPLIT distance="425" swimtime="00:06:16.82" />
                    <SPLIT distance="450" swimtime="00:06:40.42" />
                    <SPLIT distance="475" swimtime="00:07:04.24" />
                    <SPLIT distance="500" swimtime="00:07:27.63" />
                    <SPLIT distance="525" swimtime="00:07:50.46" />
                    <SPLIT distance="550" swimtime="00:08:14.18" />
                    <SPLIT distance="575" swimtime="00:08:37.14" />
                    <SPLIT distance="600" swimtime="00:09:00.04" />
                    <SPLIT distance="625" swimtime="00:09:22.87" />
                    <SPLIT distance="650" swimtime="00:10:30.48" />
                    <SPLIT distance="675" swimtime="00:10:08.15" />
                    <SPLIT distance="700" swimtime="00:11:14.29" />
                    <SPLIT distance="725" swimtime="00:10:52.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="363" swimtime="00:01:02.96" resultid="109833" heatid="110684" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.48" />
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                    <SPLIT distance="75" swimtime="00:00:46.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="257" reactiontime="+91" swimtime="00:00:34.25" resultid="109834" heatid="110744" lane="7" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="323" swimtime="00:02:24.82" resultid="109835" heatid="110774" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.51" />
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="75" swimtime="00:00:49.98" />
                    <SPLIT distance="100" swimtime="00:01:08.73" />
                    <SPLIT distance="125" swimtime="00:01:27.99" />
                    <SPLIT distance="150" swimtime="00:01:47.73" />
                    <SPLIT distance="175" swimtime="00:02:07.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-13" firstname="Michał" gender="M" lastname="Kieres" nation="POL" athleteid="109964">
              <RESULTS>
                <RESULT eventid="98830" points="298" reactiontime="+94" swimtime="00:02:44.03" resultid="109965" heatid="110627" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.89" />
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="125" swimtime="00:01:41.51" />
                    <SPLIT distance="150" swimtime="00:02:04.40" />
                    <SPLIT distance="175" swimtime="00:02:25.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="378" reactiontime="+52" swimtime="00:02:46.56" resultid="109966" heatid="110670" lane="0" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.60" />
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="75" swimtime="00:00:56.94" />
                    <SPLIT distance="100" swimtime="00:01:18.34" />
                    <SPLIT distance="125" swimtime="00:01:39.98" />
                    <SPLIT distance="150" swimtime="00:02:02.43" />
                    <SPLIT distance="175" swimtime="00:02:23.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="329" reactiontime="+90" swimtime="00:01:13.32" resultid="109967" heatid="110703" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.92" />
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="75" swimtime="00:00:55.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="391" swimtime="00:01:16.02" resultid="109968" heatid="110734" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.05" />
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="75" swimtime="00:00:55.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="339" reactiontime="+62" swimtime="00:05:37.57" resultid="109969" heatid="110791" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.58" />
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="75" swimtime="00:00:51.56" />
                    <SPLIT distance="100" swimtime="00:01:11.45" />
                    <SPLIT distance="125" swimtime="00:01:34.93" />
                    <SPLIT distance="150" swimtime="00:01:58.27" />
                    <SPLIT distance="175" swimtime="00:02:21.74" />
                    <SPLIT distance="200" swimtime="00:02:45.77" />
                    <SPLIT distance="225" swimtime="00:03:08.54" />
                    <SPLIT distance="250" swimtime="00:03:31.56" />
                    <SPLIT distance="275" swimtime="00:03:55.09" />
                    <SPLIT distance="300" swimtime="00:04:18.91" />
                    <SPLIT distance="325" swimtime="00:04:39.99" />
                    <SPLIT distance="350" swimtime="00:04:59.76" />
                    <SPLIT distance="375" swimtime="00:05:19.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="334" reactiontime="+82" swimtime="00:01:09.79" resultid="109970" heatid="110803" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.51" />
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="75" swimtime="00:00:50.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="401" reactiontime="+75" swimtime="00:00:34.22" resultid="109971" heatid="110831" lane="5" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-21" firstname="Tomasz" gender="M" lastname="Kozłowski" nation="POL" athleteid="109813">
              <RESULTS>
                <RESULT eventid="98956" points="162" reactiontime="+71" swimtime="00:03:40.91" resultid="109814" heatid="110666" lane="2" entrytime="00:03:53.69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.76" />
                    <SPLIT distance="50" swimtime="00:00:49.28" />
                    <SPLIT distance="75" swimtime="00:01:16.53" />
                    <SPLIT distance="100" swimtime="00:01:45.54" />
                    <SPLIT distance="125" swimtime="00:02:14.92" />
                    <SPLIT distance="150" swimtime="00:02:43.76" />
                    <SPLIT distance="175" swimtime="00:03:12.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="176" reactiontime="+90" swimtime="00:01:39.19" resultid="109815" heatid="110728" lane="1" entrytime="00:01:47.36">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.65" />
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                    <SPLIT distance="75" swimtime="00:01:13.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="109816" heatid="110811" lane="4" entrytime="00:03:43.85" />
                <RESULT eventid="99425" points="177" swimtime="00:00:44.91" resultid="109817" heatid="110826" lane="0" entrytime="00:00:45.71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-07" firstname="Elżbieta" gender="F" lastname="Buczyńska" nation="POL" athleteid="109976">
              <RESULTS>
                <RESULT eventid="98863" points="180" reactiontime="+112" swimtime="00:14:08.66" resultid="109977" heatid="110634" lane="2" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.50" />
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                    <SPLIT distance="75" swimtime="00:01:06.94" />
                    <SPLIT distance="100" swimtime="00:01:31.89" />
                    <SPLIT distance="125" swimtime="00:01:58.30" />
                    <SPLIT distance="150" swimtime="00:02:24.38" />
                    <SPLIT distance="175" swimtime="00:02:51.16" />
                    <SPLIT distance="200" swimtime="00:03:18.20" />
                    <SPLIT distance="225" swimtime="00:03:45.38" />
                    <SPLIT distance="250" swimtime="00:04:12.54" />
                    <SPLIT distance="275" swimtime="00:04:39.53" />
                    <SPLIT distance="300" swimtime="00:05:07.02" />
                    <SPLIT distance="325" swimtime="00:05:34.03" />
                    <SPLIT distance="350" swimtime="00:06:01.71" />
                    <SPLIT distance="375" swimtime="00:06:29.01" />
                    <SPLIT distance="400" swimtime="00:06:56.46" />
                    <SPLIT distance="425" swimtime="00:07:23.47" />
                    <SPLIT distance="450" swimtime="00:07:50.88" />
                    <SPLIT distance="475" swimtime="00:08:18.54" />
                    <SPLIT distance="500" swimtime="00:08:45.75" />
                    <SPLIT distance="525" swimtime="00:09:13.00" />
                    <SPLIT distance="550" swimtime="00:09:40.56" />
                    <SPLIT distance="575" swimtime="00:10:08.29" />
                    <SPLIT distance="600" swimtime="00:10:35.85" />
                    <SPLIT distance="625" swimtime="00:11:03.22" />
                    <SPLIT distance="650" swimtime="00:11:30.72" />
                    <SPLIT distance="675" swimtime="00:11:58.33" />
                    <SPLIT distance="700" swimtime="00:12:25.43" />
                    <SPLIT distance="725" swimtime="00:12:52.51" />
                    <SPLIT distance="750" swimtime="00:13:19.73" />
                    <SPLIT distance="775" swimtime="00:13:45.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="208" reactiontime="+82" swimtime="00:01:25.90" resultid="109978" heatid="110672" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.46" />
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="75" swimtime="00:01:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="212" reactiontime="+91" swimtime="00:01:44.46" resultid="109979" heatid="110722" lane="5" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.43" />
                    <SPLIT distance="50" swimtime="00:00:50.30" />
                    <SPLIT distance="75" swimtime="00:01:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="175" swimtime="00:03:18.04" resultid="109980" heatid="110766" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.39" />
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                    <SPLIT distance="75" swimtime="00:01:08.17" />
                    <SPLIT distance="100" swimtime="00:01:33.92" />
                    <SPLIT distance="125" swimtime="00:02:00.25" />
                    <SPLIT distance="150" swimtime="00:02:26.56" />
                    <SPLIT distance="175" swimtime="00:02:53.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="184" reactiontime="+93" swimtime="00:06:51.73" resultid="109981" heatid="110841" lane="7" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.54" />
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                    <SPLIT distance="75" swimtime="00:01:07.54" />
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                    <SPLIT distance="125" swimtime="00:01:57.78" />
                    <SPLIT distance="150" swimtime="00:02:23.90" />
                    <SPLIT distance="175" swimtime="00:02:50.07" />
                    <SPLIT distance="200" swimtime="00:03:17.47" />
                    <SPLIT distance="225" swimtime="00:03:43.51" />
                    <SPLIT distance="250" swimtime="00:04:11.30" />
                    <SPLIT distance="275" swimtime="00:04:38.76" />
                    <SPLIT distance="300" swimtime="00:05:05.65" />
                    <SPLIT distance="325" swimtime="00:05:33.03" />
                    <SPLIT distance="350" swimtime="00:06:00.05" />
                    <SPLIT distance="375" swimtime="00:06:26.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="99059" points="239" reactiontime="+87" swimtime="00:02:25.82" resultid="110004" heatid="110716" lane="2">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.50" />
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="75" swimtime="00:00:51.86" />
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                    <SPLIT distance="125" swimtime="00:01:31.28" />
                    <SPLIT distance="150" swimtime="00:01:55.58" />
                    <SPLIT distance="175" swimtime="00:02:10.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109939" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="109964" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="109958" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="109830" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="99059" points="393" reactiontime="+90" swimtime="00:02:03.48" resultid="110005" heatid="110718" lane="4" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.90" />
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="75" swimtime="00:00:50.64" />
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="125" swimtime="00:01:21.74" />
                    <SPLIT distance="150" swimtime="00:01:36.69" />
                    <SPLIT distance="175" swimtime="00:01:49.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109844" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="109951" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="109862" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="109932" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="99059" points="276" reactiontime="+92" swimtime="00:02:18.97" resultid="110006" heatid="110717" lane="1" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.34" />
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="75" swimtime="00:00:54.82" />
                    <SPLIT distance="100" swimtime="00:01:16.17" />
                    <SPLIT distance="125" swimtime="00:01:31.39" />
                    <SPLIT distance="150" swimtime="00:01:49.66" />
                    <SPLIT distance="175" swimtime="00:02:03.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109942" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="109853" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="109880" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="109972" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="10">
              <RESULTS>
                <RESULT eventid="99250" points="305" reactiontime="+67" swimtime="00:02:02.70" resultid="110010" heatid="110782" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                    <SPLIT distance="75" swimtime="00:01:16.71" />
                    <SPLIT distance="100" swimtime="00:01:00.49" />
                    <SPLIT distance="150" swimtime="00:01:34.50" />
                    <SPLIT distance="175" swimtime="00:01:47.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109830" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="109841" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="109958" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="109939" number="4" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="11">
              <RESULTS>
                <RESULT eventid="99250" points="506" reactiontime="+79" swimtime="00:01:43.62" resultid="110009" heatid="110784" lane="1" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.64" />
                    <SPLIT distance="50" swimtime="00:00:25.82" />
                    <SPLIT distance="75" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:00:52.14" />
                    <SPLIT distance="125" swimtime="00:01:05.30" />
                    <SPLIT distance="150" swimtime="00:01:19.14" />
                    <SPLIT distance="175" swimtime="00:01:30.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109862" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="109951" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="109932" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="109887" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="12">
              <RESULTS>
                <RESULT eventid="99250" points="309" reactiontime="+77" swimtime="00:02:02.08" resultid="110011" heatid="110783" lane="8" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.81" />
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="75" swimtime="00:00:47.06" />
                    <SPLIT distance="100" swimtime="00:01:02.54" />
                    <SPLIT distance="125" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:01:32.96" />
                    <SPLIT distance="175" swimtime="00:01:46.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109964" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="109880" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="109942" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="109844" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="13">
              <RESULTS>
                <RESULT eventid="99250" points="182" reactiontime="+102" swimtime="00:02:25.71" resultid="110012" heatid="110781" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.87" />
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="75" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:01.55" />
                    <SPLIT distance="125" swimtime="00:01:19.41" />
                    <SPLIT distance="150" swimtime="00:01:41.03" />
                    <SPLIT distance="175" swimtime="00:02:02.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109972" number="1" reactiontime="+102" />
                    <RELAYPOSITION athleteid="109853" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="109982" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="109813" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="99036" points="355" reactiontime="+90" swimtime="00:02:26.80" resultid="110002" heatid="110715" lane="1" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.49" />
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="75" swimtime="00:00:57.10" />
                    <SPLIT distance="100" swimtime="00:01:20.22" />
                    <SPLIT distance="125" swimtime="00:01:34.71" />
                    <SPLIT distance="150" swimtime="00:01:52.35" />
                    <SPLIT distance="175" swimtime="00:02:08.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109925" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="109920" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="109985" number="3" reactiontime="-2" />
                    <RELAYPOSITION athleteid="109821" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="5">
              <RESULTS>
                <RESULT eventid="99036" points="198" reactiontime="+78" swimtime="00:02:58.50" resultid="110003" heatid="110714" lane="4">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.89" />
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                    <SPLIT distance="75" swimtime="00:01:08.92" />
                    <SPLIT distance="100" swimtime="00:01:39.84" />
                    <SPLIT distance="125" swimtime="00:01:58.02" />
                    <SPLIT distance="150" swimtime="00:02:20.08" />
                    <SPLIT distance="175" swimtime="00:02:38.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109836" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="109907" number="2" />
                    <RELAYPOSITION athleteid="109871" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="109976" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="9">
              <RESULTS>
                <RESULT eventid="99234" points="377" reactiontime="+90" swimtime="00:02:10.39" resultid="110007" heatid="110780" lane="1" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.60" />
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="75" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:02.86" />
                    <SPLIT distance="125" swimtime="00:01:19.50" />
                    <SPLIT distance="150" swimtime="00:01:37.35" />
                    <SPLIT distance="175" swimtime="00:01:53.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109925" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="109985" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="109871" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="109920" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="10">
              <RESULTS>
                <RESULT eventid="99234" points="137" reactiontime="+92" swimtime="00:03:02.50" resultid="110008" heatid="110779" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.27" />
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="75" swimtime="00:00:56.44" />
                    <SPLIT distance="100" swimtime="00:01:14.98" />
                    <SPLIT distance="125" swimtime="00:01:43.61" />
                    <SPLIT distance="150" swimtime="00:02:16.11" />
                    <SPLIT distance="175" swimtime="00:02:38.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109976" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="109836" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="109907" number="3" />
                    <RELAYPOSITION athleteid="109911" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="397" reactiontime="+58" swimtime="00:01:52.32" resultid="109998" heatid="110631" lane="5" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:55.96" />
                    <SPLIT distance="75" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:26.68" />
                    <SPLIT distance="125" swimtime="00:01:10.65" />
                    <SPLIT distance="175" swimtime="00:01:39.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109887" number="1" reactiontime="+58" />
                    <RELAYPOSITION athleteid="109925" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="109985" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="109862" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="253" swimtime="00:02:10.56" resultid="110000" heatid="110631" lane="9" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="75" swimtime="00:00:44.18" />
                    <SPLIT distance="100" swimtime="00:01:02.67" />
                    <SPLIT distance="125" swimtime="00:01:21.06" />
                    <SPLIT distance="150" swimtime="00:01:39.90" />
                    <SPLIT distance="175" swimtime="00:01:54.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109932" number="1" />
                    <RELAYPOSITION athleteid="109821" number="2" />
                    <RELAYPOSITION athleteid="109976" number="3" />
                    <RELAYPOSITION athleteid="109844" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="98846" points="77" swimtime="00:03:13.96" resultid="110001" heatid="110629" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.40" />
                    <SPLIT distance="75" swimtime="00:01:22.35" />
                    <SPLIT distance="100" swimtime="00:01:47.34" />
                    <SPLIT distance="125" swimtime="00:02:07.93" />
                    <SPLIT distance="150" swimtime="00:02:28.32" />
                    <SPLIT distance="175" swimtime="00:02:49.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109907" number="1" />
                    <RELAYPOSITION athleteid="109911" number="2" />
                    <RELAYPOSITION athleteid="109982" number="3" reactiontime="+81" />
                    <RELAYPOSITION athleteid="109813" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="98846" points="281" reactiontime="+97" swimtime="00:02:06.00" resultid="109999" heatid="110631" lane="1" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.04" />
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="75" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:00.08" />
                    <SPLIT distance="125" swimtime="00:01:16.46" />
                    <SPLIT distance="150" swimtime="00:01:33.78" />
                    <SPLIT distance="175" swimtime="00:01:49.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109951" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="109972" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="109871" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="109920" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="13">
              <RESULTS>
                <RESULT eventid="99441" points="374" reactiontime="+74" swimtime="00:02:05.56" resultid="110013" heatid="110837" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.45" />
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="75" swimtime="00:00:52.01" />
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                    <SPLIT distance="125" swimtime="00:01:23.95" />
                    <SPLIT distance="150" swimtime="00:01:41.46" />
                    <SPLIT distance="175" swimtime="00:01:53.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109925" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="109951" number="2" />
                    <RELAYPOSITION athleteid="109985" number="3" />
                    <RELAYPOSITION athleteid="109887" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="14">
              <RESULTS>
                <RESULT eventid="99441" points="235" reactiontime="+83" swimtime="00:02:26.61" resultid="110015" heatid="110837" lane="0" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="75" swimtime="00:00:56.96" />
                    <SPLIT distance="100" swimtime="00:01:51.93" />
                    <SPLIT distance="125" swimtime="00:01:36.27" />
                    <SPLIT distance="175" swimtime="00:02:08.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109844" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="109976" number="2" />
                    <RELAYPOSITION athleteid="109862" number="3" />
                    <RELAYPOSITION athleteid="109821" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="15">
              <RESULTS>
                <RESULT eventid="99441" points="238" reactiontime="+88" swimtime="00:02:25.97" resultid="110014" heatid="110836" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.75" />
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="75" swimtime="00:00:54.13" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="125" swimtime="00:01:34.04" />
                    <SPLIT distance="150" swimtime="00:01:55.49" />
                    <SPLIT distance="175" swimtime="00:02:10.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109942" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="109920" number="2" />
                    <RELAYPOSITION athleteid="109871" number="3" />
                    <RELAYPOSITION athleteid="109853" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="109325" name="AquaStars Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1978-01-01" firstname=" MARIUSZ" gender="M" lastname="GOLON " nation="POL" athleteid="109277" lastname.en="GOLON">
              <RESULTS>
                <RESULT eventid="98830" points="333" swimtime="00:02:38.11" resultid="109606" heatid="110621" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.70" />
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="75" swimtime="00:00:51.42" />
                    <SPLIT distance="100" swimtime="00:01:11.75" />
                    <SPLIT distance="125" swimtime="00:01:36.04" />
                    <SPLIT distance="150" swimtime="00:02:00.08" />
                    <SPLIT distance="175" swimtime="00:02:20.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="109607" heatid="110639" lane="3" entrytime="00:12:00.00" />
                <RESULT eventid="98924" points="319" reactiontime="+80" swimtime="00:00:32.50" resultid="109608" heatid="110654" lane="5" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="413" reactiontime="+78" swimtime="00:01:07.98" resultid="109609" heatid="110699" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="75" swimtime="00:00:50.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="377" reactiontime="+69" swimtime="00:01:16.95" resultid="109610" heatid="110727" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.65" />
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="75" swimtime="00:00:55.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="444" swimtime="00:00:28.56" resultid="109611" heatid="110746" lane="0" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="434" swimtime="00:00:33.35" resultid="109612" heatid="110827" lane="0" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="ŚLĄSK" clubid="109315" name="AZS PWSZ RACIBÓRZ">
          <CONTACT city="racibórz" email="adip45@poczta.onet.pl" name="Piechula Adolf" phone="606 114 286" state="ŚLĄSK" street="słowackiego55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-04-11" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" swrid="4992724" athleteid="109316">
              <RESULTS>
                <RESULT eventid="98830" points="200" reactiontime="+92" swimtime="00:03:07.43" resultid="109317" heatid="110622" lane="6" entrytime="00:03:04.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.40" />
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="75" swimtime="00:01:01.36" />
                    <SPLIT distance="100" swimtime="00:01:25.40" />
                    <SPLIT distance="125" swimtime="00:01:53.92" />
                    <SPLIT distance="150" swimtime="00:02:22.21" />
                    <SPLIT distance="175" swimtime="00:02:45.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="173" reactiontime="+112" swimtime="00:13:15.70" resultid="109318" heatid="110637" lane="0" entrytime="00:12:56.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.88" />
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="75" swimtime="00:01:48.58" />
                    <SPLIT distance="100" swimtime="00:01:24.79" />
                    <SPLIT distance="125" swimtime="00:02:35.47" />
                    <SPLIT distance="150" swimtime="00:02:11.49" />
                    <SPLIT distance="175" swimtime="00:03:24.21" />
                    <SPLIT distance="200" swimtime="00:02:59.66" />
                    <SPLIT distance="225" swimtime="00:04:13.31" />
                    <SPLIT distance="250" swimtime="00:03:48.62" />
                    <SPLIT distance="275" swimtime="00:05:02.94" />
                    <SPLIT distance="300" swimtime="00:04:38.01" />
                    <SPLIT distance="325" swimtime="00:05:53.24" />
                    <SPLIT distance="350" swimtime="00:05:27.70" />
                    <SPLIT distance="375" swimtime="00:06:43.79" />
                    <SPLIT distance="400" swimtime="00:06:18.39" />
                    <SPLIT distance="425" swimtime="00:07:36.45" />
                    <SPLIT distance="450" swimtime="00:07:08.86" />
                    <SPLIT distance="475" swimtime="00:08:27.61" />
                    <SPLIT distance="500" swimtime="00:08:01.64" />
                    <SPLIT distance="525" swimtime="00:09:20.79" />
                    <SPLIT distance="550" swimtime="00:08:54.72" />
                    <SPLIT distance="575" swimtime="00:10:13.73" />
                    <SPLIT distance="600" swimtime="00:09:47.43" />
                    <SPLIT distance="625" swimtime="00:11:06.46" />
                    <SPLIT distance="650" swimtime="00:10:40.63" />
                    <SPLIT distance="675" swimtime="00:11:58.94" />
                    <SPLIT distance="700" swimtime="00:11:32.81" />
                    <SPLIT distance="725" swimtime="00:12:51.07" />
                    <SPLIT distance="750" swimtime="00:12:25.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="209" reactiontime="+104" swimtime="00:03:22.70" resultid="109319" heatid="110667" lane="6" entrytime="00:03:18.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.22" />
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="75" swimtime="00:01:09.62" />
                    <SPLIT distance="100" swimtime="00:01:35.70" />
                    <SPLIT distance="125" swimtime="00:02:02.05" />
                    <SPLIT distance="150" swimtime="00:02:29.16" />
                    <SPLIT distance="175" swimtime="00:02:56.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="171" reactiontime="+105" swimtime="00:03:15.53" resultid="109320" heatid="110711" lane="5" entrytime="00:03:10.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.87" />
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="75" swimtime="00:01:07.46" />
                    <SPLIT distance="100" swimtime="00:01:32.74" />
                    <SPLIT distance="125" swimtime="00:01:58.60" />
                    <SPLIT distance="150" swimtime="00:02:24.77" />
                    <SPLIT distance="175" swimtime="00:02:50.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="186" swimtime="00:06:52.42" resultid="109322" heatid="110790" lane="9" entrytime="00:06:28.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.65" />
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                    <SPLIT distance="75" swimtime="00:01:06.40" />
                    <SPLIT distance="100" swimtime="00:01:32.33" />
                    <SPLIT distance="125" swimtime="00:01:59.09" />
                    <SPLIT distance="150" swimtime="00:02:26.48" />
                    <SPLIT distance="175" swimtime="00:02:53.66" />
                    <SPLIT distance="200" swimtime="00:03:19.63" />
                    <SPLIT distance="225" swimtime="00:03:48.83" />
                    <SPLIT distance="250" swimtime="00:04:17.83" />
                    <SPLIT distance="275" swimtime="00:04:46.63" />
                    <SPLIT distance="300" swimtime="00:05:15.37" />
                    <SPLIT distance="325" swimtime="00:05:38.87" />
                    <SPLIT distance="350" swimtime="00:06:03.53" />
                    <SPLIT distance="375" swimtime="00:06:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="183" swimtime="00:01:25.29" resultid="109323" heatid="110800" lane="6" entrytime="00:01:24.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.85" />
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                    <SPLIT distance="75" swimtime="00:00:59.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="274" swimtime="00:00:38.83" resultid="109324" heatid="110828" lane="2" entrytime="00:00:39.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="224" reactiontime="+93" swimtime="00:01:31.51" resultid="110862" heatid="110730" lane="5" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.70" />
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                    <SPLIT distance="75" swimtime="00:01:06.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="BLR" clubid="109210" name="BELARUS">
          <ATHLETES>
            <ATHLETE birthdate="1995-05-05" firstname="Yauheni" gender="M" lastname="PUZAN " nation="BLR" athleteid="109211">
              <RESULTS>
                <RESULT eventid="98798" points="533" reactiontime="+74" swimtime="00:00:24.98" resultid="109212" heatid="110612" lane="3" entrytime="00:00:24.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="496" reactiontime="+77" swimtime="00:00:56.77" resultid="109213" heatid="110689" lane="1" entrytime="00:00:55.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                    <SPLIT distance="75" swimtime="00:00:42.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="602" reactiontime="+42" swimtime="00:00:25.81" resultid="109214" heatid="110751" lane="2" entrytime="00:00:25.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="543" reactiontime="+74" swimtime="00:00:59.36" resultid="109215" heatid="110805" lane="3" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.13" />
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                    <SPLIT distance="75" swimtime="00:00:42.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="110217" name="DELFIN Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="JAKUB" gender="M" lastname="MAŃCZAK" nation="POL" swrid="4186188" athleteid="108927">
              <RESULTS>
                <RESULT eventid="99170" reactiontime="+49" status="DNF" swimtime="00:00:00.00" resultid="108928" heatid="110748" lane="4" entrytime="00:00:29.40" entrycourse="SCM" />
                <RESULT eventid="99361" points="335" reactiontime="+90" swimtime="00:01:09.71" resultid="108929" heatid="110803" lane="2" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.95" />
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="75" swimtime="00:00:51.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="289" swimtime="00:02:44.14" resultid="108930" heatid="110712" lane="2" entrytime="00:02:55.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.94" />
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="75" swimtime="00:00:56.85" />
                    <SPLIT distance="100" swimtime="00:01:18.31" />
                    <SPLIT distance="125" swimtime="00:01:40.30" />
                    <SPLIT distance="150" swimtime="00:02:02.60" />
                    <SPLIT distance="175" swimtime="00:02:24.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="372" swimtime="00:02:18.10" resultid="108931" heatid="110775" lane="6" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="75" swimtime="00:00:49.11" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="125" swimtime="00:01:24.54" />
                    <SPLIT distance="150" swimtime="00:01:42.75" />
                    <SPLIT distance="175" swimtime="00:02:01.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="107779" name="Dynamo">
          <CONTACT city="Kharkiv" email="swimmer2003@ukr.net" name="Vadym Kutsenko" phone="+38 057 7204282" street="16 Novgorodska" zip="61165" />
          <ATHLETES>
            <ATHLETE birthdate="1945-05-05" firstname="Vadym" gender="M" lastname="Kutsenko" nation="UKR" athleteid="107780">
              <RESULTS>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="107782" heatid="110698" lane="4" entrytime="00:01:21.14" entrycourse="SCM" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="107783" heatid="110774" lane="1" entrytime="00:02:28.53" entrycourse="SCM" />
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="107784" heatid="110789" lane="6" entrytime="00:06:49.52" entrycourse="LCM" />
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="107785" heatid="110847" lane="9" entrytime="00:05:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="108449" name="Gdynia Masters">
          <CONTACT email="k.mysiak@wpit.am.gdynia.pl" name="Mysiak Katarzyna" />
          <ATHLETES>
            <ATHLETE birthdate="1952-01-01" firstname="Barbara" gender="F" lastname="Chomicka" nation="POL" athleteid="108460">
              <RESULTS>
                <RESULT eventid="106294" points="96" reactiontime="+79" swimtime="00:00:56.04" resultid="108461" heatid="110646" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="48" reactiontime="+102" swimtime="00:05:27.18" resultid="108462" heatid="110707" lane="2" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.09" />
                    <SPLIT distance="50" swimtime="00:01:13.57" />
                    <SPLIT distance="75" swimtime="00:01:55.14" />
                    <SPLIT distance="100" swimtime="00:02:38.87" />
                    <SPLIT distance="125" swimtime="00:03:20.49" />
                    <SPLIT distance="150" swimtime="00:04:03.36" />
                    <SPLIT distance="175" swimtime="00:04:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="54" reactiontime="+104" swimtime="00:01:04.44" resultid="108463" heatid="110736" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="87" reactiontime="+75" swimtime="00:02:03.93" resultid="108464" heatid="110753" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="75" swimtime="00:01:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="48" reactiontime="+105" swimtime="00:02:30.03" resultid="108465" heatid="110793" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.04" />
                    <SPLIT distance="50" swimtime="00:01:09.46" />
                    <SPLIT distance="75" swimtime="00:01:50.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="83" reactiontime="+79" swimtime="00:04:32.85" resultid="108466" heatid="110806" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.70" />
                    <SPLIT distance="50" swimtime="00:01:01.97" />
                    <SPLIT distance="100" swimtime="00:02:08.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Grażyna" gender="F" lastname="Heisler" nation="POL" athleteid="108467">
              <RESULTS>
                <RESULT eventid="98777" points="158" reactiontime="+97" swimtime="00:00:42.94" resultid="108468" heatid="110587" lane="8" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="90" reactiontime="+87" swimtime="00:00:57.16" resultid="108469" heatid="110647" lane="9" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="111" swimtime="00:01:57.88" resultid="108470" heatid="110691" lane="9" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.82" />
                    <SPLIT distance="50" swimtime="00:00:54.24" />
                    <SPLIT distance="75" swimtime="00:01:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="125" reactiontime="+75" swimtime="00:02:04.46" resultid="108471" heatid="110721" lane="5" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.79" />
                    <SPLIT distance="50" swimtime="00:00:57.52" />
                    <SPLIT distance="75" swimtime="00:01:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="81" reactiontime="+43" swimtime="00:02:07.03" resultid="108472" heatid="110754" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.10" />
                    <SPLIT distance="50" swimtime="00:00:59.36" />
                    <SPLIT distance="75" swimtime="00:01:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="126" reactiontime="+109" swimtime="00:00:57.33" resultid="108473" heatid="110818" lane="1" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="108478">
              <RESULTS>
                <RESULT eventid="98798" points="116" reactiontime="+120" swimtime="00:00:41.53" resultid="108479" heatid="110597" lane="1" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="85" reactiontime="+108" swimtime="00:04:08.83" resultid="108480" heatid="110620" lane="0" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.48" />
                    <SPLIT distance="50" swimtime="00:01:00.10" />
                    <SPLIT distance="75" swimtime="00:01:33.67" />
                    <SPLIT distance="100" swimtime="00:02:08.19" />
                    <SPLIT distance="125" swimtime="00:02:41.62" />
                    <SPLIT distance="150" swimtime="00:03:15.01" />
                    <SPLIT distance="175" swimtime="00:03:42.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="89" reactiontime="+102" swimtime="00:00:49.63" resultid="108481" heatid="110653" lane="9" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="106" swimtime="00:01:47.04" resultid="108482" heatid="110697" lane="9" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.40" />
                    <SPLIT distance="50" swimtime="00:00:51.75" />
                    <SPLIT distance="75" swimtime="00:01:22.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="108" swimtime="00:01:56.60" resultid="108483" heatid="110728" lane="9" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.88" />
                    <SPLIT distance="50" swimtime="00:00:53.11" />
                    <SPLIT distance="75" swimtime="00:01:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="91" swimtime="00:03:40.32" resultid="108484" heatid="110770" lane="9" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.85" />
                    <SPLIT distance="50" swimtime="00:00:48.03" />
                    <SPLIT distance="75" swimtime="00:01:14.87" />
                    <SPLIT distance="100" swimtime="00:01:43.93" />
                    <SPLIT distance="125" swimtime="00:02:12.31" />
                    <SPLIT distance="150" swimtime="00:02:43.04" />
                    <SPLIT distance="175" swimtime="00:03:11.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="153" reactiontime="+111" swimtime="00:00:47.16" resultid="108485" heatid="110825" lane="4" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="108486">
              <RESULTS>
                <RESULT eventid="98924" points="81" reactiontime="+107" swimtime="00:00:51.30" resultid="108487" heatid="110653" lane="0" entrytime="00:00:49.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="97" swimtime="00:02:00.75" resultid="108488" heatid="110728" lane="0" entrytime="00:01:52.42">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.60" />
                    <SPLIT distance="50" swimtime="00:00:58.22" />
                    <SPLIT distance="75" swimtime="00:01:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="76" reactiontime="+87" swimtime="00:01:55.10" resultid="108489" heatid="110758" lane="7" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.67" />
                    <SPLIT distance="50" swimtime="00:00:53.64" />
                    <SPLIT distance="75" swimtime="00:01:23.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="100" swimtime="00:00:54.23" resultid="108490" heatid="110825" lane="2" entrytime="00:00:49.51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Katarzyna" gender="F" lastname="Mysiak" nation="POL" athleteid="108453">
              <RESULTS>
                <RESULT eventid="98777" points="216" reactiontime="+96" swimtime="00:00:38.72" resultid="108454" heatid="110587" lane="3" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="138" reactiontime="+87" swimtime="00:00:49.63" resultid="108455" heatid="110648" lane="0" entrytime="00:00:44.00" />
                <RESULT eventid="98907" points="173" reactiontime="+107" swimtime="00:01:31.32" resultid="108456" heatid="110672" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.30" />
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="75" swimtime="00:01:06.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="140" reactiontime="+80" swimtime="00:01:45.96" resultid="108457" heatid="110754" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.11" />
                    <SPLIT distance="75" swimtime="00:01:19.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="161" reactiontime="+99" swimtime="00:03:23.38" resultid="108458" heatid="110765" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.27" />
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                    <SPLIT distance="75" swimtime="00:01:10.66" />
                    <SPLIT distance="100" swimtime="00:01:37.19" />
                    <SPLIT distance="125" swimtime="00:02:04.18" />
                    <SPLIT distance="150" swimtime="00:02:31.36" />
                    <SPLIT distance="175" swimtime="00:02:58.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="176" reactiontime="+122" swimtime="00:06:58.46" resultid="108459" heatid="110842" lane="3" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.00" />
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                    <SPLIT distance="75" swimtime="00:01:13.06" />
                    <SPLIT distance="100" swimtime="00:01:39.97" />
                    <SPLIT distance="125" swimtime="00:03:00.88" />
                    <SPLIT distance="150" swimtime="00:02:33.45" />
                    <SPLIT distance="175" swimtime="00:03:55.25" />
                    <SPLIT distance="200" swimtime="00:03:28.15" />
                    <SPLIT distance="225" swimtime="00:04:49.52" />
                    <SPLIT distance="250" swimtime="00:04:22.64" />
                    <SPLIT distance="275" swimtime="00:05:43.03" />
                    <SPLIT distance="300" swimtime="00:05:16.80" />
                    <SPLIT distance="325" swimtime="00:06:35.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="108474">
              <RESULTS>
                <RESULT eventid="98956" points="204" swimtime="00:03:24.55" resultid="108475" heatid="110667" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.80" />
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                    <SPLIT distance="75" swimtime="00:01:10.22" />
                    <SPLIT distance="100" swimtime="00:01:36.88" />
                    <SPLIT distance="125" swimtime="00:02:04.43" />
                    <SPLIT distance="150" swimtime="00:02:32.90" />
                    <SPLIT distance="175" swimtime="00:02:58.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="241" swimtime="00:01:29.26" resultid="108476" heatid="110730" lane="0" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.18" />
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                    <SPLIT distance="75" swimtime="00:01:05.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="249" reactiontime="+103" swimtime="00:00:40.11" resultid="108477" heatid="110827" lane="1" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="141" reactiontime="+99" swimtime="00:02:38.45" resultid="108491" heatid="110629" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.25" />
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="75" swimtime="00:00:57.16" />
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="125" swimtime="00:01:38.53" />
                    <SPLIT distance="150" swimtime="00:02:01.92" />
                    <SPLIT distance="175" swimtime="00:02:19.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108453" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="108474" number="2" reactiontime="+6" />
                    <RELAYPOSITION athleteid="108467" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="108478" number="4" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="99441" points="70" reactiontime="+72" swimtime="00:03:39.05" resultid="108492" heatid="110835" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.03" />
                    <SPLIT distance="50" swimtime="00:00:57.17" />
                    <SPLIT distance="75" swimtime="00:01:22.71" />
                    <SPLIT distance="100" swimtime="00:01:17.26" />
                    <SPLIT distance="125" swimtime="00:02:21.96" />
                    <SPLIT distance="150" swimtime="00:02:57.02" />
                    <SPLIT distance="175" swimtime="00:03:15.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108467" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="108486" number="2" />
                    <RELAYPOSITION athleteid="108460" number="3" />
                    <RELAYPOSITION athleteid="108478" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="SWE" clubid="106403" name="Göteborg SIM">
          <ATHLETES>
            <ATHLETE birthdate="1951-05-11" firstname="LEONARD" gender="M" lastname="BIELICZ" nation="SWE" athleteid="106404">
              <RESULTS>
                <RESULT eventid="98798" points="392" reactiontime="+76" swimtime="00:00:27.66" resultid="106405" heatid="110608" lane="3" entrytime="00:00:27.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="394" reactiontime="+75" swimtime="00:01:01.28" resultid="106406" heatid="110686" lane="6" entrytime="00:01:01.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.00" />
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                    <SPLIT distance="75" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="407" swimtime="00:00:29.41" resultid="106407" heatid="110748" lane="6" entrytime="00:00:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="344" reactiontime="+78" swimtime="00:01:09.07" resultid="106408" heatid="110803" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.57" />
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="75" swimtime="00:00:49.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="108368" name="IKS Konstancin">
          <CONTACT name="Obiedziński" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" license="103714700078" athleteid="108369">
              <RESULTS>
                <RESULT eventid="98798" points="413" reactiontime="+79" swimtime="00:00:27.20" resultid="108370" heatid="110607" lane="2" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="318" reactiontime="+82" swimtime="00:02:40.59" resultid="108371" heatid="110625" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.39" />
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="75" swimtime="00:00:54.72" />
                    <SPLIT distance="100" swimtime="00:01:16.23" />
                    <SPLIT distance="125" swimtime="00:01:39.72" />
                    <SPLIT distance="150" swimtime="00:02:03.78" />
                    <SPLIT distance="175" swimtime="00:02:23.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="435" reactiontime="+74" swimtime="00:00:59.28" resultid="108372" heatid="110686" lane="4" entrytime="00:01:00.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                    <SPLIT distance="75" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="346" swimtime="00:01:12.14" resultid="108373" heatid="110702" lane="9" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.08" />
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="75" swimtime="00:00:55.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="319" reactiontime="+89" swimtime="00:01:21.35" resultid="108374" heatid="110731" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.60" />
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="75" swimtime="00:00:59.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="359" swimtime="00:00:30.66" resultid="108375" heatid="110747" lane="6" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="108376" heatid="110802" lane="9" entrytime="00:01:15.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="108377" heatid="110829" lane="6" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="108378" name="Kauno Takas">
          <CONTACT city="Kaunas" email="abicka@takas.lt" internet="klubastakas.lt" name="Ramune Ivanauskaite" phone="+37068297778" street="Lentvario g. 19" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1961-05-07" firstname="Jolanta" gender="F" lastname="Kozak" nation="LTU" athleteid="108393">
              <RESULTS>
                <RESULT eventid="98777" points="104" status="DNS" swimtime="00:00:49.32" resultid="108394" heatid="110586" lane="2" entrytime="00:00:58.00" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="108395" heatid="110672" lane="8" entrytime="00:01:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-14" firstname="Violeta" gender="F" lastname="Penkauskaite" nation="LTU" athleteid="108388">
              <RESULTS>
                <RESULT eventid="106294" status="DNS" swimtime="00:00:00.00" resultid="108389" heatid="110646" lane="3" entrytime="00:00:55.30" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="108390" heatid="110690" lane="4" entrytime="00:01:59.30" />
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="108391" heatid="110754" lane="2" entrytime="00:01:49.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="108392" heatid="110818" lane="7" entrytime="00:00:58.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-11-16" firstname="Violeta" gender="F" lastname="Povilaitiene" nation="LTU" athleteid="108384">
              <RESULTS>
                <RESULT eventid="98777" points="101" status="DNS" swimtime="00:00:49.89" resultid="108385" heatid="110586" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="98940" status="DNS" swimtime="00:00:00.00" resultid="108386" heatid="110661" lane="3" entrytime="00:04:30.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="108387" heatid="110818" lane="3" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-10-18" firstname="Ramune" gender="F" lastname="Ivanauskaite" nation="LTU" athleteid="108379">
              <RESULTS>
                <RESULT eventid="106294" points="198" reactiontime="+110" swimtime="00:00:44.01" resultid="108380" heatid="110648" lane="7" entrytime="00:00:42.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="239" reactiontime="+77" swimtime="00:03:36.78" resultid="108381" heatid="110662" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.25" />
                    <SPLIT distance="50" swimtime="00:00:50.32" />
                    <SPLIT distance="75" swimtime="00:01:17.41" />
                    <SPLIT distance="100" swimtime="00:01:44.41" />
                    <SPLIT distance="125" swimtime="00:02:12.10" />
                    <SPLIT distance="150" swimtime="00:02:39.95" />
                    <SPLIT distance="175" swimtime="00:03:08.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="226" reactiontime="+97" swimtime="00:01:30.27" resultid="108382" heatid="110755" lane="9" entrytime="00:01:33.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.60" />
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="75" swimtime="00:01:07.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="240" reactiontime="+101" swimtime="00:03:11.82" resultid="108383" heatid="110808" lane="9" entrytime="00:03:15.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.91" />
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                    <SPLIT distance="75" swimtime="00:01:09.51" />
                    <SPLIT distance="100" swimtime="00:01:33.54" />
                    <SPLIT distance="125" swimtime="00:01:58.06" />
                    <SPLIT distance="150" swimtime="00:02:22.60" />
                    <SPLIT distance="175" swimtime="00:02:48.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" region="KLAIPEDA" clubid="107828" name="Klaipeda Swimming Club">
          <CONTACT email="klaipeda.swimming@gmail.com" name="Tomas Zemaitis" phone="+37065244408" />
          <ATHLETES>
            <ATHLETE birthdate="1989-04-22" firstname="Martynas" gender="M" lastname="Laucka" nation="LTU" athleteid="107847">
              <RESULTS>
                <RESULT eventid="98798" points="423" reactiontime="+85" swimtime="00:00:26.97" resultid="107848" heatid="110609" lane="0" entrytime="00:00:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="402" swimtime="00:01:00.88" resultid="107849" heatid="110687" lane="2" entrytime="00:00:59.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.50" />
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="75" swimtime="00:00:45.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="328" reactiontime="+74" swimtime="00:01:20.56" resultid="107850" heatid="110732" lane="5" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.61" />
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="75" swimtime="00:00:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="320" reactiontime="+68" swimtime="00:02:25.14" resultid="107851" heatid="110774" lane="4" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.51" />
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="75" swimtime="00:00:51.28" />
                    <SPLIT distance="100" swimtime="00:01:09.86" />
                    <SPLIT distance="125" swimtime="00:01:29.19" />
                    <SPLIT distance="150" swimtime="00:01:48.81" />
                    <SPLIT distance="175" swimtime="00:02:07.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="297" reactiontime="+83" swimtime="00:00:37.83" resultid="107852" heatid="110832" lane="3" entrytime="00:00:34.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-04-10" firstname="Aidas" gender="M" lastname="Pelesinas" nation="LTU" athleteid="107842">
              <RESULTS>
                <RESULT eventid="98798" points="465" swimtime="00:00:26.15" resultid="107843" heatid="110609" lane="9" entrytime="00:00:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="426" swimtime="00:00:59.69" resultid="107844" heatid="110687" lane="0" entrytime="00:01:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="75" swimtime="00:00:44.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="327" reactiontime="+98" swimtime="00:00:31.63" resultid="107845" heatid="110746" lane="2" entrytime="00:00:31.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="420" swimtime="00:00:33.71" resultid="107846" heatid="110832" lane="9" entrytime="00:00:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-26" firstname="Ausra" gender="F" lastname="Gardziuliene" nation="LTU" athleteid="107853">
              <RESULTS>
                <RESULT eventid="98777" points="346" reactiontime="+94" swimtime="00:00:33.10" resultid="107854" heatid="110590" lane="2" entrytime="00:00:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="303" reactiontime="+91" swimtime="00:03:20.29" resultid="107855" heatid="110663" lane="5" entrytime="00:03:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.60" />
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="75" swimtime="00:01:09.75" />
                    <SPLIT distance="100" swimtime="00:01:35.09" />
                    <SPLIT distance="125" swimtime="00:02:01.30" />
                    <SPLIT distance="150" swimtime="00:02:27.68" />
                    <SPLIT distance="175" swimtime="00:02:54.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="272" swimtime="00:01:27.46" resultid="107856" heatid="110693" lane="9" entrytime="00:01:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.80" />
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="75" swimtime="00:01:05.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="331" reactiontime="+90" swimtime="00:01:30.14" resultid="107857" heatid="110724" lane="7" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.49" />
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="75" swimtime="00:01:05.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="276" reactiontime="+95" swimtime="00:00:37.42" resultid="107858" heatid="110738" lane="7" entrytime="00:00:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="347" swimtime="00:00:40.97" resultid="107859" heatid="110821" lane="6" entrytime="00:00:40.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-02-25" firstname="Arturas" gender="M" lastname="Klimas" nation="LTU" athleteid="107865">
              <RESULTS>
                <RESULT eventid="98798" points="319" reactiontime="+87" swimtime="00:00:29.63" resultid="107866" heatid="110605" lane="8" entrytime="00:00:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="319" swimtime="00:01:05.76" resultid="107867" heatid="110683" lane="6" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.08" />
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="75" swimtime="00:00:48.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="293" reactiontime="+92" swimtime="00:00:32.79" resultid="107868" heatid="110746" lane="8" entrytime="00:00:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-11-25" firstname="Egle" gender="F" lastname="Vaupsaite" nation="LTU" athleteid="107869">
              <RESULTS>
                <RESULT eventid="98814" points="284" reactiontime="+96" swimtime="00:03:05.29" resultid="107870" heatid="110616" lane="5" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.77" />
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                    <SPLIT distance="75" swimtime="00:01:06.10" />
                    <SPLIT distance="100" swimtime="00:01:29.18" />
                    <SPLIT distance="125" swimtime="00:01:53.37" />
                    <SPLIT distance="150" swimtime="00:02:17.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="325" swimtime="00:03:15.57" resultid="107871" heatid="110664" lane="9" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.17" />
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="75" swimtime="00:01:07.79" />
                    <SPLIT distance="100" swimtime="00:01:32.69" />
                    <SPLIT distance="125" swimtime="00:01:57.97" />
                    <SPLIT distance="150" swimtime="00:02:23.67" />
                    <SPLIT distance="175" swimtime="00:02:49.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="330" reactiontime="+92" swimtime="00:01:21.95" resultid="107872" heatid="110693" lane="8" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.80" />
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="75" swimtime="00:01:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="333" swimtime="00:01:29.92" resultid="107873" heatid="110724" lane="6" entrytime="00:01:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.66" />
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                    <SPLIT distance="75" swimtime="00:01:04.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="263" reactiontime="+95" swimtime="00:06:44.58" resultid="107874" heatid="110786" lane="5" entrytime="00:06:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.88" />
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                    <SPLIT distance="75" swimtime="00:01:12.19" />
                    <SPLIT distance="100" swimtime="00:01:40.26" />
                    <SPLIT distance="125" swimtime="00:03:02.02" />
                    <SPLIT distance="150" swimtime="00:02:35.11" />
                    <SPLIT distance="175" swimtime="00:03:53.67" />
                    <SPLIT distance="200" swimtime="00:03:28.23" />
                    <SPLIT distance="225" swimtime="00:04:45.54" />
                    <SPLIT distance="250" swimtime="00:04:19.56" />
                    <SPLIT distance="300" swimtime="00:05:11.79" />
                    <SPLIT distance="325" swimtime="00:05:36.35" />
                    <SPLIT distance="350" swimtime="00:06:00.10" />
                    <SPLIT distance="375" swimtime="00:06:23.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-23" firstname="Oksana" gender="F" lastname="Omelcenko" nation="LTU" athleteid="107835">
              <RESULTS>
                <RESULT eventid="98814" points="248" reactiontime="+86" swimtime="00:03:13.86" resultid="107836" heatid="110616" lane="2" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.38" />
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="75" swimtime="00:01:05.91" />
                    <SPLIT distance="100" swimtime="00:01:32.57" />
                    <SPLIT distance="125" swimtime="00:01:59.91" />
                    <SPLIT distance="150" swimtime="00:02:27.53" />
                    <SPLIT distance="175" swimtime="00:02:51.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" status="DNS" swimtime="00:00:00.00" resultid="107837" heatid="110648" lane="4" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="98972" points="266" reactiontime="+94" swimtime="00:01:28.06" resultid="107838" heatid="110692" lane="5" entrytime="00:01:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.23" />
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="75" swimtime="00:01:06.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="268" swimtime="00:00:37.78" resultid="107839" heatid="110738" lane="6" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="262" reactiontime="+58" swimtime="00:06:45.22" resultid="107840" heatid="110786" lane="6" entrytime="00:07:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.98" />
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="75" swimtime="00:01:13.39" />
                    <SPLIT distance="100" swimtime="00:01:41.01" />
                    <SPLIT distance="125" swimtime="00:02:07.82" />
                    <SPLIT distance="150" swimtime="00:02:34.01" />
                    <SPLIT distance="175" swimtime="00:03:01.09" />
                    <SPLIT distance="200" swimtime="00:03:28.75" />
                    <SPLIT distance="225" swimtime="00:03:56.33" />
                    <SPLIT distance="250" swimtime="00:04:23.69" />
                    <SPLIT distance="275" swimtime="00:04:49.98" />
                    <SPLIT distance="300" swimtime="00:05:17.11" />
                    <SPLIT distance="325" swimtime="00:05:41.02" />
                    <SPLIT distance="350" swimtime="00:06:03.84" />
                    <SPLIT distance="375" swimtime="00:06:25.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="215" reactiontime="+76" swimtime="00:03:19.02" resultid="107841" heatid="110808" lane="6" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.49" />
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                    <SPLIT distance="75" swimtime="00:01:09.77" />
                    <SPLIT distance="100" swimtime="00:01:35.50" />
                    <SPLIT distance="125" swimtime="00:02:01.43" />
                    <SPLIT distance="150" swimtime="00:02:28.30" />
                    <SPLIT distance="175" swimtime="00:02:55.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-10-21" firstname="Rasa" gender="F" lastname="Pociuviene" nation="LTU" athleteid="107860">
              <RESULTS>
                <RESULT eventid="106294" points="120" reactiontime="+95" swimtime="00:00:51.94" resultid="107861" heatid="110647" lane="7" entrytime="00:00:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="191" reactiontime="+131" swimtime="00:03:53.27" resultid="107862" heatid="110662" lane="1" entrytime="00:03:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.25" />
                    <SPLIT distance="50" swimtime="00:00:53.54" />
                    <SPLIT distance="75" swimtime="00:01:21.91" />
                    <SPLIT distance="100" swimtime="00:01:51.63" />
                    <SPLIT distance="125" swimtime="00:02:21.15" />
                    <SPLIT distance="150" swimtime="00:02:51.21" />
                    <SPLIT distance="175" swimtime="00:03:22.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="198" reactiontime="+105" swimtime="00:01:46.90" resultid="107863" heatid="110722" lane="7" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.65" />
                    <SPLIT distance="50" swimtime="00:00:50.53" />
                    <SPLIT distance="75" swimtime="00:01:18.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="207" reactiontime="+107" swimtime="00:00:48.63" resultid="107864" heatid="110820" lane="3" entrytime="00:00:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-08" firstname="Dovydas" gender="M" lastname="Eiza" nation="LTU" athleteid="107876">
              <RESULTS>
                <RESULT eventid="98798" points="334" reactiontime="+85" swimtime="00:00:29.19" resultid="107877" heatid="110601" lane="3" entrytime="00:00:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="187" reactiontime="+79" swimtime="00:00:38.79" resultid="107878" heatid="110655" lane="1" entrytime="00:00:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="309" swimtime="00:01:22.22" resultid="107879" heatid="110731" lane="9" entrytime="00:01:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.32" />
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="75" swimtime="00:00:59.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="343" reactiontime="+71" swimtime="00:00:36.06" resultid="107880" heatid="110831" lane="8" entrytime="00:00:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-10-29" firstname="Tomas" gender="M" lastname="Zemaitis" nation="LTU" athleteid="107829">
              <RESULTS>
                <RESULT eventid="98830" points="349" reactiontime="+66" swimtime="00:02:35.68" resultid="107830" heatid="110625" lane="7" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.46" />
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="75" swimtime="00:00:51.69" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="125" swimtime="00:01:35.23" />
                    <SPLIT distance="150" swimtime="00:01:59.17" />
                    <SPLIT distance="175" swimtime="00:02:17.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="321" reactiontime="+71" swimtime="00:00:32.43" resultid="107831" heatid="110657" lane="4" entrytime="00:00:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="368" reactiontime="+72" swimtime="00:01:10.68" resultid="107832" heatid="110702" lane="5" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.37" />
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="75" swimtime="00:00:54.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="365" reactiontime="+85" swimtime="00:00:30.49" resultid="107833" heatid="110747" lane="4" entrytime="00:00:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="323" reactiontime="+82" swimtime="00:01:10.56" resultid="107834" heatid="110802" lane="8" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.90" />
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="75" swimtime="00:00:50.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="420" reactiontime="+84" swimtime="00:01:50.24" resultid="107883" heatid="110781" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:28.17" />
                    <SPLIT distance="75" swimtime="00:00:42.19" />
                    <SPLIT distance="100" swimtime="00:00:57.39" />
                    <SPLIT distance="125" swimtime="00:01:10.38" />
                    <SPLIT distance="150" swimtime="00:01:24.82" />
                    <SPLIT distance="175" swimtime="00:01:36.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107847" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="107865" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="107829" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="107842" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99059" points="376" reactiontime="+89" swimtime="00:02:05.34" resultid="107884" heatid="110716" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.28" />
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="75" swimtime="00:00:48.27" />
                    <SPLIT distance="100" swimtime="00:01:00.18" />
                    <SPLIT distance="125" swimtime="00:01:22.34" />
                    <SPLIT distance="150" swimtime="00:01:40.13" />
                    <SPLIT distance="175" swimtime="00:01:52.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107829" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="107847" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="107865" number="3" />
                    <RELAYPOSITION athleteid="107842" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99234" points="284" reactiontime="+91" swimtime="00:02:23.21" resultid="107881" heatid="110779" lane="4">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.66" />
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="75" swimtime="00:00:50.36" />
                    <SPLIT distance="100" swimtime="00:01:08.13" />
                    <SPLIT distance="125" swimtime="00:01:28.63" />
                    <SPLIT distance="150" swimtime="00:01:50.03" />
                    <SPLIT distance="175" swimtime="00:02:06.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107835" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="107853" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="107860" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="107869" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99036" points="272" reactiontime="+85" swimtime="00:02:40.51" resultid="107882" heatid="110714" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.64" />
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="75" swimtime="00:01:04.19" />
                    <SPLIT distance="100" swimtime="00:01:29.82" />
                    <SPLIT distance="125" swimtime="00:01:46.63" />
                    <SPLIT distance="150" swimtime="00:01:56.16" />
                    <SPLIT distance="175" swimtime="00:02:23.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107835" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="107860" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="107853" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="107869" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="313" reactiontime="+91" swimtime="00:02:01.56" resultid="107885" heatid="110629" lane="2">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.07" />
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="75" swimtime="00:00:45.12" />
                    <SPLIT distance="100" swimtime="00:01:02.51" />
                    <SPLIT distance="125" swimtime="00:01:18.85" />
                    <SPLIT distance="150" swimtime="00:01:36.05" />
                    <SPLIT distance="175" swimtime="00:01:48.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107829" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="107853" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="107869" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="107842" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="286" reactiontime="+78" swimtime="00:02:17.37" resultid="107886" heatid="110835" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.30" />
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="75" swimtime="00:00:51.63" />
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="125" swimtime="00:01:30.95" />
                    <SPLIT distance="150" swimtime="00:01:51.54" />
                    <SPLIT distance="175" swimtime="00:02:03.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107829" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="107869" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="107853" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="107842" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="234" reactiontime="+68" swimtime="00:02:14.01" resultid="107887" heatid="110629" lane="6">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="75" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:00:57.24" />
                    <SPLIT distance="125" swimtime="00:01:14.10" />
                    <SPLIT distance="150" swimtime="00:01:32.66" />
                    <SPLIT distance="175" swimtime="00:01:52.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107835" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="107860" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="107865" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="107847" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="107888" heatid="110835" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107835" number="1" />
                    <RELAYPOSITION athleteid="107860" number="2" />
                    <RELAYPOSITION athleteid="107865" number="3" />
                    <RELAYPOSITION athleteid="107847" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" region="WIE" clubid="107786" name="KS Extreme Team Oborniki">
          <CONTACT city="OBORNIKI" email="janwol@poczta.onet.pl" name="WOLNIEWICZ JANUSZ" phone="791064667" state="WIE" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="107787">
              <RESULTS>
                <RESULT eventid="98798" points="176" reactiontime="+93" swimtime="00:00:36.15" resultid="107788" heatid="110599" lane="1" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="117" reactiontime="+92" swimtime="00:28:53.64" resultid="107789" heatid="110643" lane="8" entrytime="00:29:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.66" />
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                    <SPLIT distance="75" swimtime="00:01:10.04" />
                    <SPLIT distance="100" swimtime="00:01:35.96" />
                    <SPLIT distance="125" swimtime="00:02:02.67" />
                    <SPLIT distance="150" swimtime="00:02:29.68" />
                    <SPLIT distance="175" swimtime="00:02:57.13" />
                    <SPLIT distance="200" swimtime="00:03:25.52" />
                    <SPLIT distance="225" swimtime="00:03:53.25" />
                    <SPLIT distance="250" swimtime="00:04:21.51" />
                    <SPLIT distance="275" swimtime="00:04:49.43" />
                    <SPLIT distance="300" swimtime="00:05:17.72" />
                    <SPLIT distance="325" swimtime="00:05:45.83" />
                    <SPLIT distance="350" swimtime="00:06:14.09" />
                    <SPLIT distance="375" swimtime="00:06:42.90" />
                    <SPLIT distance="400" swimtime="00:07:11.44" />
                    <SPLIT distance="425" swimtime="00:07:40.09" />
                    <SPLIT distance="450" swimtime="00:08:09.03" />
                    <SPLIT distance="475" swimtime="00:08:38.10" />
                    <SPLIT distance="500" swimtime="00:09:07.18" />
                    <SPLIT distance="525" swimtime="00:09:35.69" />
                    <SPLIT distance="550" swimtime="00:10:04.89" />
                    <SPLIT distance="575" swimtime="00:10:33.98" />
                    <SPLIT distance="600" swimtime="00:11:03.54" />
                    <SPLIT distance="625" swimtime="00:11:33.84" />
                    <SPLIT distance="650" swimtime="00:12:03.17" />
                    <SPLIT distance="675" swimtime="00:12:32.70" />
                    <SPLIT distance="700" swimtime="00:13:02.11" />
                    <SPLIT distance="725" swimtime="00:13:33.07" />
                    <SPLIT distance="750" swimtime="00:14:02.60" />
                    <SPLIT distance="775" swimtime="00:14:32.65" />
                    <SPLIT distance="800" swimtime="00:15:01.72" />
                    <SPLIT distance="825" swimtime="00:15:30.96" />
                    <SPLIT distance="850" swimtime="00:16:00.85" />
                    <SPLIT distance="875" swimtime="00:16:30.36" />
                    <SPLIT distance="900" swimtime="00:17:00.51" />
                    <SPLIT distance="925" swimtime="00:17:30.10" />
                    <SPLIT distance="950" swimtime="00:18:00.90" />
                    <SPLIT distance="975" swimtime="00:18:30.43" />
                    <SPLIT distance="1000" swimtime="00:19:01.20" />
                    <SPLIT distance="1025" swimtime="00:19:30.39" />
                    <SPLIT distance="1050" swimtime="00:20:00.01" />
                    <SPLIT distance="1075" swimtime="00:20:28.96" />
                    <SPLIT distance="1100" swimtime="00:20:58.38" />
                    <SPLIT distance="1125" swimtime="00:21:27.40" />
                    <SPLIT distance="1150" swimtime="00:21:57.83" />
                    <SPLIT distance="1175" swimtime="00:22:27.66" />
                    <SPLIT distance="1200" swimtime="00:22:57.70" />
                    <SPLIT distance="1225" swimtime="00:23:28.37" />
                    <SPLIT distance="1250" swimtime="00:23:58.48" />
                    <SPLIT distance="1275" swimtime="00:24:28.37" />
                    <SPLIT distance="1300" swimtime="00:24:58.02" />
                    <SPLIT distance="1325" swimtime="00:25:27.88" />
                    <SPLIT distance="1350" swimtime="00:25:58.27" />
                    <SPLIT distance="1375" swimtime="00:26:28.28" />
                    <SPLIT distance="1400" swimtime="00:26:57.80" />
                    <SPLIT distance="1425" swimtime="00:27:27.73" />
                    <SPLIT distance="1450" swimtime="00:27:56.91" />
                    <SPLIT distance="1475" swimtime="00:28:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="164" reactiontime="+94" swimtime="00:01:22.08" resultid="107790" heatid="110680" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.69" />
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="75" swimtime="00:01:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="107791" heatid="110696" lane="3" entrytime="00:02:00.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="107792" heatid="110742" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="99218" points="126" swimtime="00:03:18.12" resultid="107793" heatid="110771" lane="9" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.03" />
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="75" swimtime="00:01:07.14" />
                    <SPLIT distance="100" swimtime="00:01:32.51" />
                    <SPLIT distance="125" swimtime="00:01:59.09" />
                    <SPLIT distance="150" swimtime="00:02:26.01" />
                    <SPLIT distance="175" swimtime="00:02:52.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="107794" heatid="110798" lane="3" entrytime="00:02:00.00" />
                <RESULT eventid="99473" points="115" swimtime="00:07:15.40" resultid="107795" heatid="110850" lane="9" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.53" />
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                    <SPLIT distance="75" swimtime="00:01:11.87" />
                    <SPLIT distance="100" swimtime="00:01:38.71" />
                    <SPLIT distance="125" swimtime="00:02:06.74" />
                    <SPLIT distance="150" swimtime="00:02:34.68" />
                    <SPLIT distance="175" swimtime="00:03:02.22" />
                    <SPLIT distance="200" swimtime="00:03:30.62" />
                    <SPLIT distance="225" swimtime="00:03:59.15" />
                    <SPLIT distance="250" swimtime="00:04:27.33" />
                    <SPLIT distance="275" swimtime="00:04:55.45" />
                    <SPLIT distance="300" swimtime="00:05:23.83" />
                    <SPLIT distance="325" swimtime="00:05:52.92" />
                    <SPLIT distance="350" swimtime="00:06:22.01" />
                    <SPLIT distance="375" swimtime="00:06:49.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" clubid="108223" name="KS niezrzeszeni.pl">
          <CONTACT name="K.S.niezrzeszeni.pl" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="108224">
              <RESULTS>
                <RESULT eventid="98798" points="188" reactiontime="+114" swimtime="00:00:35.32" resultid="108225" heatid="110594" lane="4">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" reactiontime="+120" status="DNF" swimtime="00:00:00.00" resultid="108226" heatid="110621" lane="1" entrytime="00:03:28.97">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.17" />
                    <SPLIT distance="50" swimtime="00:00:47.82" />
                    <SPLIT distance="75" swimtime="00:01:14.11" />
                    <SPLIT distance="100" swimtime="00:01:39.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 " eventid="98924" status="DSQ" swimtime="00:00:00.00" resultid="108227" heatid="110654" lane="3" entrytime="00:00:40.20" />
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="108228" heatid="110680" lane="6" entrytime="00:01:20.42" />
                <RESULT eventid="99091" points="150" swimtime="00:01:44.46" resultid="108229" heatid="110727" lane="0">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.77" />
                    <SPLIT distance="50" swimtime="00:00:50.84" />
                    <SPLIT distance="75" swimtime="00:01:18.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="171" reactiontime="+69" swimtime="00:01:27.97" resultid="108230" heatid="110759" lane="6" entrytime="00:01:28.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.37" />
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                    <SPLIT distance="75" swimtime="00:01:06.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="181" reactiontime="+72" swimtime="00:03:06.64" resultid="108231" heatid="110812" lane="5" entrytime="00:03:09.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.39" />
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                    <SPLIT distance="75" swimtime="00:01:07.19" />
                    <SPLIT distance="100" swimtime="00:01:30.88" />
                    <SPLIT distance="125" swimtime="00:01:55.04" />
                    <SPLIT distance="150" swimtime="00:02:19.08" />
                    <SPLIT distance="175" swimtime="00:02:43.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-08-04" firstname="Wojciech" gender="M" lastname="Staruch" nation="POL" athleteid="108232">
              <RESULTS>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="108233" heatid="110620" lane="6" entrytime="00:03:43.20" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="108234" heatid="110666" lane="3" entrytime="00:03:43.00" />
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="108235" heatid="110710" lane="3" entrytime="00:04:00.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="108236" heatid="110729" lane="9" entrytime="00:01:42.30" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="108237" heatid="110799" lane="7" entrytime="00:01:43.30" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="108238" heatid="110826" lane="8" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="DOL" clubid="107364" name="KS Rekin Świebodzice">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztof" phone="606626274" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1984-04-16" firstname="Filip" gender="M" lastname="Żemier" nation="POL" athleteid="107405">
              <RESULTS>
                <RESULT eventid="98798" points="496" reactiontime="+70" swimtime="00:00:25.58" resultid="107406" heatid="110610" lane="5" entrytime="00:00:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="467" swimtime="00:00:57.91" resultid="107407" heatid="110686" lane="9" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.05" />
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="75" swimtime="00:00:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="374" reactiontime="+81" swimtime="00:01:10.31" resultid="107408" heatid="110704" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="75" swimtime="00:00:53.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="386" reactiontime="+75" swimtime="00:00:29.92" resultid="107409" heatid="110748" lane="1" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="375" reactiontime="+81" swimtime="00:02:17.79" resultid="107410" heatid="110769" lane="8">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="75" swimtime="00:00:52.06" />
                    <SPLIT distance="100" swimtime="00:01:09.91" />
                    <SPLIT distance="125" swimtime="00:01:28.09" />
                    <SPLIT distance="150" swimtime="00:01:46.52" />
                    <SPLIT distance="175" swimtime="00:02:02.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="302" reactiontime="+85" swimtime="00:01:12.19" resultid="107411" heatid="110797" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.32" />
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="75" swimtime="00:00:51.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="339" reactiontime="+66" swimtime="00:00:36.19" resultid="107412" heatid="110830" lane="8" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-18" firstname="Marek" gender="M" lastname="Stuczyński" nation="POL" athleteid="107390">
              <RESULTS>
                <RESULT eventid="98798" points="535" reactiontime="+81" swimtime="00:00:24.95" resultid="107391" heatid="110612" lane="1" entrytime="00:00:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="533" swimtime="00:00:55.41" resultid="107392" heatid="110689" lane="9" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.63" />
                    <SPLIT distance="50" swimtime="00:00:26.46" />
                    <SPLIT distance="75" swimtime="00:00:40.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="473" reactiontime="+76" swimtime="00:01:04.98" resultid="107393" heatid="110706" lane="8" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.11" />
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                    <SPLIT distance="75" swimtime="00:00:48.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="547" reactiontime="+82" swimtime="00:01:07.97" resultid="107394" heatid="110734" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.23" />
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="75" swimtime="00:00:49.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="553" reactiontime="+73" swimtime="00:00:30.75" resultid="107395" heatid="110834" lane="7" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="107377">
              <RESULTS>
                <RESULT eventid="98777" points="342" reactiontime="+100" swimtime="00:00:33.22" resultid="107378" heatid="110590" lane="3" entrytime="00:00:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="230" reactiontime="+100" swimtime="00:03:39.46" resultid="107379" heatid="110662" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.48" />
                    <SPLIT distance="50" swimtime="00:00:49.23" />
                    <SPLIT distance="75" swimtime="00:01:16.70" />
                    <SPLIT distance="100" swimtime="00:01:45.27" />
                    <SPLIT distance="125" swimtime="00:02:13.82" />
                    <SPLIT distance="150" swimtime="00:02:43.01" />
                    <SPLIT distance="175" swimtime="00:03:11.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="311" reactiontime="+94" swimtime="00:01:15.11" resultid="107380" heatid="110674" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.91" />
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="75" swimtime="00:00:55.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="228" reactiontime="+95" swimtime="00:01:41.98" resultid="107381" heatid="110724" lane="8" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.82" />
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                    <SPLIT distance="75" swimtime="00:01:14.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="281" reactiontime="+102" swimtime="00:02:49.00" resultid="107382" heatid="110766" lane="8" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.92" />
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="75" swimtime="00:00:59.99" />
                    <SPLIT distance="100" swimtime="00:01:21.89" />
                    <SPLIT distance="125" swimtime="00:01:44.59" />
                    <SPLIT distance="150" swimtime="00:02:07.13" />
                    <SPLIT distance="175" swimtime="00:02:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="226" reactiontime="+109" swimtime="00:03:15.62" resultid="107383" heatid="110808" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.99" />
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                    <SPLIT distance="75" swimtime="00:01:11.72" />
                    <SPLIT distance="100" swimtime="00:01:36.49" />
                    <SPLIT distance="125" swimtime="00:02:01.60" />
                    <SPLIT distance="150" swimtime="00:02:27.08" />
                    <SPLIT distance="175" swimtime="00:02:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="235" swimtime="00:00:46.66" resultid="107384" heatid="110820" lane="0" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-07-17" firstname="Agnieszka" gender="F" lastname="Gajdowska" nation="POL" license="S02001100002" athleteid="107368">
              <RESULTS>
                <RESULT eventid="98777" points="641" reactiontime="+64" swimtime="00:00:26.94" resultid="107369" heatid="110593" lane="5" entrytime="00:00:26.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="479" reactiontime="+64" swimtime="00:02:35.67" resultid="107370" heatid="110618" lane="5" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.73" />
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="75" swimtime="00:00:51.43" />
                    <SPLIT distance="100" swimtime="00:01:11.18" />
                    <SPLIT distance="125" swimtime="00:01:34.72" />
                    <SPLIT distance="150" swimtime="00:01:59.10" />
                    <SPLIT distance="175" swimtime="00:02:18.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="464" reactiontime="+91" swimtime="00:00:33.14" resultid="107371" heatid="110650" lane="2" entrytime="00:00:32.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="628" reactiontime="+65" swimtime="00:00:59.44" resultid="107372" heatid="110676" lane="5" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="75" swimtime="00:00:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="521" reactiontime="+66" swimtime="00:00:30.29" resultid="107373" heatid="110740" lane="4" entrytime="00:00:29.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="557" reactiontime="+69" swimtime="00:02:14.64" resultid="107374" heatid="110768" lane="5" entrytime="00:02:14.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.65" />
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="75" swimtime="00:00:45.82" />
                    <SPLIT distance="100" swimtime="00:01:02.80" />
                    <SPLIT distance="125" swimtime="00:01:20.46" />
                    <SPLIT distance="150" swimtime="00:01:38.79" />
                    <SPLIT distance="175" swimtime="00:01:57.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="459" swimtime="00:00:37.31" resultid="107375" heatid="110823" lane="9" entrytime="00:00:37.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="527" reactiontime="+69" swimtime="00:04:50.25" resultid="107376" heatid="110839" lane="4" entrytime="00:04:45.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.13" />
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="75" swimtime="00:00:49.44" />
                    <SPLIT distance="100" swimtime="00:01:08.01" />
                    <SPLIT distance="125" swimtime="00:01:27.03" />
                    <SPLIT distance="150" swimtime="00:01:46.29" />
                    <SPLIT distance="175" swimtime="00:02:05.41" />
                    <SPLIT distance="200" swimtime="00:02:24.24" />
                    <SPLIT distance="225" swimtime="00:02:43.16" />
                    <SPLIT distance="250" swimtime="00:03:02.00" />
                    <SPLIT distance="275" swimtime="00:03:20.86" />
                    <SPLIT distance="300" swimtime="00:03:39.65" />
                    <SPLIT distance="325" swimtime="00:03:58.61" />
                    <SPLIT distance="350" swimtime="00:04:16.93" />
                    <SPLIT distance="375" swimtime="00:04:34.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-11-09" firstname="Karol" gender="M" lastname="Żemier" nation="POL" athleteid="107413">
              <RESULTS>
                <RESULT eventid="98798" points="529" reactiontime="+70" swimtime="00:00:25.04" resultid="107414" heatid="110612" lane="8" entrytime="00:00:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="555" reactiontime="+72" swimtime="00:02:13.34" resultid="107415" heatid="110628" lane="7" entrytime="00:02:19.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.45" />
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                    <SPLIT distance="75" swimtime="00:00:44.94" />
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                    <SPLIT distance="125" swimtime="00:01:21.29" />
                    <SPLIT distance="150" swimtime="00:01:41.42" />
                    <SPLIT distance="175" swimtime="00:01:58.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="542" reactiontime="+60" swimtime="00:00:27.25" resultid="107416" heatid="110660" lane="6" entrytime="00:00:27.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="594" reactiontime="+71" swimtime="00:01:00.26" resultid="107417" heatid="110706" lane="6" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                    <SPLIT distance="75" swimtime="00:00:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="525" reactiontime="+60" swimtime="00:00:27.01" resultid="107418" heatid="110741" lane="4">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="557" reactiontime="+68" swimtime="00:00:59.44" resultid="107419" heatid="110763" lane="3" entrytime="00:01:00.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                    <SPLIT distance="75" swimtime="00:00:44.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="566" reactiontime="+78" swimtime="00:00:58.54" resultid="107420" heatid="110797" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.31" />
                    <SPLIT distance="50" swimtime="00:00:27.13" />
                    <SPLIT distance="75" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="545" reactiontime="+65" swimtime="00:02:09.31" resultid="107421" heatid="110816" lane="3" entrytime="00:02:14.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.18" />
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="75" swimtime="00:00:45.75" />
                    <SPLIT distance="100" swimtime="00:01:02.35" />
                    <SPLIT distance="125" swimtime="00:01:18.86" />
                    <SPLIT distance="150" swimtime="00:01:35.82" />
                    <SPLIT distance="175" swimtime="00:01:52.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-12-12" firstname="Karolina" gender="F" lastname="Jahnz" nation="POL" athleteid="107385">
              <RESULTS>
                <RESULT eventid="98863" points="290" reactiontime="+56" swimtime="00:12:03.75" resultid="107386" heatid="110634" lane="4" entrytime="00:12:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.71" />
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="75" swimtime="00:00:59.13" />
                    <SPLIT distance="100" swimtime="00:01:21.37" />
                    <SPLIT distance="125" swimtime="00:01:44.02" />
                    <SPLIT distance="150" swimtime="00:02:06.75" />
                    <SPLIT distance="175" swimtime="00:02:29.77" />
                    <SPLIT distance="200" swimtime="00:02:52.35" />
                    <SPLIT distance="225" swimtime="00:03:15.28" />
                    <SPLIT distance="250" swimtime="00:03:38.37" />
                    <SPLIT distance="275" swimtime="00:04:01.42" />
                    <SPLIT distance="300" swimtime="00:04:24.38" />
                    <SPLIT distance="325" swimtime="00:04:47.45" />
                    <SPLIT distance="350" swimtime="00:05:10.55" />
                    <SPLIT distance="375" swimtime="00:05:33.92" />
                    <SPLIT distance="400" swimtime="00:05:57.51" />
                    <SPLIT distance="425" swimtime="00:06:20.79" />
                    <SPLIT distance="450" swimtime="00:06:44.03" />
                    <SPLIT distance="475" swimtime="00:07:07.40" />
                    <SPLIT distance="500" swimtime="00:07:30.44" />
                    <SPLIT distance="525" swimtime="00:07:53.47" />
                    <SPLIT distance="550" swimtime="00:08:16.87" />
                    <SPLIT distance="575" swimtime="00:08:40.01" />
                    <SPLIT distance="600" swimtime="00:09:03.10" />
                    <SPLIT distance="625" swimtime="00:09:26.24" />
                    <SPLIT distance="650" swimtime="00:09:48.86" />
                    <SPLIT distance="675" swimtime="00:10:11.73" />
                    <SPLIT distance="700" swimtime="00:10:34.80" />
                    <SPLIT distance="725" swimtime="00:10:57.72" />
                    <SPLIT distance="750" swimtime="00:11:20.34" />
                    <SPLIT distance="775" swimtime="00:11:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="274" swimtime="00:03:26.94" resultid="107387" heatid="110663" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.54" />
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                    <SPLIT distance="75" swimtime="00:01:13.12" />
                    <SPLIT distance="100" swimtime="00:01:39.89" />
                    <SPLIT distance="125" swimtime="00:02:06.92" />
                    <SPLIT distance="150" swimtime="00:02:33.93" />
                    <SPLIT distance="175" swimtime="00:03:00.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="281" reactiontime="+82" swimtime="00:06:35.71" resultid="107388" heatid="110785" lane="6">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.05" />
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                    <SPLIT distance="75" swimtime="00:01:10.13" />
                    <SPLIT distance="100" swimtime="00:01:36.70" />
                    <SPLIT distance="125" swimtime="00:02:01.62" />
                    <SPLIT distance="150" swimtime="00:02:25.77" />
                    <SPLIT distance="175" swimtime="00:02:50.40" />
                    <SPLIT distance="200" swimtime="00:03:15.00" />
                    <SPLIT distance="225" swimtime="00:03:42.97" />
                    <SPLIT distance="250" swimtime="00:04:10.15" />
                    <SPLIT distance="275" swimtime="00:04:37.89" />
                    <SPLIT distance="300" swimtime="00:05:05.89" />
                    <SPLIT distance="325" swimtime="00:05:29.67" />
                    <SPLIT distance="350" swimtime="00:05:52.36" />
                    <SPLIT distance="375" swimtime="00:06:14.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="305" reactiontime="+65" swimtime="00:05:48.29" resultid="107389" heatid="110841" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.88" />
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="75" swimtime="00:00:59.29" />
                    <SPLIT distance="100" swimtime="00:01:20.94" />
                    <SPLIT distance="125" swimtime="00:01:43.23" />
                    <SPLIT distance="150" swimtime="00:02:05.41" />
                    <SPLIT distance="175" swimtime="00:02:27.94" />
                    <SPLIT distance="200" swimtime="00:02:50.19" />
                    <SPLIT distance="225" swimtime="00:03:12.37" />
                    <SPLIT distance="250" swimtime="00:03:34.72" />
                    <SPLIT distance="275" swimtime="00:03:57.04" />
                    <SPLIT distance="300" swimtime="00:04:19.80" />
                    <SPLIT distance="325" swimtime="00:04:42.05" />
                    <SPLIT distance="350" swimtime="00:05:04.44" />
                    <SPLIT distance="375" swimtime="00:05:26.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-21" firstname="Alfred" gender="M" lastname="Żemier" nation="POL" athleteid="107396">
              <RESULTS>
                <RESULT eventid="98798" points="529" reactiontime="+69" swimtime="00:00:25.04" resultid="107397" heatid="110611" lane="4" entrytime="00:00:25.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="366" reactiontime="+85" swimtime="00:02:33.24" resultid="107398" heatid="110619" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.20" />
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="75" swimtime="00:00:49.76" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="125" swimtime="00:01:33.04" />
                    <SPLIT distance="150" swimtime="00:01:56.12" />
                    <SPLIT distance="175" swimtime="00:02:15.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="402" reactiontime="+67" swimtime="00:00:30.09" resultid="107399" heatid="110659" lane="4" entrytime="00:00:29.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="507" reactiontime="+83" swimtime="00:00:56.33" resultid="107400" heatid="110688" lane="4" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.76" />
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                    <SPLIT distance="75" swimtime="00:00:41.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="493" reactiontime="+77" swimtime="00:00:27.59" resultid="107401" heatid="110741" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="397" reactiontime="+72" swimtime="00:01:06.55" resultid="107402" heatid="110763" lane="9" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.12" />
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="75" swimtime="00:00:50.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="450" swimtime="00:01:03.17" resultid="107403" heatid="110798" lane="9">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.04" />
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                    <SPLIT distance="75" swimtime="00:00:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="410" reactiontime="+62" swimtime="00:00:33.98" resultid="107404" heatid="110832" lane="5" entrytime="00:00:34.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="REKIN ŚWIEBODZICE B" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="553" reactiontime="+64" swimtime="00:01:50.22" resultid="107424" heatid="110719" lane="3" entrytime="00:01:50.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="75" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:00:57.83" />
                    <SPLIT distance="125" swimtime="00:01:10.37" />
                    <SPLIT distance="150" swimtime="00:01:25.23" />
                    <SPLIT distance="175" swimtime="00:01:37.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107413" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="107390" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="107396" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="107405" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="581" reactiontime="+79" swimtime="00:01:38.95" resultid="107425" heatid="110784" lane="3" entrytime="00:01:39.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                    <SPLIT distance="50" swimtime="00:00:25.07" />
                    <SPLIT distance="75" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:00:49.52" />
                    <SPLIT distance="125" swimtime="00:01:01.03" />
                    <SPLIT distance="150" swimtime="00:01:14.14" />
                    <SPLIT distance="175" swimtime="00:01:25.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107413" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="107390" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="107396" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="107405" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="REKIN ŚWIEBODZICE B" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="346" reactiontime="+87" swimtime="00:01:57.58" resultid="107422" heatid="110632" lane="0" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.01" />
                    <SPLIT distance="50" swimtime="00:00:24.96" />
                    <SPLIT distance="75" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:00:59.22" />
                    <SPLIT distance="125" swimtime="00:01:14.89" />
                    <SPLIT distance="150" swimtime="00:01:31.84" />
                    <SPLIT distance="175" swimtime="00:01:43.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107396" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="107385" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="107377" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="107405" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="348" reactiontime="+69" swimtime="00:02:08.61" resultid="107423" heatid="110838" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.21" />
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                    <SPLIT distance="75" swimtime="00:00:52.69" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="125" swimtime="00:01:21.31" />
                    <SPLIT distance="150" swimtime="00:01:36.22" />
                    <SPLIT distance="175" swimtime="00:01:52.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107385" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="107390" number="2" />
                    <RELAYPOSITION athleteid="107396" number="3" />
                    <RELAYPOSITION athleteid="107377" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KS WAR" nation="POL" clubid="109484" name="KS Warta Poznań">
          <CONTACT city="POZNAŃ" email="jacek.thiem@gmail.com" name="THIEM JACEK" phone="502 499 565" state="WIE" street="OS. DĘBINA 19 M 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="100115700345" athleteid="109500">
              <RESULTS>
                <RESULT eventid="98891" points="208" reactiontime="+99" swimtime="00:12:27.99" resultid="109501" heatid="110637" lane="8" entrytime="00:12:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.64" />
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="75" swimtime="00:01:03.91" />
                    <SPLIT distance="100" swimtime="00:01:27.59" />
                    <SPLIT distance="125" swimtime="00:01:50.66" />
                    <SPLIT distance="150" swimtime="00:02:14.25" />
                    <SPLIT distance="175" swimtime="00:02:37.91" />
                    <SPLIT distance="200" swimtime="00:03:01.42" />
                    <SPLIT distance="225" swimtime="00:03:25.63" />
                    <SPLIT distance="250" swimtime="00:03:49.53" />
                    <SPLIT distance="275" swimtime="00:04:13.73" />
                    <SPLIT distance="300" swimtime="00:04:37.49" />
                    <SPLIT distance="325" swimtime="00:05:02.00" />
                    <SPLIT distance="350" swimtime="00:05:25.71" />
                    <SPLIT distance="375" swimtime="00:05:49.86" />
                    <SPLIT distance="400" swimtime="00:06:14.30" />
                    <SPLIT distance="425" swimtime="00:06:38.78" />
                    <SPLIT distance="450" swimtime="00:07:02.57" />
                    <SPLIT distance="475" swimtime="00:07:26.90" />
                    <SPLIT distance="500" swimtime="00:07:50.46" />
                    <SPLIT distance="525" swimtime="00:08:14.37" />
                    <SPLIT distance="550" swimtime="00:08:38.20" />
                    <SPLIT distance="575" swimtime="00:09:02.04" />
                    <SPLIT distance="600" swimtime="00:09:25.75" />
                    <SPLIT distance="625" swimtime="00:09:49.53" />
                    <SPLIT distance="650" swimtime="00:10:12.63" />
                    <SPLIT distance="675" swimtime="00:10:36.01" />
                    <SPLIT distance="700" swimtime="00:10:58.70" />
                    <SPLIT distance="725" swimtime="00:11:22.55" />
                    <SPLIT distance="750" swimtime="00:11:45.09" />
                    <SPLIT distance="775" swimtime="00:12:07.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="180" reactiontime="+110" swimtime="00:03:11.94" resultid="109502" heatid="110711" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.82" />
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                    <SPLIT distance="75" swimtime="00:01:09.76" />
                    <SPLIT distance="100" swimtime="00:01:34.55" />
                    <SPLIT distance="125" swimtime="00:01:59.12" />
                    <SPLIT distance="150" swimtime="00:02:23.28" />
                    <SPLIT distance="175" swimtime="00:02:47.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="188" reactiontime="+116" swimtime="00:00:37.99" resultid="109503" heatid="110743" lane="3" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="135" reactiontime="+92" swimtime="00:03:25.68" resultid="109504" heatid="110812" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.70" />
                    <SPLIT distance="50" swimtime="00:00:50.77" />
                    <SPLIT distance="75" swimtime="00:01:16.80" />
                    <SPLIT distance="100" swimtime="00:01:42.69" />
                    <SPLIT distance="125" swimtime="00:02:08.86" />
                    <SPLIT distance="150" swimtime="00:02:35.83" />
                    <SPLIT distance="175" swimtime="00:03:01.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-23" firstname="Przemysław" gender="M" lastname="Kuca" nation="POL" license="100115700396" athleteid="109533">
              <RESULTS>
                <RESULT eventid="98798" points="527" reactiontime="+64" swimtime="00:00:25.08" resultid="109534" heatid="110613" lane="6" entrytime="00:00:23.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="538" reactiontime="+70" swimtime="00:02:14.72" resultid="109535" heatid="110628" lane="4" entrytime="00:02:10.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.71" />
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="75" swimtime="00:00:46.98" />
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                    <SPLIT distance="125" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:01:45.33" />
                    <SPLIT distance="175" swimtime="00:02:00.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="574" reactiontime="+72" swimtime="00:00:54.07" resultid="109536" heatid="110689" lane="5" entrytime="00:00:52.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.19" />
                    <SPLIT distance="50" swimtime="00:00:25.79" />
                    <SPLIT distance="75" swimtime="00:00:39.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="571" reactiontime="+72" swimtime="00:02:10.83" resultid="109537" heatid="110713" lane="5" entrytime="00:02:05.06">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.06" />
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                    <SPLIT distance="75" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:01.69" />
                    <SPLIT distance="125" swimtime="00:01:18.55" />
                    <SPLIT distance="150" swimtime="00:01:35.84" />
                    <SPLIT distance="175" swimtime="00:01:52.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="578" reactiontime="+77" swimtime="00:01:59.24" resultid="109538" heatid="110778" lane="3" entrytime="00:01:56.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.76" />
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                    <SPLIT distance="75" swimtime="00:00:42.64" />
                    <SPLIT distance="100" swimtime="00:00:58.18" />
                    <SPLIT distance="125" swimtime="00:01:13.71" />
                    <SPLIT distance="150" swimtime="00:01:29.53" />
                    <SPLIT distance="175" swimtime="00:01:44.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="556" reactiontime="+73" swimtime="00:04:46.27" resultid="109539" heatid="110792" lane="4" entrytime="00:04:40.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.04" />
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                    <SPLIT distance="75" swimtime="00:00:45.73" />
                    <SPLIT distance="100" swimtime="00:01:03.08" />
                    <SPLIT distance="125" swimtime="00:01:23.11" />
                    <SPLIT distance="150" swimtime="00:01:41.91" />
                    <SPLIT distance="175" swimtime="00:02:00.98" />
                    <SPLIT distance="200" swimtime="00:02:19.90" />
                    <SPLIT distance="225" swimtime="00:02:40.35" />
                    <SPLIT distance="250" swimtime="00:03:01.13" />
                    <SPLIT distance="275" swimtime="00:03:22.20" />
                    <SPLIT distance="300" swimtime="00:03:43.57" />
                    <SPLIT distance="325" swimtime="00:03:59.81" />
                    <SPLIT distance="350" swimtime="00:04:15.55" />
                    <SPLIT distance="375" swimtime="00:04:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="525" swimtime="00:01:00.03" resultid="109540" heatid="110805" lane="2" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="75" swimtime="00:00:43.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="552" reactiontime="+74" swimtime="00:04:18.60" resultid="109541" heatid="110843" lane="4" entrytime="00:04:12.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="75" swimtime="00:00:45.53" />
                    <SPLIT distance="100" swimtime="00:01:01.94" />
                    <SPLIT distance="125" swimtime="00:01:18.40" />
                    <SPLIT distance="150" swimtime="00:01:35.09" />
                    <SPLIT distance="175" swimtime="00:01:51.70" />
                    <SPLIT distance="200" swimtime="00:02:08.52" />
                    <SPLIT distance="225" swimtime="00:02:24.88" />
                    <SPLIT distance="250" swimtime="00:02:41.37" />
                    <SPLIT distance="275" swimtime="00:02:57.81" />
                    <SPLIT distance="300" swimtime="00:03:14.44" />
                    <SPLIT distance="325" swimtime="00:03:31.11" />
                    <SPLIT distance="350" swimtime="00:03:47.83" />
                    <SPLIT distance="375" swimtime="00:04:04.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-22" firstname="Piotr" gender="M" lastname="Kodur" nation="POL" athleteid="109572">
              <RESULTS>
                <RESULT eventid="98830" points="476" reactiontime="+81" swimtime="00:02:20.40" resultid="109573" heatid="110623" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.69" />
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="75" swimtime="00:00:47.11" />
                    <SPLIT distance="100" swimtime="00:01:04.81" />
                    <SPLIT distance="125" swimtime="00:01:25.33" />
                    <SPLIT distance="150" swimtime="00:01:47.11" />
                    <SPLIT distance="175" swimtime="00:02:03.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="420" reactiontime="+63" swimtime="00:00:29.67" resultid="109574" heatid="110656" lane="8" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="109575" heatid="110701" lane="1" entrytime="00:01:15.00" />
                <RESULT eventid="99186" points="457" reactiontime="+73" swimtime="00:01:03.48" resultid="109576" heatid="110761" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.24" />
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                    <SPLIT distance="75" swimtime="00:00:47.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="418" swimtime="00:05:14.73" resultid="109577" heatid="110790" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="75" swimtime="00:00:48.59" />
                    <SPLIT distance="100" swimtime="00:01:07.20" />
                    <SPLIT distance="125" swimtime="00:01:28.47" />
                    <SPLIT distance="150" swimtime="00:01:48.85" />
                    <SPLIT distance="175" swimtime="00:02:09.15" />
                    <SPLIT distance="200" swimtime="00:02:28.64" />
                    <SPLIT distance="225" swimtime="00:02:52.17" />
                    <SPLIT distance="250" swimtime="00:03:15.72" />
                    <SPLIT distance="275" swimtime="00:03:39.31" />
                    <SPLIT distance="300" swimtime="00:04:02.55" />
                    <SPLIT distance="325" swimtime="00:04:22.03" />
                    <SPLIT distance="350" swimtime="00:04:40.20" />
                    <SPLIT distance="375" swimtime="00:04:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="467" swimtime="00:01:02.40" resultid="109578" heatid="110802" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                    <SPLIT distance="75" swimtime="00:00:45.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="412" reactiontime="+71" swimtime="00:02:21.90" resultid="109579" heatid="110813" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.23" />
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="75" swimtime="00:00:52.55" />
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="125" swimtime="00:01:29.03" />
                    <SPLIT distance="150" swimtime="00:01:47.00" />
                    <SPLIT distance="175" swimtime="00:02:04.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" license="100115700344" athleteid="109566">
              <RESULTS>
                <RESULT eventid="98830" points="252" reactiontime="+82" swimtime="00:02:53.56" resultid="109567" heatid="110623" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.86" />
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="75" swimtime="00:01:00.49" />
                    <SPLIT distance="100" swimtime="00:01:24.47" />
                    <SPLIT distance="125" swimtime="00:01:48.79" />
                    <SPLIT distance="150" swimtime="00:02:13.63" />
                    <SPLIT distance="175" swimtime="00:02:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="292" reactiontime="+92" swimtime="00:03:01.55" resultid="109568" heatid="110668" lane="4" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.78" />
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="75" swimtime="00:01:02.14" />
                    <SPLIT distance="100" swimtime="00:01:24.98" />
                    <SPLIT distance="125" swimtime="00:01:48.00" />
                    <SPLIT distance="150" swimtime="00:02:12.00" />
                    <SPLIT distance="175" swimtime="00:02:36.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="253" reactiontime="+96" swimtime="00:01:20.09" resultid="109569" heatid="110699" lane="3" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.33" />
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                    <SPLIT distance="75" swimtime="00:01:00.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="295" reactiontime="+89" swimtime="00:01:23.50" resultid="109570" heatid="110731" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.70" />
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="75" swimtime="00:01:01.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="306" reactiontime="+100" swimtime="00:00:37.43" resultid="109571" heatid="110828" lane="3" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" license="100115700345" athleteid="109505">
              <RESULTS>
                <RESULT eventid="98863" points="239" swimtime="00:12:52.17" resultid="109506" heatid="110634" lane="5" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.15" />
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="75" swimtime="00:01:04.60" />
                    <SPLIT distance="100" swimtime="00:01:26.91" />
                    <SPLIT distance="125" swimtime="00:01:49.65" />
                    <SPLIT distance="150" swimtime="00:02:13.32" />
                    <SPLIT distance="175" swimtime="00:02:36.85" />
                    <SPLIT distance="200" swimtime="00:03:01.35" />
                    <SPLIT distance="225" swimtime="00:03:25.37" />
                    <SPLIT distance="250" swimtime="00:03:49.80" />
                    <SPLIT distance="275" swimtime="00:04:13.57" />
                    <SPLIT distance="300" swimtime="00:04:38.39" />
                    <SPLIT distance="325" swimtime="00:05:03.10" />
                    <SPLIT distance="350" swimtime="00:05:27.73" />
                    <SPLIT distance="375" swimtime="00:05:51.94" />
                    <SPLIT distance="400" swimtime="00:06:16.71" />
                    <SPLIT distance="425" swimtime="00:06:41.37" />
                    <SPLIT distance="450" swimtime="00:07:05.78" />
                    <SPLIT distance="475" swimtime="00:07:30.32" />
                    <SPLIT distance="500" swimtime="00:07:55.14" />
                    <SPLIT distance="525" swimtime="00:08:19.37" />
                    <SPLIT distance="550" swimtime="00:08:44.15" />
                    <SPLIT distance="575" swimtime="00:09:08.88" />
                    <SPLIT distance="600" swimtime="00:09:34.46" />
                    <SPLIT distance="625" swimtime="00:09:59.28" />
                    <SPLIT distance="650" swimtime="00:10:24.28" />
                    <SPLIT distance="675" swimtime="00:10:48.94" />
                    <SPLIT distance="700" swimtime="00:11:13.91" />
                    <SPLIT distance="725" swimtime="00:11:38.70" />
                    <SPLIT distance="750" swimtime="00:12:04.52" />
                    <SPLIT distance="775" swimtime="00:12:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="168" reactiontime="+128" swimtime="00:00:46.50" resultid="109507" heatid="110647" lane="5" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="221" swimtime="00:01:24.10" resultid="109508" heatid="110673" lane="0" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.65" />
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="75" swimtime="00:01:03.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="109509" heatid="110754" lane="3" entrytime="00:01:40.00" />
                <RESULT eventid="99202" points="240" swimtime="00:02:58.13" resultid="109510" heatid="110765" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.10" />
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                    <SPLIT distance="75" swimtime="00:01:04.28" />
                    <SPLIT distance="100" swimtime="00:01:26.72" />
                    <SPLIT distance="125" swimtime="00:01:49.57" />
                    <SPLIT distance="150" swimtime="00:02:12.92" />
                    <SPLIT distance="175" swimtime="00:02:35.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="245" swimtime="00:06:14.37" resultid="109511" heatid="110841" lane="8" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.45" />
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                    <SPLIT distance="75" swimtime="00:01:05.38" />
                    <SPLIT distance="100" swimtime="00:01:28.06" />
                    <SPLIT distance="125" swimtime="00:01:50.71" />
                    <SPLIT distance="150" swimtime="00:02:13.95" />
                    <SPLIT distance="175" swimtime="00:02:37.69" />
                    <SPLIT distance="200" swimtime="00:03:01.27" />
                    <SPLIT distance="225" swimtime="00:03:25.20" />
                    <SPLIT distance="250" swimtime="00:03:49.28" />
                    <SPLIT distance="275" swimtime="00:04:13.92" />
                    <SPLIT distance="300" swimtime="00:04:38.30" />
                    <SPLIT distance="325" swimtime="00:05:02.49" />
                    <SPLIT distance="350" swimtime="00:05:26.75" />
                    <SPLIT distance="375" swimtime="00:05:50.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-22" firstname="Małgorzata" gender="F" lastname="Putowska" nation="POL" athleteid="109542">
              <RESULTS>
                <RESULT eventid="98777" points="176" reactiontime="+93" swimtime="00:00:41.40" resultid="109543" heatid="110587" lane="1" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="146" reactiontime="+88" swimtime="00:03:51.27" resultid="109544" heatid="110614" lane="5" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.17" />
                    <SPLIT distance="50" swimtime="00:00:53.95" />
                    <SPLIT distance="75" swimtime="00:02:26.21" />
                    <SPLIT distance="100" swimtime="00:01:53.02" />
                    <SPLIT distance="150" swimtime="00:02:58.96" />
                    <SPLIT distance="175" swimtime="00:03:26.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="167" swimtime="00:04:04.04" resultid="109545" heatid="110661" lane="4" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.64" />
                    <SPLIT distance="50" swimtime="00:00:54.79" />
                    <SPLIT distance="75" swimtime="00:01:26.51" />
                    <SPLIT distance="100" swimtime="00:01:58.90" />
                    <SPLIT distance="125" swimtime="00:02:32.35" />
                    <SPLIT distance="150" swimtime="00:03:04.66" />
                    <SPLIT distance="175" swimtime="00:03:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="88" reactiontime="+80" swimtime="00:04:28.46" resultid="109546" heatid="110707" lane="5" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.86" />
                    <SPLIT distance="50" swimtime="00:00:54.54" />
                    <SPLIT distance="75" swimtime="00:01:28.88" />
                    <SPLIT distance="100" swimtime="00:02:04.68" />
                    <SPLIT distance="125" swimtime="00:02:41.17" />
                    <SPLIT distance="150" swimtime="00:03:17.88" />
                    <SPLIT distance="175" swimtime="00:03:54.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="120" reactiontime="+77" swimtime="00:01:51.31" resultid="109547" heatid="110754" lane="6" entrytime="00:01:47.73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.30" />
                    <SPLIT distance="50" swimtime="00:00:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="134" swimtime="00:08:26.36" resultid="109548" heatid="110785" lane="4" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.16" />
                    <SPLIT distance="50" swimtime="00:00:55.30" />
                    <SPLIT distance="75" swimtime="00:01:29.31" />
                    <SPLIT distance="100" swimtime="00:02:07.30" />
                    <SPLIT distance="125" swimtime="00:02:38.23" />
                    <SPLIT distance="150" swimtime="00:03:09.99" />
                    <SPLIT distance="175" swimtime="00:03:41.46" />
                    <SPLIT distance="200" swimtime="00:04:12.36" />
                    <SPLIT distance="225" swimtime="00:04:46.81" />
                    <SPLIT distance="250" swimtime="00:05:22.16" />
                    <SPLIT distance="275" swimtime="00:05:57.45" />
                    <SPLIT distance="300" swimtime="00:06:32.06" />
                    <SPLIT distance="325" swimtime="00:07:00.68" />
                    <SPLIT distance="350" swimtime="00:07:29.44" />
                    <SPLIT distance="375" swimtime="00:07:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="77" swimtime="00:02:07.93" resultid="109549" heatid="110794" lane="0" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.22" />
                    <SPLIT distance="50" swimtime="00:00:55.85" />
                    <SPLIT distance="75" swimtime="00:01:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="122" reactiontime="+82" swimtime="00:04:00.39" resultid="109550" heatid="110807" lane="9" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.71" />
                    <SPLIT distance="50" swimtime="00:00:54.19" />
                    <SPLIT distance="75" swimtime="00:01:23.51" />
                    <SPLIT distance="100" swimtime="00:02:59.50" />
                    <SPLIT distance="125" swimtime="00:02:27.61" />
                    <SPLIT distance="175" swimtime="00:03:31.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Grażyna" gender="F" lastname="Drela" nation="POL" athleteid="109525">
              <RESULTS>
                <RESULT eventid="98777" points="320" reactiontime="+79" swimtime="00:00:33.95" resultid="109526" heatid="110589" lane="8" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="258" reactiontime="+83" swimtime="00:03:11.30" resultid="109527" heatid="110615" lane="4" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.63" />
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="75" swimtime="00:01:05.33" />
                    <SPLIT distance="100" swimtime="00:01:30.68" />
                    <SPLIT distance="125" swimtime="00:01:55.84" />
                    <SPLIT distance="150" swimtime="00:02:22.83" />
                    <SPLIT distance="175" swimtime="00:02:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="306" reactiontime="+82" swimtime="00:03:19.62" resultid="109528" heatid="110663" lane="7" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.78" />
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                    <SPLIT distance="75" swimtime="00:01:10.05" />
                    <SPLIT distance="100" swimtime="00:01:35.40" />
                    <SPLIT distance="125" swimtime="00:02:01.26" />
                    <SPLIT distance="150" swimtime="00:02:27.89" />
                    <SPLIT distance="175" swimtime="00:02:53.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="296" reactiontime="+90" swimtime="00:01:25.00" resultid="109529" heatid="110693" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.41" />
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="75" swimtime="00:01:03.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="308" reactiontime="+96" swimtime="00:01:32.32" resultid="109530" heatid="110723" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.70" />
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                    <SPLIT distance="75" swimtime="00:01:07.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="249" reactiontime="+94" swimtime="00:00:38.73" resultid="109531" heatid="110737" lane="3" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="304" swimtime="00:00:42.80" resultid="109532" heatid="110821" lane="0" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" license="100115700384" athleteid="109551">
              <RESULTS>
                <RESULT eventid="98830" points="520" reactiontime="+79" swimtime="00:02:16.30" resultid="109552" heatid="110628" lane="3" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="75" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:04.52" />
                    <SPLIT distance="125" swimtime="00:01:23.94" />
                    <SPLIT distance="150" swimtime="00:01:43.97" />
                    <SPLIT distance="175" swimtime="00:02:00.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="535" reactiontime="+81" swimtime="00:17:24.34" resultid="109553" heatid="110641" lane="4" entrytime="00:17:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.37" />
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="75" swimtime="00:00:47.75" />
                    <SPLIT distance="100" swimtime="00:01:04.88" />
                    <SPLIT distance="125" swimtime="00:01:22.08" />
                    <SPLIT distance="150" swimtime="00:01:39.32" />
                    <SPLIT distance="175" swimtime="00:01:56.59" />
                    <SPLIT distance="200" swimtime="00:02:14.11" />
                    <SPLIT distance="225" swimtime="00:02:31.59" />
                    <SPLIT distance="250" swimtime="00:02:48.97" />
                    <SPLIT distance="275" swimtime="00:03:06.44" />
                    <SPLIT distance="300" swimtime="00:03:23.98" />
                    <SPLIT distance="325" swimtime="00:03:41.58" />
                    <SPLIT distance="350" swimtime="00:03:59.27" />
                    <SPLIT distance="375" swimtime="00:04:16.77" />
                    <SPLIT distance="400" swimtime="00:04:34.28" />
                    <SPLIT distance="425" swimtime="00:04:51.84" />
                    <SPLIT distance="450" swimtime="00:05:09.56" />
                    <SPLIT distance="475" swimtime="00:05:27.18" />
                    <SPLIT distance="500" swimtime="00:05:44.72" />
                    <SPLIT distance="525" swimtime="00:06:02.20" />
                    <SPLIT distance="550" swimtime="00:06:19.71" />
                    <SPLIT distance="575" swimtime="00:06:37.47" />
                    <SPLIT distance="600" swimtime="00:06:54.94" />
                    <SPLIT distance="625" swimtime="00:07:12.34" />
                    <SPLIT distance="650" swimtime="00:07:29.91" />
                    <SPLIT distance="675" swimtime="00:07:47.54" />
                    <SPLIT distance="700" swimtime="00:08:05.06" />
                    <SPLIT distance="725" swimtime="00:08:22.59" />
                    <SPLIT distance="750" swimtime="00:08:40.10" />
                    <SPLIT distance="775" swimtime="00:08:57.70" />
                    <SPLIT distance="800" swimtime="00:09:15.37" />
                    <SPLIT distance="825" swimtime="00:09:32.97" />
                    <SPLIT distance="850" swimtime="00:09:50.75" />
                    <SPLIT distance="875" swimtime="00:10:08.53" />
                    <SPLIT distance="900" swimtime="00:10:26.27" />
                    <SPLIT distance="925" swimtime="00:10:43.99" />
                    <SPLIT distance="950" swimtime="00:11:01.71" />
                    <SPLIT distance="975" swimtime="00:11:19.43" />
                    <SPLIT distance="1000" swimtime="00:11:36.83" />
                    <SPLIT distance="1025" swimtime="00:11:54.37" />
                    <SPLIT distance="1050" swimtime="00:12:12.11" />
                    <SPLIT distance="1075" swimtime="00:12:29.83" />
                    <SPLIT distance="1100" swimtime="00:12:47.29" />
                    <SPLIT distance="1125" swimtime="00:13:04.80" />
                    <SPLIT distance="1150" swimtime="00:13:22.38" />
                    <SPLIT distance="1175" swimtime="00:13:39.89" />
                    <SPLIT distance="1200" swimtime="00:13:57.59" />
                    <SPLIT distance="1225" swimtime="00:14:15.22" />
                    <SPLIT distance="1250" swimtime="00:14:32.72" />
                    <SPLIT distance="1275" swimtime="00:14:50.46" />
                    <SPLIT distance="1300" swimtime="00:15:08.00" />
                    <SPLIT distance="1325" swimtime="00:15:25.30" />
                    <SPLIT distance="1350" swimtime="00:15:42.79" />
                    <SPLIT distance="1375" swimtime="00:16:00.24" />
                    <SPLIT distance="1400" swimtime="00:16:17.88" />
                    <SPLIT distance="1425" swimtime="00:16:35.41" />
                    <SPLIT distance="1450" swimtime="00:16:52.68" />
                    <SPLIT distance="1475" swimtime="00:17:09.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="481" reactiontime="+71" swimtime="00:02:33.76" resultid="109554" heatid="110670" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.56" />
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="75" swimtime="00:00:53.48" />
                    <SPLIT distance="100" swimtime="00:01:13.39" />
                    <SPLIT distance="125" swimtime="00:01:33.60" />
                    <SPLIT distance="150" swimtime="00:01:53.73" />
                    <SPLIT distance="175" swimtime="00:02:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="518" reactiontime="+78" swimtime="00:02:15.17" resultid="109555" heatid="110713" lane="3" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.58" />
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                    <SPLIT distance="75" swimtime="00:00:46.34" />
                    <SPLIT distance="100" swimtime="00:01:03.60" />
                    <SPLIT distance="125" swimtime="00:01:20.64" />
                    <SPLIT distance="150" swimtime="00:01:38.26" />
                    <SPLIT distance="175" swimtime="00:01:56.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="535" reactiontime="+70" swimtime="00:02:02.38" resultid="109556" heatid="110778" lane="7" entrytime="00:01:59.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                    <SPLIT distance="75" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:00:59.51" />
                    <SPLIT distance="125" swimtime="00:01:15.28" />
                    <SPLIT distance="150" swimtime="00:01:31.35" />
                    <SPLIT distance="175" swimtime="00:01:47.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="487" reactiontime="+74" swimtime="00:04:59.20" resultid="109557" heatid="110792" lane="5" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                    <SPLIT distance="75" swimtime="00:00:47.47" />
                    <SPLIT distance="100" swimtime="00:01:05.03" />
                    <SPLIT distance="125" swimtime="00:01:25.74" />
                    <SPLIT distance="150" swimtime="00:01:45.90" />
                    <SPLIT distance="175" swimtime="00:02:05.80" />
                    <SPLIT distance="200" swimtime="00:02:25.81" />
                    <SPLIT distance="225" swimtime="00:02:46.98" />
                    <SPLIT distance="250" swimtime="00:03:08.41" />
                    <SPLIT distance="275" swimtime="00:03:29.94" />
                    <SPLIT distance="300" swimtime="00:03:51.52" />
                    <SPLIT distance="325" swimtime="00:04:09.32" />
                    <SPLIT distance="350" swimtime="00:04:26.35" />
                    <SPLIT distance="375" swimtime="00:04:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="484" swimtime="00:01:01.69" resultid="109558" heatid="110805" lane="9" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="75" swimtime="00:00:44.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="548" reactiontime="+74" swimtime="00:04:19.23" resultid="109559" heatid="110843" lane="3" entrytime="00:04:19.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="75" swimtime="00:00:46.03" />
                    <SPLIT distance="100" swimtime="00:01:02.71" />
                    <SPLIT distance="125" swimtime="00:01:19.31" />
                    <SPLIT distance="150" swimtime="00:01:36.06" />
                    <SPLIT distance="175" swimtime="00:01:52.75" />
                    <SPLIT distance="200" swimtime="00:02:09.70" />
                    <SPLIT distance="225" swimtime="00:02:26.30" />
                    <SPLIT distance="250" swimtime="00:02:43.08" />
                    <SPLIT distance="275" swimtime="00:02:59.48" />
                    <SPLIT distance="300" swimtime="00:03:15.95" />
                    <SPLIT distance="325" swimtime="00:03:32.12" />
                    <SPLIT distance="350" swimtime="00:03:48.27" />
                    <SPLIT distance="375" swimtime="00:04:04.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="Tomaszewski" nation="POL" athleteid="109560">
              <RESULTS>
                <RESULT eventid="98798" points="472" swimtime="00:00:26.02" resultid="109561" heatid="110608" lane="9" entrytime="00:00:27.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="438" reactiontime="+68" swimtime="00:00:29.25" resultid="109562" heatid="110659" lane="2" entrytime="00:00:30.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="462" reactiontime="+68" swimtime="00:01:03.24" resultid="109563" heatid="110762" lane="6" entrytime="00:01:09.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.19" />
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                    <SPLIT distance="75" swimtime="00:00:46.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="435" reactiontime="+41" swimtime="00:02:11.10" resultid="109564" heatid="110774" lane="6" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="75" swimtime="00:00:45.86" />
                    <SPLIT distance="100" swimtime="00:01:02.88" />
                    <SPLIT distance="125" swimtime="00:01:19.44" />
                    <SPLIT distance="150" swimtime="00:01:36.85" />
                    <SPLIT distance="175" swimtime="00:01:54.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="390" reactiontime="+70" swimtime="00:02:24.55" resultid="109565" heatid="110815" lane="6" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.92" />
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="75" swimtime="00:00:50.00" />
                    <SPLIT distance="100" swimtime="00:01:08.46" />
                    <SPLIT distance="125" swimtime="00:01:27.77" />
                    <SPLIT distance="150" swimtime="00:01:46.44" />
                    <SPLIT distance="175" swimtime="00:02:05.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-05-14" firstname="Przemysław" gender="M" lastname="Isalski" nation="POL" athleteid="109520">
              <RESULTS>
                <RESULT eventid="98891" points="371" reactiontime="+84" swimtime="00:10:16.92" resultid="109521" heatid="110636" lane="8" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.81" />
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="75" swimtime="00:00:51.87" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="125" swimtime="00:01:29.00" />
                    <SPLIT distance="150" swimtime="00:01:47.92" />
                    <SPLIT distance="175" swimtime="00:02:06.89" />
                    <SPLIT distance="200" swimtime="00:02:26.13" />
                    <SPLIT distance="225" swimtime="00:02:45.22" />
                    <SPLIT distance="250" swimtime="00:03:04.85" />
                    <SPLIT distance="275" swimtime="00:03:24.32" />
                    <SPLIT distance="300" swimtime="00:03:43.97" />
                    <SPLIT distance="325" swimtime="00:04:03.43" />
                    <SPLIT distance="350" swimtime="00:04:23.32" />
                    <SPLIT distance="375" swimtime="00:04:42.88" />
                    <SPLIT distance="400" swimtime="00:05:02.49" />
                    <SPLIT distance="425" swimtime="00:05:21.91" />
                    <SPLIT distance="450" swimtime="00:05:41.46" />
                    <SPLIT distance="475" swimtime="00:06:00.90" />
                    <SPLIT distance="500" swimtime="00:06:20.57" />
                    <SPLIT distance="525" swimtime="00:06:40.21" />
                    <SPLIT distance="550" swimtime="00:07:00.00" />
                    <SPLIT distance="575" swimtime="00:07:19.78" />
                    <SPLIT distance="600" swimtime="00:07:39.88" />
                    <SPLIT distance="625" swimtime="00:07:59.12" />
                    <SPLIT distance="650" swimtime="00:08:19.20" />
                    <SPLIT distance="675" swimtime="00:08:38.84" />
                    <SPLIT distance="700" swimtime="00:08:58.72" />
                    <SPLIT distance="725" swimtime="00:09:18.70" />
                    <SPLIT distance="750" swimtime="00:09:38.55" />
                    <SPLIT distance="775" swimtime="00:09:57.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="360" reactiontime="+88" swimtime="00:02:49.31" resultid="109522" heatid="110668" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.89" />
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="75" swimtime="00:01:00.63" />
                    <SPLIT distance="100" swimtime="00:01:22.28" />
                    <SPLIT distance="125" swimtime="00:01:43.90" />
                    <SPLIT distance="150" swimtime="00:02:05.69" />
                    <SPLIT distance="175" swimtime="00:02:27.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="393" swimtime="00:02:15.66" resultid="109523" heatid="110775" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.66" />
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="75" swimtime="00:00:47.32" />
                    <SPLIT distance="100" swimtime="00:01:04.18" />
                    <SPLIT distance="125" swimtime="00:01:21.30" />
                    <SPLIT distance="150" swimtime="00:01:39.07" />
                    <SPLIT distance="175" swimtime="00:01:57.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="395" reactiontime="+94" swimtime="00:04:49.24" resultid="109524" heatid="110845" lane="1" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="75" swimtime="00:00:49.83" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="125" swimtime="00:01:25.90" />
                    <SPLIT distance="150" swimtime="00:01:44.44" />
                    <SPLIT distance="175" swimtime="00:02:02.80" />
                    <SPLIT distance="200" swimtime="00:02:21.20" />
                    <SPLIT distance="225" swimtime="00:02:39.77" />
                    <SPLIT distance="250" swimtime="00:02:58.25" />
                    <SPLIT distance="275" swimtime="00:03:16.86" />
                    <SPLIT distance="300" swimtime="00:03:35.47" />
                    <SPLIT distance="325" swimtime="00:03:53.97" />
                    <SPLIT distance="350" swimtime="00:04:12.43" />
                    <SPLIT distance="375" swimtime="00:04:30.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-03" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" license="100115700350" athleteid="109580">
              <RESULTS>
                <RESULT eventid="106277" points="420" reactiontime="+91" swimtime="00:01:00.00" resultid="109581" heatid="110686" lane="1" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.95" />
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                    <SPLIT distance="75" swimtime="00:00:44.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="402" reactiontime="+76" swimtime="00:02:14.61" resultid="109582" heatid="110776" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.81" />
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="75" swimtime="00:00:48.19" />
                    <SPLIT distance="100" swimtime="00:01:05.64" />
                    <SPLIT distance="125" swimtime="00:01:23.17" />
                    <SPLIT distance="150" swimtime="00:01:40.73" />
                    <SPLIT distance="175" swimtime="00:01:58.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="109583" heatid="110802" lane="2" entrytime="00:01:12.00" />
                <RESULT eventid="99473" points="377" swimtime="00:04:53.60" resultid="109584" heatid="110844" lane="2" entrytime="00:04:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="75" swimtime="00:00:50.61" />
                    <SPLIT distance="100" swimtime="00:01:09.07" />
                    <SPLIT distance="125" swimtime="00:01:27.83" />
                    <SPLIT distance="150" swimtime="00:01:46.92" />
                    <SPLIT distance="175" swimtime="00:02:05.86" />
                    <SPLIT distance="200" swimtime="00:02:25.06" />
                    <SPLIT distance="225" swimtime="00:02:44.25" />
                    <SPLIT distance="250" swimtime="00:03:03.54" />
                    <SPLIT distance="275" swimtime="00:03:22.27" />
                    <SPLIT distance="300" swimtime="00:03:41.31" />
                    <SPLIT distance="325" swimtime="00:03:59.84" />
                    <SPLIT distance="350" swimtime="00:04:18.60" />
                    <SPLIT distance="375" swimtime="00:04:36.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" license="100115700346" athleteid="109512">
              <RESULTS>
                <RESULT eventid="98798" points="359" reactiontime="+83" swimtime="00:00:28.49" resultid="109513" heatid="110604" lane="4" entrytime="00:00:29.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="328" reactiontime="+92" swimtime="00:10:42.34" resultid="109514" heatid="110636" lane="6" entrytime="00:10:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.79" />
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="75" swimtime="00:00:54.90" />
                    <SPLIT distance="100" swimtime="00:01:14.64" />
                    <SPLIT distance="125" swimtime="00:01:34.46" />
                    <SPLIT distance="150" swimtime="00:01:54.65" />
                    <SPLIT distance="175" swimtime="00:02:14.62" />
                    <SPLIT distance="200" swimtime="00:02:34.50" />
                    <SPLIT distance="225" swimtime="00:02:54.44" />
                    <SPLIT distance="250" swimtime="00:03:14.91" />
                    <SPLIT distance="275" swimtime="00:03:35.36" />
                    <SPLIT distance="300" swimtime="00:03:56.05" />
                    <SPLIT distance="325" swimtime="00:04:16.77" />
                    <SPLIT distance="350" swimtime="00:04:37.06" />
                    <SPLIT distance="375" swimtime="00:04:57.44" />
                    <SPLIT distance="400" swimtime="00:05:18.05" />
                    <SPLIT distance="425" swimtime="00:05:38.41" />
                    <SPLIT distance="450" swimtime="00:05:58.88" />
                    <SPLIT distance="475" swimtime="00:06:19.67" />
                    <SPLIT distance="500" swimtime="00:06:40.49" />
                    <SPLIT distance="525" swimtime="00:07:00.63" />
                    <SPLIT distance="550" swimtime="00:07:21.31" />
                    <SPLIT distance="575" swimtime="00:07:41.71" />
                    <SPLIT distance="600" swimtime="00:08:02.46" />
                    <SPLIT distance="625" swimtime="00:08:22.50" />
                    <SPLIT distance="650" swimtime="00:08:43.38" />
                    <SPLIT distance="675" swimtime="00:09:03.57" />
                    <SPLIT distance="700" swimtime="00:09:23.62" />
                    <SPLIT distance="725" swimtime="00:09:43.61" />
                    <SPLIT distance="750" swimtime="00:10:04.47" />
                    <SPLIT distance="775" swimtime="00:10:23.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="322" reactiontime="+86" swimtime="00:00:32.39" resultid="109515" heatid="110657" lane="3" entrytime="00:00:33.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="332" reactiontime="+101" swimtime="00:01:13.13" resultid="109516" heatid="110701" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.30" />
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="75" swimtime="00:00:55.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="309" reactiontime="+79" swimtime="00:01:12.31" resultid="109517" heatid="110761" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.80" />
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="75" swimtime="00:00:55.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="300" reactiontime="+72" swimtime="00:02:37.70" resultid="109518" heatid="110814" lane="6" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="75" swimtime="00:00:57.51" />
                    <SPLIT distance="100" swimtime="00:01:17.69" />
                    <SPLIT distance="125" swimtime="00:01:37.91" />
                    <SPLIT distance="150" swimtime="00:01:58.71" />
                    <SPLIT distance="175" swimtime="00:02:18.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="330" swimtime="00:05:07.14" resultid="109519" heatid="110846" lane="6" entrytime="00:05:12.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.45" />
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="75" swimtime="00:00:53.08" />
                    <SPLIT distance="100" swimtime="00:01:12.17" />
                    <SPLIT distance="125" swimtime="00:01:31.25" />
                    <SPLIT distance="150" swimtime="00:01:50.75" />
                    <SPLIT distance="175" swimtime="00:02:10.44" />
                    <SPLIT distance="200" swimtime="00:02:30.46" />
                    <SPLIT distance="225" swimtime="00:02:49.89" />
                    <SPLIT distance="250" swimtime="00:03:09.62" />
                    <SPLIT distance="275" swimtime="00:03:29.05" />
                    <SPLIT distance="300" swimtime="00:03:49.29" />
                    <SPLIT distance="325" swimtime="00:04:08.96" />
                    <SPLIT distance="350" swimtime="00:04:29.13" />
                    <SPLIT distance="375" swimtime="00:04:48.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="482" reactiontime="+64" swimtime="00:01:55.37" resultid="109586" heatid="110719" lane="6" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.99" />
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                    <SPLIT distance="75" swimtime="00:00:43.58" />
                    <SPLIT distance="100" swimtime="00:01:00.71" />
                    <SPLIT distance="125" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:28.17" />
                    <SPLIT distance="175" swimtime="00:01:41.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109560" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="109572" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="109551" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="109520" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="99059" points="287" reactiontime="+78" swimtime="00:02:17.06" resultid="109587" heatid="110718" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.76" />
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="75" swimtime="00:00:50.38" />
                    <SPLIT distance="100" swimtime="00:01:11.41" />
                    <SPLIT distance="125" swimtime="00:01:28.83" />
                    <SPLIT distance="150" swimtime="00:01:49.59" />
                    <SPLIT distance="175" swimtime="00:02:02.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109512" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="109566" number="2" />
                    <RELAYPOSITION athleteid="109500" number="3" />
                    <RELAYPOSITION athleteid="109580" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="99250" points="477" reactiontime="+75" swimtime="00:01:45.65" resultid="109588" heatid="110783" lane="5" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.75" />
                    <SPLIT distance="50" swimtime="00:00:26.32" />
                    <SPLIT distance="75" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:00:53.18" />
                    <SPLIT distance="125" swimtime="00:01:05.66" />
                    <SPLIT distance="150" swimtime="00:01:19.86" />
                    <SPLIT distance="175" swimtime="00:01:32.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109560" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="109572" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="109551" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="109520" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="99250" points="312" reactiontime="+104" swimtime="00:02:01.78" resultid="109589" heatid="110782" lane="1" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="75" swimtime="00:00:44.22" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="125" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:01:33.58" />
                    <SPLIT distance="175" swimtime="00:01:47.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109512" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="109566" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="109500" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="109580" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="222" swimtime="00:02:16.24" resultid="109585" heatid="110630" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.01" />
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="75" swimtime="00:00:56.74" />
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="125" swimtime="00:01:28.96" />
                    <SPLIT distance="150" swimtime="00:01:44.43" />
                    <SPLIT distance="175" swimtime="00:01:59.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109505" number="1" />
                    <RELAYPOSITION athleteid="109525" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="109512" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="109580" number="4" reactiontime="-1" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="99441" points="254" reactiontime="+122" swimtime="00:02:22.85" resultid="109590" heatid="110837" lane="8" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.30" />
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                    <SPLIT distance="75" swimtime="00:01:06.43" />
                    <SPLIT distance="100" swimtime="00:01:29.00" />
                    <SPLIT distance="125" swimtime="00:01:42.37" />
                    <SPLIT distance="150" swimtime="00:01:57.56" />
                    <SPLIT distance="175" swimtime="00:02:09.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109505" number="1" reactiontime="+122" />
                    <RELAYPOSITION athleteid="109525" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="109551" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="109560" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="PO" clubid="106624" name="KU AZS UAM Poznań">
          <CONTACT city="Poznań" email="kukowalazs@gmail.com" name="Kowalik" phone="603965223" state="WLKP" street="Zagajnikowa 9" zip="61-602" />
          <ATHLETES>
            <ATHLETE birthdate="1981-12-27" firstname="Bartosz" gender="M" lastname="Jankowiak" nation="POL" athleteid="106630">
              <RESULTS>
                <RESULT eventid="98798" points="311" reactiontime="+58" swimtime="00:00:29.90" resultid="106631" heatid="110603" lane="4" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="256" swimtime="00:11:38.25" resultid="106632" heatid="110636" lane="9" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.75" />
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="75" swimtime="00:00:55.80" />
                    <SPLIT distance="100" swimtime="00:01:16.71" />
                    <SPLIT distance="125" swimtime="00:01:37.37" />
                    <SPLIT distance="150" swimtime="00:01:59.09" />
                    <SPLIT distance="175" swimtime="00:02:20.90" />
                    <SPLIT distance="200" swimtime="00:02:42.86" />
                    <SPLIT distance="225" swimtime="00:03:05.01" />
                    <SPLIT distance="250" swimtime="00:03:27.53" />
                    <SPLIT distance="275" swimtime="00:03:49.99" />
                    <SPLIT distance="300" swimtime="00:04:12.37" />
                    <SPLIT distance="325" swimtime="00:04:34.89" />
                    <SPLIT distance="350" swimtime="00:04:57.68" />
                    <SPLIT distance="375" swimtime="00:05:19.90" />
                    <SPLIT distance="400" swimtime="00:05:42.67" />
                    <SPLIT distance="425" swimtime="00:06:05.11" />
                    <SPLIT distance="450" swimtime="00:06:27.65" />
                    <SPLIT distance="475" swimtime="00:06:50.15" />
                    <SPLIT distance="500" swimtime="00:07:12.34" />
                    <SPLIT distance="525" swimtime="00:07:34.70" />
                    <SPLIT distance="550" swimtime="00:07:57.05" />
                    <SPLIT distance="575" swimtime="00:08:19.38" />
                    <SPLIT distance="600" swimtime="00:08:41.93" />
                    <SPLIT distance="625" swimtime="00:09:04.37" />
                    <SPLIT distance="650" swimtime="00:09:26.77" />
                    <SPLIT distance="675" swimtime="00:09:49.41" />
                    <SPLIT distance="700" swimtime="00:10:11.75" />
                    <SPLIT distance="725" swimtime="00:10:33.89" />
                    <SPLIT distance="750" swimtime="00:10:56.60" />
                    <SPLIT distance="775" swimtime="00:11:18.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="282" swimtime="00:01:08.53" resultid="106633" heatid="110683" lane="9" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.75" />
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="75" swimtime="00:00:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="259" swimtime="00:02:35.84" resultid="106634" heatid="110773" lane="0" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="75" swimtime="00:00:52.34" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="125" swimtime="00:01:33.54" />
                    <SPLIT distance="150" swimtime="00:01:54.85" />
                    <SPLIT distance="175" swimtime="00:02:16.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="272" reactiontime="+86" swimtime="00:05:27.54" resultid="106635" heatid="110847" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.50" />
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="75" swimtime="00:00:55.76" />
                    <SPLIT distance="100" swimtime="00:01:16.32" />
                    <SPLIT distance="125" swimtime="00:01:37.02" />
                    <SPLIT distance="150" swimtime="00:01:58.01" />
                    <SPLIT distance="175" swimtime="00:02:18.99" />
                    <SPLIT distance="200" swimtime="00:02:40.26" />
                    <SPLIT distance="225" swimtime="00:03:01.40" />
                    <SPLIT distance="250" swimtime="00:03:22.53" />
                    <SPLIT distance="275" swimtime="00:03:43.81" />
                    <SPLIT distance="300" swimtime="00:04:05.02" />
                    <SPLIT distance="325" swimtime="00:04:26.35" />
                    <SPLIT distance="350" swimtime="00:04:47.81" />
                    <SPLIT distance="375" swimtime="00:05:09.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-11" firstname="Magdalena" gender="F" lastname="Mieścicka" nation="POL" athleteid="106642">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="106643" heatid="110588" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="99004" status="DNS" swimtime="00:00:00.00" resultid="106644" heatid="110708" lane="0" entrytime="00:03:30.00" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="106645" heatid="110737" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="106646" heatid="110794" lane="2" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-25" firstname="Przemysław" gender="M" lastname="Tomczak" nation="POL" athleteid="106647">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="106648" heatid="110599" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="106649" heatid="110681" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="106650" heatid="110772" lane="0" entrytime="00:02:50.00" />
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="106651" heatid="110850" lane="2" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-02-17" firstname="Jerzy" gender="M" lastname="Gniazdowski" nation="POL" athleteid="106671">
              <RESULTS>
                <RESULT eventid="98798" points="468" reactiontime="+70" swimtime="00:00:26.08" resultid="106672" heatid="110612" lane="0" entrytime="00:00:25.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="474" reactiontime="+60" swimtime="00:00:57.63" resultid="106673" heatid="110688" lane="5" entrytime="00:00:56.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.58" />
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                    <SPLIT distance="75" swimtime="00:00:42.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="465" reactiontime="+58" swimtime="00:02:08.21" resultid="106674" heatid="110777" lane="5" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="75" swimtime="00:00:45.20" />
                    <SPLIT distance="100" swimtime="00:01:01.77" />
                    <SPLIT distance="125" swimtime="00:01:18.39" />
                    <SPLIT distance="150" swimtime="00:01:35.14" />
                    <SPLIT distance="175" swimtime="00:01:51.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="436" reactiontime="+58" swimtime="00:04:39.83" resultid="106675" heatid="110844" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="75" swimtime="00:00:47.22" />
                    <SPLIT distance="100" swimtime="00:01:04.89" />
                    <SPLIT distance="125" swimtime="00:01:22.16" />
                    <SPLIT distance="150" swimtime="00:01:39.77" />
                    <SPLIT distance="175" swimtime="00:01:57.71" />
                    <SPLIT distance="200" swimtime="00:02:15.92" />
                    <SPLIT distance="225" swimtime="00:02:33.50" />
                    <SPLIT distance="250" swimtime="00:02:51.53" />
                    <SPLIT distance="275" swimtime="00:03:09.42" />
                    <SPLIT distance="300" swimtime="00:03:27.60" />
                    <SPLIT distance="325" swimtime="00:03:45.97" />
                    <SPLIT distance="350" swimtime="00:04:04.37" />
                    <SPLIT distance="375" swimtime="00:04:22.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-05" firstname="Piotr" gender="M" lastname="Kowalik" nation="POL" license="103315700017" athleteid="106652">
              <RESULTS>
                <RESULT eventid="98798" points="520" reactiontime="+63" swimtime="00:00:25.19" resultid="106653" heatid="110613" lane="5" entrytime="00:00:23.79">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="534" reactiontime="+62" swimtime="00:00:27.38" resultid="106654" heatid="110660" lane="4" entrytime="00:00:26.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="645" reactiontime="+57" swimtime="00:00:25.23" resultid="106655" heatid="110751" lane="4" entrytime="00:00:24.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="616" reactiontime="+55" swimtime="00:00:56.90" resultid="106656" heatid="110805" lane="4" entrytime="00:00:54.68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.51" />
                    <SPLIT distance="50" swimtime="00:00:25.47" />
                    <SPLIT distance="75" swimtime="00:00:40.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="Sterczyński" nation="POL" license="103315200002" athleteid="106657">
              <RESULTS>
                <RESULT eventid="98830" points="462" reactiontime="+76" swimtime="00:02:21.80" resultid="106658" heatid="110628" lane="0" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.35" />
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="75" swimtime="00:00:47.85" />
                    <SPLIT distance="100" swimtime="00:01:05.66" />
                    <SPLIT distance="125" swimtime="00:01:25.99" />
                    <SPLIT distance="150" swimtime="00:01:47.49" />
                    <SPLIT distance="175" swimtime="00:02:05.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="394" reactiontime="+72" swimtime="00:00:30.30" resultid="106659" heatid="110659" lane="3" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="496" swimtime="00:01:03.97" resultid="106660" heatid="110706" lane="0" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.05" />
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="75" swimtime="00:00:47.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="462" reactiontime="+71" swimtime="00:00:28.18" resultid="106661" heatid="110749" lane="5" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="425" reactiontime="+74" swimtime="00:01:05.02" resultid="106662" heatid="110763" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="75" swimtime="00:00:48.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="411" reactiontime="+72" swimtime="00:02:22.04" resultid="106663" heatid="110816" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.63" />
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="75" swimtime="00:00:50.30" />
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                    <SPLIT distance="125" swimtime="00:01:26.60" />
                    <SPLIT distance="150" swimtime="00:01:45.24" />
                    <SPLIT distance="175" swimtime="00:02:04.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-15" firstname="Marcin" gender="M" lastname="Tomczak" nation="POL" athleteid="106636">
              <RESULTS>
                <RESULT eventid="98798" points="320" reactiontime="+92" swimtime="00:00:29.59" resultid="106637" heatid="110607" lane="1" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" status="DNS" swimtime="00:00:00.00" resultid="106638" heatid="110641" lane="0" entrytime="00:21:00.00" />
                <RESULT eventid="106277" points="297" swimtime="00:01:07.29" resultid="106639" heatid="110685" lane="9" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.26" />
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="75" swimtime="00:00:48.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="306" reactiontime="+76" swimtime="00:02:27.36" resultid="106640" heatid="110774" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.09" />
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="75" swimtime="00:00:52.06" />
                    <SPLIT distance="100" swimtime="00:01:10.83" />
                    <SPLIT distance="125" swimtime="00:01:29.96" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                    <SPLIT distance="175" swimtime="00:02:08.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="304" reactiontime="+101" swimtime="00:05:15.43" resultid="106641" heatid="110846" lane="3" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="75" swimtime="00:00:53.60" />
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="125" swimtime="00:01:31.78" />
                    <SPLIT distance="150" swimtime="00:01:51.43" />
                    <SPLIT distance="175" swimtime="00:02:11.43" />
                    <SPLIT distance="200" swimtime="00:02:31.69" />
                    <SPLIT distance="225" swimtime="00:02:52.08" />
                    <SPLIT distance="250" swimtime="00:03:12.28" />
                    <SPLIT distance="275" swimtime="00:03:32.55" />
                    <SPLIT distance="300" swimtime="00:03:53.14" />
                    <SPLIT distance="325" swimtime="00:04:13.82" />
                    <SPLIT distance="350" swimtime="00:04:34.76" />
                    <SPLIT distance="375" swimtime="00:04:55.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="Sterczyńska" nation="POL" license="103315100003" athleteid="106664">
              <RESULTS>
                <RESULT eventid="98777" points="606" reactiontime="+72" swimtime="00:00:27.45" resultid="106665" heatid="110593" lane="7" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="483" reactiontime="+77" swimtime="00:00:32.70" resultid="106666" heatid="110650" lane="7" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="592" reactiontime="+82" swimtime="00:01:00.63" resultid="106667" heatid="110676" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.01" />
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="75" swimtime="00:00:44.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="525" swimtime="00:01:17.30" resultid="106668" heatid="110725" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.71" />
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="75" swimtime="00:00:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="500" reactiontime="+68" swimtime="00:00:30.71" resultid="106669" heatid="110740" lane="3" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="538" reactiontime="+73" swimtime="00:00:35.41" resultid="106670" heatid="110823" lane="5" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="Sztafeta dowolna mężczyzn" number="2">
              <RESULTS>
                <RESULT eventid="99250" points="436" reactiontime="+68" swimtime="00:01:48.89" resultid="106678" heatid="110784" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.00" />
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                    <SPLIT distance="75" swimtime="00:00:43.15" />
                    <SPLIT distance="100" swimtime="00:00:58.79" />
                    <SPLIT distance="125" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:24.78" />
                    <SPLIT distance="175" swimtime="00:01:36.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106630" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="106636" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="106657" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="106652" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="Sztafeta Zmienna mężczyzn" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="393" reactiontime="+71" swimtime="00:02:03.48" resultid="106679" heatid="110719" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.89" />
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                    <SPLIT distance="75" swimtime="00:00:48.07" />
                    <SPLIT distance="100" swimtime="00:01:09.92" />
                    <SPLIT distance="125" swimtime="00:01:21.13" />
                    <SPLIT distance="150" swimtime="00:01:34.98" />
                    <SPLIT distance="175" swimtime="00:01:48.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106630" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="106636" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="106657" number="3" reactiontime="+20" />
                    <RELAYPOSITION athleteid="106652" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="Sztafeta dowolna mix" number="1">
              <RESULTS>
                <RESULT eventid="98846" status="DNS" swimtime="00:00:00.00" resultid="106677" heatid="110632" lane="2" entrytime="00:01:50.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106642" number="1" />
                    <RELAYPOSITION athleteid="106664" number="2" />
                    <RELAYPOSITION athleteid="106657" number="3" />
                    <RELAYPOSITION athleteid="106652" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="Sztafeta Zmienna mix" number="1">
              <RESULTS>
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="106676" heatid="110838" lane="8" entrytime="00:02:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106657" number="1" />
                    <RELAYPOSITION athleteid="106664" number="2" />
                    <RELAYPOSITION athleteid="106652" number="3" />
                    <RELAYPOSITION athleteid="106642" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="LAT" clubid="106409" name="LATVIA">
          <ATHLETES>
            <ATHLETE birthdate="1955-05-17" firstname="RAIMONDS" gender="M" lastname="GARENCIKS" nation="LAT" athleteid="106410">
              <RESULTS>
                <RESULT eventid="106256" points="262" reactiontime="+117" swimtime="00:22:03.86" resultid="106411" heatid="110642" lane="4" entrytime="00:21:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.07" />
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="75" swimtime="00:00:58.86" />
                    <SPLIT distance="100" swimtime="00:01:19.70" />
                    <SPLIT distance="125" swimtime="00:01:40.73" />
                    <SPLIT distance="150" swimtime="00:02:01.81" />
                    <SPLIT distance="175" swimtime="00:02:23.84" />
                    <SPLIT distance="200" swimtime="00:02:45.37" />
                    <SPLIT distance="225" swimtime="00:03:06.82" />
                    <SPLIT distance="250" swimtime="00:03:28.76" />
                    <SPLIT distance="275" swimtime="00:03:50.37" />
                    <SPLIT distance="300" swimtime="00:04:12.34" />
                    <SPLIT distance="325" swimtime="00:04:34.63" />
                    <SPLIT distance="350" swimtime="00:04:56.22" />
                    <SPLIT distance="375" swimtime="00:05:18.78" />
                    <SPLIT distance="400" swimtime="00:05:40.79" />
                    <SPLIT distance="425" swimtime="00:06:03.04" />
                    <SPLIT distance="450" swimtime="00:06:25.41" />
                    <SPLIT distance="475" swimtime="00:06:47.28" />
                    <SPLIT distance="500" swimtime="00:07:09.66" />
                    <SPLIT distance="525" swimtime="00:07:31.84" />
                    <SPLIT distance="550" swimtime="00:07:54.06" />
                    <SPLIT distance="575" swimtime="00:09:01.50" />
                    <SPLIT distance="600" swimtime="00:08:38.95" />
                    <SPLIT distance="625" swimtime="00:09:46.37" />
                    <SPLIT distance="650" swimtime="00:09:23.94" />
                    <SPLIT distance="675" swimtime="00:10:31.27" />
                    <SPLIT distance="700" swimtime="00:10:08.71" />
                    <SPLIT distance="725" swimtime="00:11:15.88" />
                    <SPLIT distance="750" swimtime="00:10:53.86" />
                    <SPLIT distance="775" swimtime="00:12:01.51" />
                    <SPLIT distance="800" swimtime="00:11:39.01" />
                    <SPLIT distance="825" swimtime="00:12:46.49" />
                    <SPLIT distance="850" swimtime="00:12:23.86" />
                    <SPLIT distance="875" swimtime="00:13:31.08" />
                    <SPLIT distance="900" swimtime="00:13:08.92" />
                    <SPLIT distance="925" swimtime="00:14:15.92" />
                    <SPLIT distance="950" swimtime="00:13:53.77" />
                    <SPLIT distance="1000" swimtime="00:14:38.60" />
                    <SPLIT distance="1025" swimtime="00:15:01.14" />
                    <SPLIT distance="1050" swimtime="00:15:23.46" />
                    <SPLIT distance="1075" swimtime="00:15:45.95" />
                    <SPLIT distance="1100" swimtime="00:16:08.50" />
                    <SPLIT distance="1125" swimtime="00:16:30.91" />
                    <SPLIT distance="1150" swimtime="00:16:53.52" />
                    <SPLIT distance="1175" swimtime="00:17:16.02" />
                    <SPLIT distance="1200" swimtime="00:17:38.19" />
                    <SPLIT distance="1225" swimtime="00:18:00.30" />
                    <SPLIT distance="1250" swimtime="00:18:22.22" />
                    <SPLIT distance="1275" swimtime="00:18:44.29" />
                    <SPLIT distance="1300" swimtime="00:19:06.33" />
                    <SPLIT distance="1325" swimtime="00:19:28.41" />
                    <SPLIT distance="1350" swimtime="00:19:50.87" />
                    <SPLIT distance="1375" swimtime="00:20:13.03" />
                    <SPLIT distance="1400" swimtime="00:20:35.41" />
                    <SPLIT distance="1425" swimtime="00:20:58.09" />
                    <SPLIT distance="1450" swimtime="00:21:20.80" />
                    <SPLIT distance="1475" swimtime="00:21:42.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="255" swimtime="00:02:36.50" resultid="106412" heatid="110773" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.92" />
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="75" swimtime="00:00:54.54" />
                    <SPLIT distance="100" swimtime="00:01:14.05" />
                    <SPLIT distance="125" swimtime="00:01:34.10" />
                    <SPLIT distance="150" swimtime="00:01:54.92" />
                    <SPLIT distance="175" swimtime="00:02:16.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="260" swimtime="00:05:32.19" resultid="106413" heatid="110847" lane="6" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.02" />
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="75" swimtime="00:00:57.48" />
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                    <SPLIT distance="125" swimtime="00:01:38.74" />
                    <SPLIT distance="150" swimtime="00:01:59.87" />
                    <SPLIT distance="175" swimtime="00:02:21.07" />
                    <SPLIT distance="200" swimtime="00:02:42.18" />
                    <SPLIT distance="225" swimtime="00:03:03.54" />
                    <SPLIT distance="250" swimtime="00:03:24.94" />
                    <SPLIT distance="275" swimtime="00:03:46.53" />
                    <SPLIT distance="300" swimtime="00:04:08.19" />
                    <SPLIT distance="325" swimtime="00:04:29.96" />
                    <SPLIT distance="350" swimtime="00:04:51.33" />
                    <SPLIT distance="375" swimtime="00:05:12.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06614" nation="POL" region="WAR" clubid="107159" name="Legia Warszawa">
          <CONTACT email="janek@plywanielegia.pl" name="Peńsko" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1986-03-05" firstname="Robert" gender="M" lastname="Majchrzak" nation="POL" athleteid="107194">
              <RESULTS>
                <RESULT eventid="98798" points="189" reactiontime="+105" swimtime="00:00:35.25" resultid="107195" heatid="110597" lane="3" entrytime="00:00:39.59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-28" firstname="Jan" gender="M" lastname="Chmura" nation="POL" athleteid="107179">
              <RESULTS>
                <RESULT eventid="98798" points="492" reactiontime="+66" swimtime="00:00:25.66" resultid="107180" heatid="110610" lane="7" entrytime="00:00:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="107181" heatid="110700" lane="4" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-02" firstname="Władysław" gender="M" lastname="Surała" nation="POL" athleteid="107211">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="107212" heatid="110597" lane="2" entrytime="00:00:39.61" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-16" firstname="Jacek" gender="M" lastname="Kaczyński" nation="POL" athleteid="107198">
              <RESULTS>
                <RESULT eventid="98798" points="617" reactiontime="+75" swimtime="00:00:23.79" resultid="107199" heatid="110613" lane="4" entrytime="00:00:23.51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="622" reactiontime="+42" swimtime="00:00:25.53" resultid="107200" heatid="110751" lane="6" entrytime="00:00:25.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-09" firstname="Łukasz" gender="M" lastname="Drzewiński" nation="POL" athleteid="107253">
              <RESULTS>
                <RESULT eventid="98891" status="DNS" swimtime="00:00:00.00" resultid="107254" heatid="110637" lane="6" />
                <RESULT eventid="98924" points="365" reactiontime="+76" swimtime="00:00:31.07" resultid="107255" heatid="110659" lane="6" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="400" reactiontime="+64" swimtime="00:02:43.49" resultid="107256" heatid="110670" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.57" />
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="75" swimtime="00:00:53.45" />
                    <SPLIT distance="100" swimtime="00:01:13.74" />
                    <SPLIT distance="125" swimtime="00:01:34.68" />
                    <SPLIT distance="150" swimtime="00:01:57.30" />
                    <SPLIT distance="175" swimtime="00:02:19.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="449" swimtime="00:01:12.59" resultid="107257" heatid="110734" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.89" />
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="75" swimtime="00:00:52.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="485" reactiontime="+76" swimtime="00:00:27.74" resultid="107258" heatid="110750" lane="1" entrytime="00:00:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-03-22" firstname="Mariusz" gender="M" lastname="Mikołajewski" nation="POL" athleteid="107186">
              <RESULTS>
                <RESULT eventid="98798" points="593" reactiontime="+74" swimtime="00:00:24.11" resultid="107187" heatid="110612" lane="6" entrytime="00:00:24.69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="577" reactiontime="+78" swimtime="00:02:11.63" resultid="107188" heatid="110628" lane="2" entrytime="00:02:19.69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.79" />
                    <SPLIT distance="50" swimtime="00:00:27.84" />
                    <SPLIT distance="75" swimtime="00:00:45.41" />
                    <SPLIT distance="100" swimtime="00:01:02.62" />
                    <SPLIT distance="125" swimtime="00:01:21.23" />
                    <SPLIT distance="150" swimtime="00:01:40.30" />
                    <SPLIT distance="175" swimtime="00:01:56.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="489" reactiontime="+76" swimtime="00:00:28.19" resultid="107189" heatid="110660" lane="7" entrytime="00:00:28.69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="642" reactiontime="+86" swimtime="00:00:58.71" resultid="107190" heatid="110706" lane="3" entrytime="00:01:00.69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.05" />
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                    <SPLIT distance="75" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="578" reactiontime="+79" swimtime="00:00:26.17" resultid="107191" heatid="110741" lane="2">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-03-27" firstname="Agata" gender="F" lastname="Korc" nation="POL" athleteid="107217">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="107218" heatid="110593" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="106294" status="DNS" swimtime="00:00:00.00" resultid="107219" heatid="110650" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="107220" heatid="110695" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="107221" heatid="110740" lane="2" entrytime="00:00:30.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-10-11" firstname="Marta" gender="F" lastname="Majchrzak" nation="POL" athleteid="107259">
              <RESULTS>
                <RESULT eventid="98777" points="395" reactiontime="+91" swimtime="00:00:31.66" resultid="107260" heatid="110592" lane="1" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-09" firstname="Paweł" gender="M" lastname="Korzeniowski" nation="POL" athleteid="107240">
              <RESULTS>
                <RESULT eventid="98988" points="744" reactiontime="+74" swimtime="00:00:55.89" resultid="107241" heatid="110706" lane="4" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.22" />
                    <SPLIT distance="50" swimtime="00:00:25.65" />
                    <SPLIT distance="75" swimtime="00:00:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="682" reactiontime="+74" swimtime="00:02:03.33" resultid="107242" heatid="110713" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.27" />
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                    <SPLIT distance="75" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:01:00.25" />
                    <SPLIT distance="125" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:31.89" />
                    <SPLIT distance="175" swimtime="00:01:47.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="677" reactiontime="+71" swimtime="00:01:03.31" resultid="107243" heatid="110734" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="75" swimtime="00:00:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="687" reactiontime="+76" swimtime="00:01:52.57" resultid="107244" heatid="110778" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.07" />
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                    <SPLIT distance="75" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:00:55.23" />
                    <SPLIT distance="125" swimtime="00:01:10.03" />
                    <SPLIT distance="150" swimtime="00:01:25.03" />
                    <SPLIT distance="175" swimtime="00:01:39.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-07" firstname="Agnieszka" gender="F" lastname="Kaczmarek" nation="POL" athleteid="107225">
              <RESULTS>
                <RESULT eventid="98814" points="461" reactiontime="+93" swimtime="00:02:37.68" resultid="107226" heatid="110618" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.29" />
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="75" swimtime="00:00:52.70" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="125" swimtime="00:01:35.06" />
                    <SPLIT distance="150" swimtime="00:01:58.28" />
                    <SPLIT distance="175" swimtime="00:02:18.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="482" reactiontime="+73" swimtime="00:00:32.73" resultid="107227" heatid="110650" lane="6" entrytime="00:00:32.08">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="454" reactiontime="+78" swimtime="00:01:11.60" resultid="107229" heatid="110752" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.90" />
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="75" swimtime="00:00:52.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="443" reactiontime="+94" swimtime="00:02:25.29" resultid="107230" heatid="110768" lane="3" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.57" />
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="75" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:08.91" />
                    <SPLIT distance="125" swimtime="00:01:27.77" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                    <SPLIT distance="175" swimtime="00:02:06.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="441" reactiontime="+84" swimtime="00:02:36.58" resultid="107231" heatid="110809" lane="4" entrytime="00:02:35.08">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.89" />
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="75" swimtime="00:00:56.49" />
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                    <SPLIT distance="125" swimtime="00:01:37.44" />
                    <SPLIT distance="150" swimtime="00:01:58.09" />
                    <SPLIT distance="175" swimtime="00:02:17.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="412" reactiontime="+92" swimtime="00:05:15.09" resultid="107232" heatid="110839" lane="7" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.42" />
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="75" swimtime="00:00:52.86" />
                    <SPLIT distance="100" swimtime="00:01:12.33" />
                    <SPLIT distance="125" swimtime="00:01:31.94" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                    <SPLIT distance="175" swimtime="00:02:12.04" />
                    <SPLIT distance="200" swimtime="00:02:32.70" />
                    <SPLIT distance="225" swimtime="00:02:52.97" />
                    <SPLIT distance="250" swimtime="00:03:13.16" />
                    <SPLIT distance="275" swimtime="00:03:33.74" />
                    <SPLIT distance="300" swimtime="00:03:54.15" />
                    <SPLIT distance="325" swimtime="00:04:14.62" />
                    <SPLIT distance="350" swimtime="00:04:35.44" />
                    <SPLIT distance="375" swimtime="00:04:56.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="475" reactiontime="+95" swimtime="00:01:05.21" resultid="109605" heatid="110676" lane="7" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.24" />
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="75" swimtime="00:00:48.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-12" firstname="Filip" gender="M" lastname="Rowiński" nation="POL" athleteid="107175">
              <RESULTS>
                <RESULT eventid="98798" points="524" reactiontime="+65" swimtime="00:00:25.13" resultid="107176" heatid="110612" lane="5" entrytime="00:00:24.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="605" reactiontime="+66" swimtime="00:01:05.75" resultid="107177" heatid="110734" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.64" />
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="75" swimtime="00:00:47.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="657" reactiontime="+68" swimtime="00:00:29.04" resultid="107178" heatid="110834" lane="4" entrytime="00:00:28.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Marta" gender="F" lastname="Wilczęga" nation="POL" athleteid="110853" />
            <ATHLETE birthdate="1976-11-12" firstname="Marcin" gender="M" lastname="Podhorecki" nation="POL" athleteid="107215">
              <RESULTS>
                <RESULT eventid="98798" points="213" reactiontime="+87" swimtime="00:00:33.92" resultid="107216" heatid="110597" lane="6" entrytime="00:00:39.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-28" firstname="Tomasz" gender="M" lastname="Wilczęga" nation="POL" athleteid="107245">
              <RESULTS>
                <RESULT eventid="98798" points="509" reactiontime="+72" swimtime="00:00:25.36" resultid="107246" heatid="110611" lane="3" entrytime="00:00:25.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="107247" heatid="110687" lane="3" entrytime="00:00:59.00" />
                <RESULT eventid="98988" points="454" reactiontime="+61" swimtime="00:01:05.91" resultid="107248" heatid="110703" lane="5" entrytime="00:01:08.51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="75" swimtime="00:00:51.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="488" reactiontime="+64" swimtime="00:00:27.68" resultid="107249" heatid="110750" lane="8" entrytime="00:00:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-21" firstname="Krzysztof" gender="M" lastname="Spyra" nation="POL" athleteid="107250">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="107251" heatid="110609" lane="5" entrytime="00:00:26.50" />
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="107252" heatid="110687" lane="9" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" athleteid="107182">
              <RESULTS>
                <RESULT eventid="98798" points="483" reactiontime="+50" swimtime="00:00:25.82" resultid="107183" heatid="110611" lane="0" entrytime="00:00:25.91">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="428" reactiontime="+78" swimtime="00:01:07.21" resultid="107184" heatid="110703" lane="4" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.81" />
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="75" swimtime="00:00:50.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="411" reactiontime="+73" swimtime="00:00:29.31" resultid="107185" heatid="110749" lane="7" entrytime="00:00:28.95">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-26" firstname="Olga" gender="F" lastname="Surała" nation="POL" athleteid="107208">
              <RESULTS>
                <RESULT eventid="106294" points="447" reactiontime="+73" swimtime="00:00:33.57" resultid="107209" heatid="110650" lane="8" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="450" reactiontime="+71" swimtime="00:01:13.93" resultid="107210" heatid="110695" lane="8" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.26" />
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="75" swimtime="00:00:55.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-30" firstname="Aleksandra" gender="F" lastname="Cichowska-Majchrzak" nation="POL" athleteid="107206">
              <RESULTS>
                <RESULT eventid="98777" points="412" reactiontime="+73" swimtime="00:00:31.22" resultid="107207" heatid="110591" lane="5" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-10-13" firstname="Rafał" gender="M" lastname="Majchrzak" nation="POL" athleteid="107192">
              <RESULTS>
                <RESULT eventid="98798" points="229" reactiontime="+96" swimtime="00:00:33.10" resultid="107193" heatid="110597" lane="5" entrytime="00:00:39.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-01" firstname="Michał" gender="M" lastname="Kucharski" nation="POL" athleteid="107213">
              <RESULTS>
                <RESULT eventid="98798" points="161" reactiontime="+123" swimtime="00:00:37.19" resultid="107214" heatid="110597" lane="4" entrytime="00:00:39.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-27" firstname="Jan" gender="M" lastname="Peńsko" nation="POL" swrid="4060705" athleteid="107167">
              <RESULTS>
                <RESULT eventid="98830" points="544" reactiontime="+93" swimtime="00:02:14.27" resultid="107168" heatid="110619" lane="2">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                    <SPLIT distance="75" swimtime="00:00:45.42" />
                    <SPLIT distance="100" swimtime="00:01:02.94" />
                    <SPLIT distance="125" swimtime="00:01:22.05" />
                    <SPLIT distance="150" swimtime="00:01:42.38" />
                    <SPLIT distance="175" swimtime="00:01:59.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="521" reactiontime="+87" swimtime="00:09:11.03" resultid="107169" heatid="110635" lane="4" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.56" />
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="75" swimtime="00:00:48.65" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="125" swimtime="00:01:23.52" />
                    <SPLIT distance="150" swimtime="00:01:40.67" />
                    <SPLIT distance="175" swimtime="00:01:57.95" />
                    <SPLIT distance="200" swimtime="00:02:15.24" />
                    <SPLIT distance="225" swimtime="00:02:32.66" />
                    <SPLIT distance="250" swimtime="00:02:50.41" />
                    <SPLIT distance="275" swimtime="00:03:08.01" />
                    <SPLIT distance="300" swimtime="00:03:25.33" />
                    <SPLIT distance="325" swimtime="00:03:42.90" />
                    <SPLIT distance="350" swimtime="00:04:00.47" />
                    <SPLIT distance="375" swimtime="00:04:18.30" />
                    <SPLIT distance="400" swimtime="00:04:35.81" />
                    <SPLIT distance="425" swimtime="00:04:53.10" />
                    <SPLIT distance="450" swimtime="00:05:10.32" />
                    <SPLIT distance="475" swimtime="00:05:27.62" />
                    <SPLIT distance="500" swimtime="00:05:44.81" />
                    <SPLIT distance="525" swimtime="00:06:01.98" />
                    <SPLIT distance="550" swimtime="00:06:19.23" />
                    <SPLIT distance="575" swimtime="00:06:36.61" />
                    <SPLIT distance="600" swimtime="00:06:53.91" />
                    <SPLIT distance="625" swimtime="00:07:11.45" />
                    <SPLIT distance="650" swimtime="00:07:28.79" />
                    <SPLIT distance="675" swimtime="00:07:46.37" />
                    <SPLIT distance="700" swimtime="00:08:03.94" />
                    <SPLIT distance="725" swimtime="00:08:21.06" />
                    <SPLIT distance="750" swimtime="00:08:37.84" />
                    <SPLIT distance="775" swimtime="00:08:54.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="498" reactiontime="+77" swimtime="00:00:28.02" resultid="107170" heatid="110651" lane="8">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="484" reactiontime="+81" swimtime="00:02:18.21" resultid="107171" heatid="110709" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.96" />
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="75" swimtime="00:00:49.00" />
                    <SPLIT distance="100" swimtime="00:01:06.94" />
                    <SPLIT distance="125" swimtime="00:01:24.90" />
                    <SPLIT distance="150" swimtime="00:01:42.78" />
                    <SPLIT distance="175" swimtime="00:01:59.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="500" reactiontime="+75" swimtime="00:01:01.62" resultid="107172" heatid="110757" lane="8">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.60" />
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="75" swimtime="00:00:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="519" swimtime="00:04:52.86" resultid="107173" heatid="110788" lane="0">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.12" />
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="75" swimtime="00:00:50.11" />
                    <SPLIT distance="100" swimtime="00:01:09.30" />
                    <SPLIT distance="125" swimtime="00:01:29.46" />
                    <SPLIT distance="150" swimtime="00:01:48.14" />
                    <SPLIT distance="175" swimtime="00:02:06.16" />
                    <SPLIT distance="200" swimtime="00:02:24.41" />
                    <SPLIT distance="225" swimtime="00:02:44.73" />
                    <SPLIT distance="250" swimtime="00:03:05.08" />
                    <SPLIT distance="275" swimtime="00:03:25.55" />
                    <SPLIT distance="300" swimtime="00:03:46.50" />
                    <SPLIT distance="325" swimtime="00:04:04.09" />
                    <SPLIT distance="350" swimtime="00:04:20.54" />
                    <SPLIT distance="375" swimtime="00:04:36.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="456" reactiontime="+90" swimtime="00:02:17.16" resultid="107174" heatid="110816" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.70" />
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="75" swimtime="00:00:50.55" />
                    <SPLIT distance="100" swimtime="00:01:08.46" />
                    <SPLIT distance="125" swimtime="00:01:26.01" />
                    <SPLIT distance="150" swimtime="00:01:43.21" />
                    <SPLIT distance="175" swimtime="00:02:00.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-09" firstname="Jakub" gender="M" lastname="Dobies" nation="POL" athleteid="107196">
              <RESULTS>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="107197" heatid="110834" lane="2" entrytime="00:00:30.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" swrid="4043251" athleteid="107233">
              <RESULTS>
                <RESULT eventid="98924" points="607" reactiontime="+65" swimtime="00:00:26.23" resultid="107234" heatid="110660" lane="5" entrytime="00:00:26.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="543" reactiontime="+70" swimtime="00:02:13.06" resultid="107235" heatid="110709" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.55" />
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="75" swimtime="00:00:47.88" />
                    <SPLIT distance="100" swimtime="00:01:04.53" />
                    <SPLIT distance="125" swimtime="00:01:21.96" />
                    <SPLIT distance="150" swimtime="00:01:39.50" />
                    <SPLIT distance="175" swimtime="00:01:56.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="582" reactiontime="+78" swimtime="00:00:26.11" resultid="107236" heatid="110741" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="572" reactiontime="+65" swimtime="00:00:58.90" resultid="107237" heatid="110763" lane="4" entrytime="00:00:58.53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.15" />
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                    <SPLIT distance="75" swimtime="00:00:44.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="593" swimtime="00:00:57.63" resultid="107238" heatid="110797" lane="6">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                    <SPLIT distance="75" swimtime="00:00:42.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="504" reactiontime="+67" swimtime="00:02:12.73" resultid="107239" heatid="110816" lane="5" entrytime="00:02:10.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.07" />
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="75" swimtime="00:00:47.27" />
                    <SPLIT distance="100" swimtime="00:01:03.97" />
                    <SPLIT distance="125" swimtime="00:01:21.10" />
                    <SPLIT distance="150" swimtime="00:01:37.94" />
                    <SPLIT distance="175" swimtime="00:01:55.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="522" swimtime="00:09:10.58" resultid="110360" heatid="110639" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-11" firstname="Katarzyna" gender="F" lastname="Ptasińska" nation="POL" athleteid="107201">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="107202" heatid="110593" lane="2" entrytime="00:00:27.99" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="107203" heatid="110676" lane="6" entrytime="00:01:00.00" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="107204" heatid="110740" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="107205" heatid="110768" lane="1" entrytime="00:02:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-09-28" firstname="Jędrzej" gender="M" lastname="Sieczych" nation="POL" athleteid="107222">
              <RESULTS>
                <RESULT eventid="98798" points="382" reactiontime="+82" swimtime="00:00:27.92" resultid="107223" heatid="110606" lane="0" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="307" reactiontime="+72" swimtime="00:01:15.05" resultid="107224" heatid="110701" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="75" swimtime="00:00:57.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="633" reactiontime="+56" swimtime="00:01:36.20" resultid="107266" heatid="110784" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.29" />
                    <SPLIT distance="50" swimtime="00:00:25.20" />
                    <SPLIT distance="75" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:00:48.40" />
                    <SPLIT distance="125" swimtime="00:00:59.90" />
                    <SPLIT distance="150" swimtime="00:01:13.11" />
                    <SPLIT distance="175" swimtime="00:01:23.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107245" number="1" reactiontime="+56" />
                    <RELAYPOSITION athleteid="107186" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="107175" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="107198" number="4" reactiontime="+1" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="629" reactiontime="+62" swimtime="00:01:45.59" resultid="107268" heatid="110719" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.11" />
                    <SPLIT distance="50" swimtime="00:00:26.33" />
                    <SPLIT distance="75" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:00:57.93" />
                    <SPLIT distance="125" swimtime="00:01:08.18" />
                    <SPLIT distance="150" swimtime="00:01:21.17" />
                    <SPLIT distance="175" swimtime="00:01:32.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107233" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="107253" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="107240" number="3" reactiontime="+20" />
                    <RELAYPOSITION athleteid="107167" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99250" points="634" reactiontime="+73" swimtime="00:01:36.11" resultid="107265" heatid="110784" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:25.24" />
                    <SPLIT distance="75" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:00:48.95" />
                    <SPLIT distance="125" swimtime="00:01:00.93" />
                    <SPLIT distance="150" swimtime="00:01:14.52" />
                    <SPLIT distance="175" swimtime="00:01:24.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107167" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="107233" number="2" reactiontime="+2" />
                    <RELAYPOSITION athleteid="107182" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="107240" number="4" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="620" reactiontime="+73" swimtime="00:01:46.13" resultid="107267" heatid="110719" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                    <SPLIT distance="75" swimtime="00:00:40.40" />
                    <SPLIT distance="100" swimtime="00:00:56.40" />
                    <SPLIT distance="125" swimtime="00:01:07.51" />
                    <SPLIT distance="150" swimtime="00:01:21.54" />
                    <SPLIT distance="175" swimtime="00:01:33.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107186" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="107175" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="107198" number="3" reactiontime="+13" />
                    <RELAYPOSITION athleteid="107245" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99234" points="399" reactiontime="+61" swimtime="00:02:07.91" resultid="107269" heatid="110780" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.87" />
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="75" swimtime="00:00:44.05" />
                    <SPLIT distance="100" swimtime="00:01:00.52" />
                    <SPLIT distance="125" swimtime="00:01:18.09" />
                    <SPLIT distance="150" swimtime="00:01:38.74" />
                    <SPLIT distance="175" swimtime="00:01:52.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107259" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="107208" number="2" />
                    <RELAYPOSITION athleteid="107206" number="3" />
                    <RELAYPOSITION athleteid="107225" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99036" points="350" reactiontime="+72" swimtime="00:02:27.50" resultid="107270" heatid="110715" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.18" />
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="75" swimtime="00:00:57.12" />
                    <SPLIT distance="100" swimtime="00:01:24.25" />
                    <SPLIT distance="125" swimtime="00:01:38.19" />
                    <SPLIT distance="150" swimtime="00:01:55.82" />
                    <SPLIT distance="175" swimtime="00:02:11.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107208" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="107225" number="2" />
                    <RELAYPOSITION athleteid="107206" number="3" />
                    <RELAYPOSITION athleteid="107259" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" status="WDR" swimtime="00:00:00.00" resultid="107261" heatid="110632" lane="4" entrytime="00:01:45.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107186" number="1" />
                    <RELAYPOSITION athleteid="107175" number="2" />
                    <RELAYPOSITION athleteid="107208" number="3" />
                    <RELAYPOSITION athleteid="107201" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="434" reactiontime="+68" swimtime="00:01:59.52" resultid="107264" heatid="110838" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.67" />
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="75" swimtime="00:00:46.48" />
                    <SPLIT distance="100" swimtime="00:01:02.41" />
                    <SPLIT distance="125" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:01:28.53" />
                    <SPLIT distance="175" swimtime="00:01:43.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107167" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="107175" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="107225" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="107208" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT comment="O4/ III ZMIANA" eventid="98846" reactiontime="+75" status="DSQ" swimtime="00:00:00.00" resultid="107262" heatid="110632" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                    <SPLIT distance="75" swimtime="00:01:06.06" />
                    <SPLIT distance="100" swimtime="00:01:24.84" />
                    <SPLIT distance="125" swimtime="00:01:38.19" />
                    <SPLIT distance="150" swimtime="00:01:53.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107198" number="1" reactiontime="+75" status="DSQ" />
                    <RELAYPOSITION athleteid="107179" number="2" reactiontime="+64" status="DSQ" />
                    <RELAYPOSITION athleteid="107225" number="3" reactiontime="-4" status="DSQ" />
                    <RELAYPOSITION athleteid="110853" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="107263" heatid="110838" lane="4" entrytime="00:01:50.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107225" number="1" />
                    <RELAYPOSITION athleteid="107196" number="2" />
                    <RELAYPOSITION athleteid="107233" number="3" />
                    <RELAYPOSITION athleteid="107206" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="98846" points="247" reactiontime="+69" swimtime="00:02:11.62" resultid="107271" heatid="110631" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.27" />
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="75" swimtime="00:00:47.29" />
                    <SPLIT distance="100" swimtime="00:01:05.76" />
                    <SPLIT distance="125" swimtime="00:01:21.87" />
                    <SPLIT distance="150" swimtime="00:01:40.21" />
                    <SPLIT distance="175" swimtime="00:01:55.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107206" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="107194" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="107192" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="107259" number="4" reactiontime="+6" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="107958" name="Masters Białystok">
          <CONTACT email="mbzgloszenia@gmail.com" name="Dominika Michalik" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="107959">
              <RESULTS>
                <RESULT eventid="106254" points="465" reactiontime="+65" swimtime="00:19:46.81" resultid="107960" heatid="110640" lane="5" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.44" />
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="75" swimtime="00:00:53.55" />
                    <SPLIT distance="100" swimtime="00:01:12.76" />
                    <SPLIT distance="125" swimtime="00:01:31.87" />
                    <SPLIT distance="150" swimtime="00:01:51.21" />
                    <SPLIT distance="175" swimtime="00:02:10.52" />
                    <SPLIT distance="200" swimtime="00:02:30.23" />
                    <SPLIT distance="225" swimtime="00:02:49.62" />
                    <SPLIT distance="250" swimtime="00:03:09.04" />
                    <SPLIT distance="275" swimtime="00:03:28.78" />
                    <SPLIT distance="300" swimtime="00:03:48.65" />
                    <SPLIT distance="325" swimtime="00:04:08.28" />
                    <SPLIT distance="350" swimtime="00:04:28.20" />
                    <SPLIT distance="375" swimtime="00:04:47.82" />
                    <SPLIT distance="400" swimtime="00:05:07.70" />
                    <SPLIT distance="425" swimtime="00:05:27.78" />
                    <SPLIT distance="450" swimtime="00:05:47.56" />
                    <SPLIT distance="475" swimtime="00:06:07.29" />
                    <SPLIT distance="500" swimtime="00:06:27.07" />
                    <SPLIT distance="525" swimtime="00:06:46.55" />
                    <SPLIT distance="550" swimtime="00:07:06.35" />
                    <SPLIT distance="575" swimtime="00:07:26.05" />
                    <SPLIT distance="600" swimtime="00:07:45.98" />
                    <SPLIT distance="625" swimtime="00:08:05.81" />
                    <SPLIT distance="650" swimtime="00:08:25.75" />
                    <SPLIT distance="675" swimtime="00:08:45.51" />
                    <SPLIT distance="700" swimtime="00:09:05.41" />
                    <SPLIT distance="725" swimtime="00:09:25.25" />
                    <SPLIT distance="750" swimtime="00:09:45.19" />
                    <SPLIT distance="775" swimtime="00:10:05.14" />
                    <SPLIT distance="800" swimtime="00:10:24.90" />
                    <SPLIT distance="825" swimtime="00:10:45.11" />
                    <SPLIT distance="850" swimtime="00:11:05.21" />
                    <SPLIT distance="875" swimtime="00:11:25.45" />
                    <SPLIT distance="900" swimtime="00:11:45.33" />
                    <SPLIT distance="925" swimtime="00:12:05.36" />
                    <SPLIT distance="950" swimtime="00:12:25.47" />
                    <SPLIT distance="975" swimtime="00:12:45.74" />
                    <SPLIT distance="1000" swimtime="00:13:06.00" />
                    <SPLIT distance="1025" swimtime="00:13:26.17" />
                    <SPLIT distance="1050" swimtime="00:13:46.85" />
                    <SPLIT distance="1075" swimtime="00:14:06.97" />
                    <SPLIT distance="1100" swimtime="00:14:27.15" />
                    <SPLIT distance="1125" swimtime="00:14:47.38" />
                    <SPLIT distance="1150" swimtime="00:15:07.43" />
                    <SPLIT distance="1175" swimtime="00:15:27.46" />
                    <SPLIT distance="1200" swimtime="00:15:47.98" />
                    <SPLIT distance="1225" swimtime="00:16:07.45" />
                    <SPLIT distance="1250" swimtime="00:16:27.64" />
                    <SPLIT distance="1275" swimtime="00:16:47.62" />
                    <SPLIT distance="1300" swimtime="00:17:07.91" />
                    <SPLIT distance="1325" swimtime="00:17:27.86" />
                    <SPLIT distance="1350" swimtime="00:17:48.20" />
                    <SPLIT distance="1375" swimtime="00:18:08.09" />
                    <SPLIT distance="1400" swimtime="00:18:28.47" />
                    <SPLIT distance="1425" swimtime="00:18:48.89" />
                    <SPLIT distance="1450" swimtime="00:19:08.86" />
                    <SPLIT distance="1475" swimtime="00:19:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="448" swimtime="00:01:06.49" resultid="107961" heatid="110676" lane="9" entrytime="00:01:05.27">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.60" />
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="75" swimtime="00:00:49.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="482" reactiontime="+85" swimtime="00:02:21.29" resultid="107962" heatid="110768" lane="2" entrytime="00:02:19.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.66" />
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="75" swimtime="00:00:50.58" />
                    <SPLIT distance="100" swimtime="00:01:08.74" />
                    <SPLIT distance="125" swimtime="00:01:27.18" />
                    <SPLIT distance="150" swimtime="00:01:45.62" />
                    <SPLIT distance="175" swimtime="00:02:04.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="496" reactiontime="+77" swimtime="00:04:56.12" resultid="107963" heatid="110839" lane="5" entrytime="00:04:57.46">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.34" />
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="75" swimtime="00:00:52.39" />
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                    <SPLIT distance="125" swimtime="00:01:29.56" />
                    <SPLIT distance="150" swimtime="00:01:48.39" />
                    <SPLIT distance="175" swimtime="00:02:07.53" />
                    <SPLIT distance="200" swimtime="00:02:26.64" />
                    <SPLIT distance="225" swimtime="00:02:45.69" />
                    <SPLIT distance="250" swimtime="00:03:04.67" />
                    <SPLIT distance="275" swimtime="00:03:23.68" />
                    <SPLIT distance="300" swimtime="00:03:43.00" />
                    <SPLIT distance="325" swimtime="00:04:01.86" />
                    <SPLIT distance="350" swimtime="00:04:20.73" />
                    <SPLIT distance="375" swimtime="00:04:39.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Elżbieta" gender="F" lastname="Piwowarczyk" nation="POL" athleteid="107985">
              <RESULTS>
                <RESULT eventid="98777" points="335" reactiontime="+75" swimtime="00:00:33.46" resultid="107986" heatid="110589" lane="4" entrytime="00:00:34.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="268" reactiontime="+79" swimtime="00:03:08.83" resultid="107987" heatid="110616" lane="8" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.34" />
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                    <SPLIT distance="75" swimtime="00:01:06.09" />
                    <SPLIT distance="100" swimtime="00:01:30.69" />
                    <SPLIT distance="125" swimtime="00:01:58.51" />
                    <SPLIT distance="150" swimtime="00:02:26.61" />
                    <SPLIT distance="175" swimtime="00:02:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="248" reactiontime="+77" swimtime="00:00:40.81" resultid="107988" heatid="110648" lane="6" entrytime="00:00:40.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="323" swimtime="00:01:14.16" resultid="107989" heatid="110674" lane="9" entrytime="00:01:16.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.13" />
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                    <SPLIT distance="75" swimtime="00:00:54.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="247" reactiontime="+80" swimtime="00:01:27.60" resultid="107990" heatid="110755" lane="7" entrytime="00:01:29.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.95" />
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="75" swimtime="00:01:05.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="296" reactiontime="+94" swimtime="00:02:46.15" resultid="107991" heatid="110766" lane="1" entrytime="00:02:55.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.80" />
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="75" swimtime="00:00:57.93" />
                    <SPLIT distance="100" swimtime="00:01:19.14" />
                    <SPLIT distance="125" swimtime="00:01:40.68" />
                    <SPLIT distance="150" swimtime="00:02:02.75" />
                    <SPLIT distance="175" swimtime="00:02:24.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="255" reactiontime="+83" swimtime="00:03:07.85" resultid="107992" heatid="110808" lane="8" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.62" />
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="75" swimtime="00:01:07.83" />
                    <SPLIT distance="100" swimtime="00:01:31.52" />
                    <SPLIT distance="125" swimtime="00:01:55.56" />
                    <SPLIT distance="150" swimtime="00:02:19.62" />
                    <SPLIT distance="175" swimtime="00:02:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="276" reactiontime="+89" swimtime="00:06:00.18" resultid="107993" heatid="110841" lane="3" entrytime="00:06:05.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.22" />
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="75" swimtime="00:00:59.39" />
                    <SPLIT distance="100" swimtime="00:01:21.10" />
                    <SPLIT distance="125" swimtime="00:01:43.26" />
                    <SPLIT distance="150" swimtime="00:02:05.82" />
                    <SPLIT distance="175" swimtime="00:02:28.67" />
                    <SPLIT distance="200" swimtime="00:02:51.67" />
                    <SPLIT distance="225" swimtime="00:03:14.89" />
                    <SPLIT distance="250" swimtime="00:03:38.43" />
                    <SPLIT distance="275" swimtime="00:04:02.29" />
                    <SPLIT distance="300" swimtime="00:04:26.22" />
                    <SPLIT distance="325" swimtime="00:04:50.07" />
                    <SPLIT distance="350" swimtime="00:05:13.97" />
                    <SPLIT distance="375" swimtime="00:05:37.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Maciej" gender="M" lastname="Daszuta" nation="POL" athleteid="107964">
              <RESULTS>
                <RESULT eventid="98798" points="388" reactiontime="+70" swimtime="00:00:27.76" resultid="107965" heatid="110607" lane="4" entrytime="00:00:27.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="345" reactiontime="+68" swimtime="00:00:31.67" resultid="107966" heatid="110658" lane="6" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="333" reactiontime="+69" swimtime="00:01:13.05" resultid="107967" heatid="110702" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="75" swimtime="00:00:55.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="371" swimtime="00:01:17.37" resultid="107968" heatid="110732" lane="0" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.02" />
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="75" swimtime="00:00:56.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="107969" heatid="110761" lane="3" entrytime="00:01:14.00" />
                <RESULT comment="K4" eventid="99425" reactiontime="+66" status="DSQ" swimtime="00:00:00.00" resultid="107970" heatid="110832" lane="4" entrytime="00:00:34.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosław" gender="M" lastname="Matusik" nation="POL" athleteid="107971">
              <RESULTS>
                <RESULT eventid="98798" status="WDR" swimtime="00:00:00.00" resultid="107972" entrytime="00:00:33.00" />
                <RESULT eventid="98988" status="WDR" swimtime="00:00:00.00" resultid="107973" entrytime="00:01:24.80" />
                <RESULT eventid="99091" status="WDR" swimtime="00:00:00.00" resultid="107974" entrytime="00:01:29.80" />
                <RESULT eventid="99170" status="WDR" swimtime="00:00:00.00" resultid="107975" entrytime="00:00:35.90" />
                <RESULT eventid="99361" status="WDR" swimtime="00:00:00.00" resultid="107976" entrytime="00:01:45.00" />
                <RESULT eventid="99425" status="WDR" swimtime="00:00:00.00" resultid="107977" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LBL" clubid="107994" name="Masters Chełm">
          <CONTACT city="Chełm" email="wepa56@interia.pl" name="Wepa Wiesław" phone="663903089" state="LBL" street="Grunwaldzka 36" zip="22-100" />
          <ATHLETES>
            <ATHLETE birthdate="1941-10-11" firstname="Janusz" gender="M" lastname="G0lik" nation="POL" athleteid="107995">
              <RESULTS>
                <RESULT eventid="98956" points="99" reactiontime="+97" swimtime="00:04:19.90" resultid="107996" heatid="110666" lane="8" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.24" />
                    <SPLIT distance="50" swimtime="00:00:59.63" />
                    <SPLIT distance="75" swimtime="00:01:32.90" />
                    <SPLIT distance="100" swimtime="00:02:06.95" />
                    <SPLIT distance="125" swimtime="00:02:40.69" />
                    <SPLIT distance="150" swimtime="00:03:14.74" />
                    <SPLIT distance="175" swimtime="00:03:47.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="63" reactiontime="+107" swimtime="00:04:31.62" resultid="107997" heatid="110710" lane="7" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.39" />
                    <SPLIT distance="50" swimtime="00:01:02.17" />
                    <SPLIT distance="75" swimtime="00:01:37.26" />
                    <SPLIT distance="100" swimtime="00:02:12.75" />
                    <SPLIT distance="125" swimtime="00:02:50.07" />
                    <SPLIT distance="150" swimtime="00:03:26.37" />
                    <SPLIT distance="175" swimtime="00:04:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="157" reactiontime="+113" swimtime="00:01:43.06" resultid="107998" heatid="110728" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.43" />
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                    <SPLIT distance="75" swimtime="00:01:14.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="89" reactiontime="+95" swimtime="00:00:48.77" resultid="107999" heatid="110742" lane="3" entrytime="00:00:46.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="76" reactiontime="+104" swimtime="00:01:54.29" resultid="108000" heatid="110799" lane="8" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.82" />
                    <SPLIT distance="50" swimtime="00:00:56.41" />
                    <SPLIT distance="75" swimtime="00:01:25.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="154" swimtime="00:00:47.01" resultid="108001" heatid="110826" lane="6" entrytime="00:00:44.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KRA" nation="POL" region="MAL" clubid="108493" name="Masters Korona Kraków">
          <CONTACT city="Kraków" email="masterskorona@wp.pl" name="Mariola Kuliœ" phone="500677133" state="MA£" />
          <ATHLETES>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="108524">
              <RESULTS>
                <RESULT eventid="98814" points="316" reactiontime="+89" swimtime="00:02:58.82" resultid="108525" heatid="110616" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.01" />
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="75" swimtime="00:01:00.97" />
                    <SPLIT distance="100" swimtime="00:01:24.03" />
                    <SPLIT distance="125" swimtime="00:01:50.11" />
                    <SPLIT distance="150" swimtime="00:02:16.58" />
                    <SPLIT distance="175" swimtime="00:02:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="327" reactiontime="+67" swimtime="00:01:22.18" resultid="108526" heatid="110692" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.52" />
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="75" swimtime="00:01:02.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="306" reactiontime="+96" swimtime="00:06:24.84" resultid="108527" heatid="110786" lane="4" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.96" />
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="75" swimtime="00:01:00.98" />
                    <SPLIT distance="100" swimtime="00:01:23.46" />
                    <SPLIT distance="125" swimtime="00:01:49.83" />
                    <SPLIT distance="150" swimtime="00:02:14.97" />
                    <SPLIT distance="175" swimtime="00:02:40.17" />
                    <SPLIT distance="200" swimtime="00:03:05.24" />
                    <SPLIT distance="225" swimtime="00:03:32.76" />
                    <SPLIT distance="250" swimtime="00:04:00.47" />
                    <SPLIT distance="275" swimtime="00:04:28.20" />
                    <SPLIT distance="300" swimtime="00:04:56.39" />
                    <SPLIT distance="325" swimtime="00:05:19.39" />
                    <SPLIT distance="350" swimtime="00:05:41.27" />
                    <SPLIT distance="375" swimtime="00:06:03.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="311" swimtime="00:01:20.54" resultid="108528" heatid="110795" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.39" />
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="75" swimtime="00:00:58.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="108494" lastname.en="Kuliś">
              <RESULTS>
                <RESULT eventid="98777" points="501" reactiontime="+84" swimtime="00:00:29.25" resultid="108495" heatid="110592" lane="2" entrytime="00:00:29.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="394" reactiontime="+65" swimtime="00:00:34.99" resultid="108496" heatid="110649" lane="8" entrytime="00:00:38.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="427" swimtime="00:01:15.21" resultid="108497" heatid="110695" lane="9" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.08" />
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="75" swimtime="00:00:56.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="432" swimtime="00:00:32.25" resultid="108498" heatid="110740" lane="0" entrytime="00:00:32.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="372" reactiontime="+78" swimtime="00:01:16.50" resultid="108499" heatid="110756" lane="1" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.11" />
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="75" swimtime="00:00:56.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="508" swimtime="00:00:36.09" resultid="108500" heatid="110823" lane="6" entrytime="00:00:36.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-03" firstname="Marcin" gender="M" lastname="Wyżga" nation="POL" athleteid="108552">
              <RESULTS>
                <RESULT eventid="98798" points="374" reactiontime="+86" swimtime="00:00:28.10" resultid="108553" heatid="110605" lane="1" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="263" reactiontime="+69" swimtime="00:00:34.68" resultid="108554" heatid="110657" lane="8" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="353" reactiontime="+77" swimtime="00:00:30.82" resultid="108555" heatid="110746" lane="5" entrytime="00:00:31.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="336" reactiontime="+81" swimtime="00:00:36.31" resultid="108556" heatid="110829" lane="7" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-24" firstname="Bogusław" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="108574">
              <RESULTS>
                <RESULT eventid="98798" points="53" reactiontime="+104" swimtime="00:00:53.65" resultid="108575" heatid="110595" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="37" reactiontime="+88" swimtime="00:01:06.48" resultid="108576" heatid="110651" lane="7">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="43" reactiontime="+106" swimtime="00:02:07.65" resultid="108577" heatid="110677" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.54" />
                    <SPLIT distance="50" swimtime="00:00:56.45" />
                    <SPLIT distance="75" swimtime="00:01:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="45" reactiontime="+104" swimtime="00:02:35.38" resultid="108578" heatid="110726" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.16" />
                    <SPLIT distance="50" swimtime="00:01:13.88" />
                    <SPLIT distance="75" swimtime="00:01:54.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="42" reactiontime="+123" swimtime="00:04:44.39" resultid="108579" heatid="110769" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.72" />
                    <SPLIT distance="50" swimtime="00:01:00.30" />
                    <SPLIT distance="75" swimtime="00:01:35.28" />
                    <SPLIT distance="100" swimtime="00:02:13.63" />
                    <SPLIT distance="125" swimtime="00:02:51.56" />
                    <SPLIT distance="150" swimtime="00:03:30.33" />
                    <SPLIT distance="175" swimtime="00:04:08.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="35" reactiontime="+101" swimtime="00:05:20.30" resultid="108580" heatid="110810" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.78" />
                    <SPLIT distance="50" swimtime="00:01:14.54" />
                    <SPLIT distance="75" swimtime="00:01:53.63" />
                    <SPLIT distance="100" swimtime="00:02:35.98" />
                    <SPLIT distance="125" swimtime="00:03:18.08" />
                    <SPLIT distance="150" swimtime="00:04:00.45" />
                    <SPLIT distance="175" swimtime="00:04:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="50" reactiontime="+112" swimtime="00:01:08.23" resultid="108581" heatid="110824" lane="8">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-16" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="108582">
              <RESULTS>
                <RESULT eventid="98798" points="73" reactiontime="+69" swimtime="00:00:48.47" resultid="108583" heatid="110595" lane="4" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="28" reactiontime="+120" swimtime="00:05:58.31" resultid="108584" heatid="110619" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.71" />
                    <SPLIT distance="50" swimtime="00:01:27.05" />
                    <SPLIT distance="75" swimtime="00:02:10.59" />
                    <SPLIT distance="100" swimtime="00:02:57.15" />
                    <SPLIT distance="125" swimtime="00:03:55.93" />
                    <SPLIT distance="150" swimtime="00:04:53.68" />
                    <SPLIT distance="175" swimtime="00:05:24.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="57" reactiontime="+113" swimtime="00:01:56.30" resultid="108585" heatid="110678" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.18" />
                    <SPLIT distance="50" swimtime="00:00:51.74" />
                    <SPLIT distance="75" swimtime="00:01:24.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="30" reactiontime="+112" swimtime="00:02:41.33" resultid="108586" heatid="110696" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.68" />
                    <SPLIT distance="50" swimtime="00:01:15.00" />
                    <SPLIT distance="75" swimtime="00:02:14.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="14" swimtime="00:01:30.21" resultid="108587" heatid="110742" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="51" swimtime="00:04:27.20" resultid="108588" heatid="110769" lane="6" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.71" />
                    <SPLIT distance="50" swimtime="00:00:56.27" />
                    <SPLIT distance="75" swimtime="00:01:28.55" />
                    <SPLIT distance="100" swimtime="00:02:04.61" />
                    <SPLIT distance="125" swimtime="00:02:40.34" />
                    <SPLIT distance="150" swimtime="00:03:17.02" />
                    <SPLIT distance="175" swimtime="00:03:53.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="108589" heatid="110810" lane="4" entrytime="00:05:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="108529">
              <RESULTS>
                <RESULT eventid="98798" points="210" reactiontime="+118" swimtime="00:00:34.07" resultid="108530" heatid="110601" lane="1" entrytime="00:00:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="124" reactiontime="+125" swimtime="00:03:39.72" resultid="108531" heatid="110620" lane="4" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.53" />
                    <SPLIT distance="50" swimtime="00:00:47.67" />
                    <SPLIT distance="75" swimtime="00:01:17.83" />
                    <SPLIT distance="100" swimtime="00:01:46.80" />
                    <SPLIT distance="125" swimtime="00:02:21.10" />
                    <SPLIT distance="150" swimtime="00:02:52.22" />
                    <SPLIT distance="175" swimtime="00:03:18.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="211" reactiontime="+107" swimtime="00:01:15.39" resultid="108532" heatid="110681" lane="5" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.92" />
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="75" swimtime="00:00:56.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="63" reactiontime="+140" swimtime="00:04:32.63" resultid="108533" heatid="110710" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.69" />
                    <SPLIT distance="50" swimtime="00:01:01.71" />
                    <SPLIT distance="75" swimtime="00:01:38.11" />
                    <SPLIT distance="100" swimtime="00:02:12.27" />
                    <SPLIT distance="125" swimtime="00:02:46.56" />
                    <SPLIT distance="150" swimtime="00:03:21.42" />
                    <SPLIT distance="175" swimtime="00:03:57.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="165" reactiontime="+137" swimtime="00:03:00.82" resultid="108534" heatid="110771" lane="3" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.58" />
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="75" swimtime="00:01:03.48" />
                    <SPLIT distance="100" swimtime="00:01:25.97" />
                    <SPLIT distance="125" swimtime="00:01:49.44" />
                    <SPLIT distance="150" swimtime="00:02:12.79" />
                    <SPLIT distance="175" swimtime="00:02:37.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="99" reactiontime="+153" swimtime="00:08:27.79" resultid="108535" heatid="110788" lane="3" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.42" />
                    <SPLIT distance="50" swimtime="00:00:56.12" />
                    <SPLIT distance="75" swimtime="00:01:30.05" />
                    <SPLIT distance="100" swimtime="00:02:02.68" />
                    <SPLIT distance="125" swimtime="00:02:37.00" />
                    <SPLIT distance="150" swimtime="00:03:13.02" />
                    <SPLIT distance="175" swimtime="00:03:48.91" />
                    <SPLIT distance="200" swimtime="00:04:26.15" />
                    <SPLIT distance="225" swimtime="00:04:59.68" />
                    <SPLIT distance="250" swimtime="00:05:35.45" />
                    <SPLIT distance="275" swimtime="00:06:11.38" />
                    <SPLIT distance="300" swimtime="00:06:47.63" />
                    <SPLIT distance="325" swimtime="00:07:14.49" />
                    <SPLIT distance="350" swimtime="00:07:40.02" />
                    <SPLIT distance="375" swimtime="00:08:03.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="86" swimtime="00:01:49.60" resultid="108536" heatid="110799" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.92" />
                    <SPLIT distance="50" swimtime="00:00:49.97" />
                    <SPLIT distance="75" swimtime="00:01:18.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="142" reactiontime="+141" swimtime="00:06:46.76" resultid="108537" heatid="110850" lane="4" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.96" />
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                    <SPLIT distance="75" swimtime="00:01:13.43" />
                    <SPLIT distance="100" swimtime="00:01:39.97" />
                    <SPLIT distance="125" swimtime="00:02:06.32" />
                    <SPLIT distance="150" swimtime="00:02:32.97" />
                    <SPLIT distance="175" swimtime="00:02:58.66" />
                    <SPLIT distance="200" swimtime="00:03:24.39" />
                    <SPLIT distance="225" swimtime="00:04:40.99" />
                    <SPLIT distance="250" swimtime="00:04:16.24" />
                    <SPLIT distance="300" swimtime="00:05:07.14" />
                    <SPLIT distance="325" swimtime="00:05:32.31" />
                    <SPLIT distance="350" swimtime="00:05:58.25" />
                    <SPLIT distance="375" swimtime="00:06:23.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="Frączek" nation="POL" athleteid="108563">
              <RESULTS>
                <RESULT eventid="98777" points="527" reactiontime="+81" swimtime="00:00:28.76" resultid="108564" heatid="110593" lane="4" entrytime="00:00:26.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="337" reactiontime="+73" swimtime="00:00:36.88" resultid="108565" heatid="110649" lane="2" entrytime="00:00:37.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="463" swimtime="00:01:05.79" resultid="108566" heatid="110676" lane="0" entrytime="00:01:05.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.88" />
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="75" swimtime="00:00:47.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="421" reactiontime="+85" swimtime="00:00:32.51" resultid="108567" heatid="110739" lane="4" entrytime="00:00:32.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="108568" heatid="110767" lane="3" entrytime="00:02:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-05" firstname="Mateo" gender="M" lastname="Morlupi" nation="POL" athleteid="108590">
              <RESULTS>
                <RESULT eventid="98798" points="252" swimtime="00:00:32.07" resultid="108591" heatid="110601" lane="9" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="197" reactiontime="+89" swimtime="00:01:17.22" resultid="108592" heatid="110681" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.03" />
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="242" reactiontime="+86" swimtime="00:01:29.18" resultid="108593" heatid="110729" lane="4" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.90" />
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                    <SPLIT distance="75" swimtime="00:01:04.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="269" swimtime="00:00:39.09" resultid="108594" heatid="110829" lane="0" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-30" firstname="Piotr" gender="M" lastname="Łysiak" nation="POL" athleteid="108557">
              <RESULTS>
                <RESULT eventid="98798" points="339" reactiontime="+69" swimtime="00:00:29.04" resultid="108558" heatid="110606" lane="6" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="266" reactiontime="+63" swimtime="00:00:34.52" resultid="108559" heatid="110656" lane="6" entrytime="00:00:34.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="324" swimtime="00:02:55.33" resultid="108560" heatid="110669" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.85" />
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="75" swimtime="00:01:01.85" />
                    <SPLIT distance="100" swimtime="00:01:23.91" />
                    <SPLIT distance="125" swimtime="00:01:45.82" />
                    <SPLIT distance="150" swimtime="00:02:08.72" />
                    <SPLIT distance="175" swimtime="00:02:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="340" reactiontime="+92" swimtime="00:01:19.67" resultid="108561" heatid="110732" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.82" />
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="75" swimtime="00:00:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="108562" heatid="110827" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-26" firstname="Józef" gender="M" lastname="Śmigielski" nation="POL" athleteid="108518">
              <RESULTS>
                <RESULT eventid="98798" points="75" reactiontime="+113" swimtime="00:00:47.91" resultid="108519" heatid="110595" lane="5" entrytime="00:00:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="43" reactiontime="+112" swimtime="00:01:03.12" resultid="108520" heatid="110652" lane="0" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="108521" heatid="110678" lane="6" entrytime="00:01:57.00" />
                <RESULT eventid="99186" points="55" reactiontime="+124" swimtime="00:02:08.51" resultid="108522" heatid="110758" lane="0" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.48" />
                    <SPLIT distance="50" swimtime="00:01:01.37" />
                    <SPLIT distance="75" swimtime="00:01:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="60" reactiontime="+99" swimtime="00:04:29.81" resultid="108523" heatid="110811" lane="8" entrytime="00:04:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.18" />
                    <SPLIT distance="50" swimtime="00:01:02.47" />
                    <SPLIT distance="75" swimtime="00:01:35.83" />
                    <SPLIT distance="100" swimtime="00:02:11.64" />
                    <SPLIT distance="125" swimtime="00:02:45.88" />
                    <SPLIT distance="150" swimtime="00:03:21.43" />
                    <SPLIT distance="175" swimtime="00:03:56.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="108501">
              <RESULTS>
                <RESULT eventid="98777" points="321" swimtime="00:00:33.91" resultid="108502" heatid="110590" lane="9" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="267" swimtime="00:12:23.86" resultid="108503" heatid="110634" lane="9" entrytime="00:12:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.90" />
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="75" swimtime="00:01:01.57" />
                    <SPLIT distance="100" swimtime="00:01:24.18" />
                    <SPLIT distance="125" swimtime="00:01:46.97" />
                    <SPLIT distance="150" swimtime="00:02:10.69" />
                    <SPLIT distance="175" swimtime="00:02:34.16" />
                    <SPLIT distance="200" swimtime="00:02:57.54" />
                    <SPLIT distance="225" swimtime="00:03:21.23" />
                    <SPLIT distance="250" swimtime="00:03:44.86" />
                    <SPLIT distance="275" swimtime="00:04:08.59" />
                    <SPLIT distance="300" swimtime="00:04:32.25" />
                    <SPLIT distance="325" swimtime="00:04:56.43" />
                    <SPLIT distance="350" swimtime="00:05:20.33" />
                    <SPLIT distance="375" swimtime="00:05:44.72" />
                    <SPLIT distance="400" swimtime="00:06:08.64" />
                    <SPLIT distance="425" swimtime="00:06:32.40" />
                    <SPLIT distance="450" swimtime="00:06:56.30" />
                    <SPLIT distance="475" swimtime="00:07:19.90" />
                    <SPLIT distance="500" swimtime="00:07:44.11" />
                    <SPLIT distance="525" swimtime="00:08:07.82" />
                    <SPLIT distance="550" swimtime="00:08:31.61" />
                    <SPLIT distance="575" swimtime="00:08:55.62" />
                    <SPLIT distance="600" swimtime="00:09:19.52" />
                    <SPLIT distance="625" swimtime="00:09:43.00" />
                    <SPLIT distance="650" swimtime="00:10:06.53" />
                    <SPLIT distance="675" swimtime="00:10:29.59" />
                    <SPLIT distance="700" swimtime="00:10:53.08" />
                    <SPLIT distance="725" swimtime="00:11:16.66" />
                    <SPLIT distance="750" swimtime="00:11:40.07" />
                    <SPLIT distance="775" swimtime="00:12:02.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="314" reactiontime="+81" swimtime="00:01:14.87" resultid="108504" heatid="110674" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.23" />
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="75" swimtime="00:00:55.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" status="DNS" swimtime="00:00:00.00" resultid="108505" heatid="110708" lane="1" entrytime="00:03:25.00" />
                <RESULT eventid="99154" points="257" swimtime="00:00:38.33" resultid="108506" heatid="110738" lane="9" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="276" swimtime="00:02:50.04" resultid="108507" heatid="110767" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="75" swimtime="00:01:00.10" />
                    <SPLIT distance="100" swimtime="00:01:21.46" />
                    <SPLIT distance="125" swimtime="00:01:43.86" />
                    <SPLIT distance="150" swimtime="00:02:06.41" />
                    <SPLIT distance="175" swimtime="00:02:29.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="228" swimtime="00:01:29.33" resultid="108508" heatid="110794" lane="4" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.84" />
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                    <SPLIT distance="75" swimtime="00:01:03.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="277" swimtime="00:05:59.53" resultid="108509" heatid="110840" lane="9" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.66" />
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                    <SPLIT distance="75" swimtime="00:01:01.47" />
                    <SPLIT distance="100" swimtime="00:01:23.78" />
                    <SPLIT distance="125" swimtime="00:01:46.39" />
                    <SPLIT distance="150" swimtime="00:02:09.72" />
                    <SPLIT distance="175" swimtime="00:02:32.81" />
                    <SPLIT distance="200" swimtime="00:02:56.06" />
                    <SPLIT distance="225" swimtime="00:03:18.74" />
                    <SPLIT distance="250" swimtime="00:03:41.69" />
                    <SPLIT distance="275" swimtime="00:04:04.74" />
                    <SPLIT distance="300" swimtime="00:04:28.07" />
                    <SPLIT distance="325" swimtime="00:04:51.34" />
                    <SPLIT distance="350" swimtime="00:05:14.95" />
                    <SPLIT distance="375" swimtime="00:05:37.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="108547">
              <RESULTS>
                <RESULT eventid="106294" points="249" reactiontime="+86" swimtime="00:00:40.78" resultid="108548" heatid="110648" lane="2" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="226" reactiontime="+107" swimtime="00:01:33.00" resultid="108549" heatid="110692" lane="1" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.18" />
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                    <SPLIT distance="75" swimtime="00:01:12.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="270" reactiontime="+95" swimtime="00:00:37.72" resultid="108550" heatid="110737" lane="4" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="216" reactiontime="+88" swimtime="00:03:18.60" resultid="108551" heatid="110807" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.51" />
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="75" swimtime="00:01:11.40" />
                    <SPLIT distance="100" swimtime="00:01:37.23" />
                    <SPLIT distance="125" swimtime="00:02:04.00" />
                    <SPLIT distance="150" swimtime="00:02:30.41" />
                    <SPLIT distance="175" swimtime="00:02:55.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-08" firstname="Tomasz" gender="M" lastname="Czerniecki" nation="POL" athleteid="108569">
              <RESULTS>
                <RESULT eventid="98798" points="496" reactiontime="+69" swimtime="00:00:25.59" resultid="108570" heatid="110611" lane="5" entrytime="00:00:25.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="496" reactiontime="+79" swimtime="00:00:56.76" resultid="108571" heatid="110677" lane="4">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.95" />
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="75" swimtime="00:00:41.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="424" swimtime="00:01:07.40" resultid="108572" heatid="110705" lane="9" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="75" swimtime="00:00:51.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="394" reactiontime="+78" swimtime="00:00:29.73" resultid="108573" heatid="110748" lane="5" entrytime="00:00:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="108510">
              <RESULTS>
                <RESULT eventid="98798" points="100" reactiontime="+115" swimtime="00:00:43.62" resultid="108511" heatid="110596" lane="0" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="97" reactiontime="+123" swimtime="00:30:43.76" resultid="108512" heatid="110643" lane="1" entrytime="00:32:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.06" />
                    <SPLIT distance="50" swimtime="00:00:57.46" />
                    <SPLIT distance="75" swimtime="00:01:27.57" />
                    <SPLIT distance="100" swimtime="00:01:58.18" />
                    <SPLIT distance="125" swimtime="00:02:29.34" />
                    <SPLIT distance="150" swimtime="00:03:01.46" />
                    <SPLIT distance="175" swimtime="00:03:32.40" />
                    <SPLIT distance="200" swimtime="00:04:03.73" />
                    <SPLIT distance="225" swimtime="00:04:34.52" />
                    <SPLIT distance="250" swimtime="00:05:06.24" />
                    <SPLIT distance="275" swimtime="00:05:36.71" />
                    <SPLIT distance="300" swimtime="00:06:07.53" />
                    <SPLIT distance="325" swimtime="00:06:38.21" />
                    <SPLIT distance="350" swimtime="00:07:09.34" />
                    <SPLIT distance="375" swimtime="00:07:40.55" />
                    <SPLIT distance="400" swimtime="00:08:11.97" />
                    <SPLIT distance="425" swimtime="00:08:42.93" />
                    <SPLIT distance="450" swimtime="00:09:14.70" />
                    <SPLIT distance="475" swimtime="00:09:45.26" />
                    <SPLIT distance="500" swimtime="00:10:16.72" />
                    <SPLIT distance="525" swimtime="00:10:47.71" />
                    <SPLIT distance="550" swimtime="00:11:18.76" />
                    <SPLIT distance="575" swimtime="00:11:49.10" />
                    <SPLIT distance="600" swimtime="00:12:19.54" />
                    <SPLIT distance="625" swimtime="00:12:49.85" />
                    <SPLIT distance="650" swimtime="00:13:21.42" />
                    <SPLIT distance="675" swimtime="00:13:51.92" />
                    <SPLIT distance="700" swimtime="00:14:23.07" />
                    <SPLIT distance="725" swimtime="00:14:54.27" />
                    <SPLIT distance="750" swimtime="00:15:25.74" />
                    <SPLIT distance="775" swimtime="00:15:56.19" />
                    <SPLIT distance="800" swimtime="00:16:27.94" />
                    <SPLIT distance="825" swimtime="00:16:58.35" />
                    <SPLIT distance="850" swimtime="00:17:29.48" />
                    <SPLIT distance="875" swimtime="00:18:00.13" />
                    <SPLIT distance="900" swimtime="00:18:30.35" />
                    <SPLIT distance="925" swimtime="00:19:01.33" />
                    <SPLIT distance="950" swimtime="00:19:32.43" />
                    <SPLIT distance="975" swimtime="00:20:03.04" />
                    <SPLIT distance="1000" swimtime="00:20:34.78" />
                    <SPLIT distance="1025" swimtime="00:21:05.62" />
                    <SPLIT distance="1050" swimtime="00:21:37.58" />
                    <SPLIT distance="1075" swimtime="00:22:07.96" />
                    <SPLIT distance="1100" swimtime="00:22:38.63" />
                    <SPLIT distance="1125" swimtime="00:23:08.79" />
                    <SPLIT distance="1150" swimtime="00:23:40.51" />
                    <SPLIT distance="1175" swimtime="00:24:10.98" />
                    <SPLIT distance="1200" swimtime="00:24:41.92" />
                    <SPLIT distance="1225" swimtime="00:25:12.24" />
                    <SPLIT distance="1250" swimtime="00:25:43.18" />
                    <SPLIT distance="1275" swimtime="00:26:13.08" />
                    <SPLIT distance="1300" swimtime="00:26:44.04" />
                    <SPLIT distance="1325" swimtime="00:27:14.49" />
                    <SPLIT distance="1350" swimtime="00:27:45.44" />
                    <SPLIT distance="1375" swimtime="00:28:14.71" />
                    <SPLIT distance="1400" swimtime="00:28:43.97" />
                    <SPLIT distance="1425" swimtime="00:29:14.22" />
                    <SPLIT distance="1450" swimtime="00:29:45.59" />
                    <SPLIT distance="1475" swimtime="00:30:15.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="99" reactiontime="+110" swimtime="00:01:36.95" resultid="108513" heatid="110679" lane="8" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.20" />
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                    <SPLIT distance="75" swimtime="00:01:10.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="67" reactiontime="+125" swimtime="00:02:16.75" resultid="108514" heatid="110727" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.87" />
                    <SPLIT distance="50" swimtime="00:01:03.78" />
                    <SPLIT distance="75" swimtime="00:01:39.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="88" reactiontime="+119" swimtime="00:03:42.81" resultid="108515" heatid="110769" lane="3" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.77" />
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                    <SPLIT distance="75" swimtime="00:01:19.68" />
                    <SPLIT distance="100" swimtime="00:01:47.92" />
                    <SPLIT distance="125" swimtime="00:02:16.99" />
                    <SPLIT distance="150" swimtime="00:02:45.71" />
                    <SPLIT distance="175" swimtime="00:03:15.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="68" reactiontime="+119" swimtime="00:01:01.73" resultid="108516" heatid="110824" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="84" swimtime="00:08:04.09" resultid="108517" heatid="110851" lane="0" entrytime="00:07:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.61" />
                    <SPLIT distance="50" swimtime="00:00:57.49" />
                    <SPLIT distance="75" swimtime="00:01:27.28" />
                    <SPLIT distance="100" swimtime="00:01:58.06" />
                    <SPLIT distance="125" swimtime="00:02:30.22" />
                    <SPLIT distance="150" swimtime="00:03:01.58" />
                    <SPLIT distance="175" swimtime="00:03:32.85" />
                    <SPLIT distance="200" swimtime="00:04:04.30" />
                    <SPLIT distance="225" swimtime="00:04:35.08" />
                    <SPLIT distance="250" swimtime="00:05:06.02" />
                    <SPLIT distance="275" swimtime="00:05:37.07" />
                    <SPLIT distance="300" swimtime="00:06:07.29" />
                    <SPLIT distance="325" swimtime="00:06:38.23" />
                    <SPLIT distance="350" swimtime="00:07:08.87" />
                    <SPLIT distance="375" swimtime="00:07:37.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="108538">
              <RESULTS>
                <RESULT eventid="98777" points="47" reactiontime="+102" swimtime="00:01:04.33" resultid="108539" heatid="110586" lane="7" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="43" reactiontime="+106" swimtime="00:05:46.50" resultid="108540" heatid="110614" lane="7" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:37.26" />
                    <SPLIT distance="50" swimtime="00:01:21.37" />
                    <SPLIT distance="75" swimtime="00:02:09.23" />
                    <SPLIT distance="100" swimtime="00:02:58.88" />
                    <SPLIT distance="125" swimtime="00:03:43.76" />
                    <SPLIT distance="150" swimtime="00:04:28.73" />
                    <SPLIT distance="175" swimtime="00:05:07.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="47" swimtime="00:02:20.58" resultid="108541" heatid="110672" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.14" />
                    <SPLIT distance="50" swimtime="00:01:05.94" />
                    <SPLIT distance="75" swimtime="00:01:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="45" reactiontime="+113" swimtime="00:02:38.78" resultid="108542" heatid="110690" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.94" />
                    <SPLIT distance="50" swimtime="00:01:18.69" />
                    <SPLIT distance="75" swimtime="00:02:01.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="62" reactiontime="+121" swimtime="00:02:37.19" resultid="108543" heatid="110721" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.11" />
                    <SPLIT distance="50" swimtime="00:01:12.94" />
                    <SPLIT distance="75" swimtime="00:01:55.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="29" swimtime="00:01:18.82" resultid="108544" heatid="110736" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="25" swimtime="00:03:04.92" resultid="108545" heatid="110793" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:39.47" />
                    <SPLIT distance="50" swimtime="00:01:26.23" />
                    <SPLIT distance="75" swimtime="00:02:15.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="82" swimtime="00:01:06.19" resultid="108546" heatid="110818" lane="0" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Masters Korona Kraków C" number="1">
              <RESULTS>
                <RESULT eventid="99059" status="DNS" swimtime="00:00:00.00" resultid="108603" heatid="110718" lane="2" entrytime="00:02:07.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108557" number="1" />
                    <RELAYPOSITION athleteid="108590" number="2" />
                    <RELAYPOSITION athleteid="108552" number="3" />
                    <RELAYPOSITION athleteid="108569" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" name="Masters Korona Kraków F" number="1">
              <RESULTS>
                <RESULT comment="S4/ III ZMIANA" eventid="99059" reactiontime="+101" status="DSQ" swimtime="00:00:00.00" resultid="108595" heatid="110716" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.17" />
                    <SPLIT distance="50" swimtime="00:01:00.54" />
                    <SPLIT distance="75" swimtime="00:01:29.03" />
                    <SPLIT distance="100" swimtime="00:02:01.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108518" number="1" reactiontime="+101" status="DSQ" />
                    <RELAYPOSITION athleteid="108510" number="2" reactiontime="+54" status="DSQ" />
                    <RELAYPOSITION athleteid="108529" number="3" reactiontime="-69" status="DSQ" />
                    <RELAYPOSITION athleteid="108582" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="101" reactiontime="+134" swimtime="00:02:56.82" resultid="108596" heatid="110781" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.67" />
                    <SPLIT distance="50" swimtime="00:00:51.09" />
                    <SPLIT distance="75" swimtime="00:01:13.19" />
                    <SPLIT distance="100" swimtime="00:01:39.44" />
                    <SPLIT distance="125" swimtime="00:01:56.46" />
                    <SPLIT distance="150" swimtime="00:02:04.85" />
                    <SPLIT distance="175" swimtime="00:02:33.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108518" number="1" reactiontime="+134" />
                    <RELAYPOSITION athleteid="108582" number="2" reactiontime="+96" />
                    <RELAYPOSITION athleteid="108529" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="108510" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Masters Korona Kraków D" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="386" reactiontime="+58" swimtime="00:02:22.80" resultid="108599" heatid="110715" lane="6" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.67" />
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="75" swimtime="00:00:53.58" />
                    <SPLIT distance="100" swimtime="00:01:12.99" />
                    <SPLIT distance="125" swimtime="00:01:29.51" />
                    <SPLIT distance="150" swimtime="00:01:48.54" />
                    <SPLIT distance="175" swimtime="00:02:05.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108501" number="1" reactiontime="+58" />
                    <RELAYPOSITION athleteid="108494" number="2" />
                    <RELAYPOSITION athleteid="108524" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="108563" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99234" points="420" swimtime="00:02:05.84" resultid="108600" heatid="110780" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.37" />
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                    <SPLIT distance="75" swimtime="00:00:45.89" />
                    <SPLIT distance="100" swimtime="00:01:03.09" />
                    <SPLIT distance="125" swimtime="00:01:20.07" />
                    <SPLIT distance="150" swimtime="00:01:37.53" />
                    <SPLIT distance="175" swimtime="00:01:51.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108494" number="1" />
                    <RELAYPOSITION athleteid="108524" number="2" />
                    <RELAYPOSITION athleteid="108501" number="3" />
                    <RELAYPOSITION athleteid="108563" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Masters Korona Kraków " number="2">
              <RESULTS>
                <RESULT eventid="99441" points="282" reactiontime="+79" swimtime="00:02:17.95" resultid="108602" heatid="110838" lane="1" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.21" />
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="75" swimtime="00:00:51.36" />
                    <SPLIT distance="100" swimtime="00:01:11.18" />
                    <SPLIT distance="125" swimtime="00:01:26.49" />
                    <SPLIT distance="150" swimtime="00:01:44.19" />
                    <SPLIT distance="175" swimtime="00:02:00.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108557" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="108494" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="108563" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="108529" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Masters Korona Kraków C" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="413" reactiontime="+73" swimtime="00:01:50.87" resultid="108601" heatid="110632" lane="8" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                    <SPLIT distance="75" swimtime="00:00:42.30" />
                    <SPLIT distance="100" swimtime="00:00:56.53" />
                    <SPLIT distance="125" swimtime="00:01:10.41" />
                    <SPLIT distance="150" swimtime="00:01:25.19" />
                    <SPLIT distance="175" swimtime="00:01:37.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108494" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="108557" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="108563" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="108569" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Masters Korona Kraków D" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="250" reactiontime="+67" swimtime="00:02:11.11" resultid="108597" heatid="110630" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.07" />
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="75" swimtime="00:00:45.80" />
                    <SPLIT distance="100" swimtime="00:01:03.67" />
                    <SPLIT distance="125" swimtime="00:01:19.83" />
                    <SPLIT distance="150" swimtime="00:01:37.75" />
                    <SPLIT distance="175" swimtime="00:01:54.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108552" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="108501" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="108524" number="3" reactiontime="+15" />
                    <RELAYPOSITION athleteid="108529" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="108598" heatid="110836" lane="9" entrytime="00:03:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108501" number="1" />
                    <RELAYPOSITION athleteid="108590" number="2" />
                    <RELAYPOSITION athleteid="108524" number="3" />
                    <RELAYPOSITION athleteid="108529" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="106946" name="Masters Swim">
          <CONTACT email="basen@wladcywody.pl" name="Wereszczyński" phone="723897862" street="Kłodzka" zip="55-040" />
          <ATHLETES>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="106956">
              <RESULTS>
                <RESULT eventid="98777" points="241" reactiontime="+71" swimtime="00:00:37.34" resultid="106957" heatid="110588" lane="5" entrytime="00:00:37.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="147" reactiontime="+93" swimtime="00:03:50.38" resultid="106958" heatid="110615" lane="0" entrytime="00:03:47.93">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.09" />
                    <SPLIT distance="50" swimtime="00:00:54.92" />
                    <SPLIT distance="75" swimtime="00:01:25.39" />
                    <SPLIT distance="100" swimtime="00:01:56.42" />
                    <SPLIT distance="125" swimtime="00:02:26.74" />
                    <SPLIT distance="150" swimtime="00:02:57.87" />
                    <SPLIT distance="175" swimtime="00:03:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="122" reactiontime="+102" swimtime="00:00:51.72" resultid="106959" heatid="110647" lane="2" entrytime="00:00:48.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="201" reactiontime="+84" swimtime="00:01:26.83" resultid="106960" heatid="110673" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.95" />
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                    <SPLIT distance="75" swimtime="00:01:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="233" swimtime="00:01:41.28" resultid="106961" heatid="110722" lane="6" entrytime="00:01:43.47">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.33" />
                    <SPLIT distance="50" swimtime="00:00:48.18" />
                    <SPLIT distance="75" swimtime="00:01:15.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="106962" heatid="110765" lane="9" entrytime="00:03:25.31" />
                <RESULT eventid="99409" points="254" reactiontime="+63" swimtime="00:00:45.44" resultid="106963" heatid="110820" lane="7" entrytime="00:00:45.74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-13" firstname="Maciej" gender="M" lastname="Dąbrowski" nation="POL" athleteid="106947">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="106948" heatid="110604" lane="3" entrytime="00:00:29.50" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="106949" heatid="110624" lane="1" entrytime="00:02:47.00" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="106950" heatid="110656" lane="2" entrytime="00:00:34.50" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="106951" heatid="110701" lane="4" entrytime="00:01:14.50" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="106952" heatid="110745" lane="0" entrytime="00:00:33.50" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="106953" heatid="110761" lane="0" entrytime="00:01:17.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="106954" heatid="110801" lane="8" entrytime="00:01:18.00" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="106955" heatid="110814" lane="0" entrytime="00:02:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="107702" name="Masters Team Biała Podlaska">
          <CONTACT city="Biała Podlaska" email="wilhelmg@poczta.onet.pl" name="Gromisz" zip="21-500" />
          <ATHLETES>
            <ATHLETE birthdate="1981-11-29" firstname="Iga" gender="F" lastname="Olszanowska" nation="POL" athleteid="107703">
              <RESULTS>
                <RESULT eventid="98777" points="475" reactiontime="+99" swimtime="00:00:29.78" resultid="107704" heatid="110593" lane="0" entrytime="00:00:28.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="389" reactiontime="+79" swimtime="00:02:46.81" resultid="107705" heatid="110618" lane="0" entrytime="00:02:44.31">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.52" />
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="75" swimtime="00:00:56.45" />
                    <SPLIT distance="100" swimtime="00:01:18.72" />
                    <SPLIT distance="125" swimtime="00:01:41.72" />
                    <SPLIT distance="150" swimtime="00:02:06.46" />
                    <SPLIT distance="175" swimtime="00:02:27.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="472" reactiontime="+90" swimtime="00:01:05.38" resultid="107706" heatid="110676" lane="8" entrytime="00:01:05.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.07" />
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="75" swimtime="00:00:48.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="416" reactiontime="+86" swimtime="00:01:15.89" resultid="107707" heatid="110695" lane="2" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.34" />
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="75" swimtime="00:00:57.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="464" swimtime="00:00:31.47" resultid="107708" heatid="110740" lane="6" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="399" reactiontime="+91" swimtime="00:02:30.45" resultid="107709" heatid="110768" lane="8" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.99" />
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="75" swimtime="00:00:52.48" />
                    <SPLIT distance="100" swimtime="00:01:11.89" />
                    <SPLIT distance="125" swimtime="00:01:31.51" />
                    <SPLIT distance="150" swimtime="00:01:51.55" />
                    <SPLIT distance="175" swimtime="00:02:11.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="401" reactiontime="+95" swimtime="00:01:14.04" resultid="107710" heatid="110796" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.51" />
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="75" swimtime="00:00:53.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="415" reactiontime="+96" swimtime="00:00:38.59" resultid="107711" heatid="110822" lane="8" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-12-27" firstname="Renata" gender="F" lastname="Kasprowicz" nation="POL" athleteid="107712">
              <RESULTS>
                <RESULT eventid="98777" points="448" reactiontime="+80" swimtime="00:00:30.35" resultid="107713" heatid="110592" lane="3" entrytime="00:00:29.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="355" reactiontime="+61" swimtime="00:03:09.94" resultid="107714" heatid="110664" lane="7" entrytime="00:03:00.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.05" />
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="75" swimtime="00:01:03.36" />
                    <SPLIT distance="100" swimtime="00:01:27.16" />
                    <SPLIT distance="125" swimtime="00:01:51.78" />
                    <SPLIT distance="150" swimtime="00:02:17.67" />
                    <SPLIT distance="175" swimtime="00:02:43.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="364" reactiontime="+78" swimtime="00:01:19.33" resultid="107715" heatid="110694" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.94" />
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="75" swimtime="00:01:00.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="396" swimtime="00:01:24.88" resultid="107716" heatid="110725" lane="0" entrytime="00:01:23.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.64" />
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="75" swimtime="00:01:01.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="384" reactiontime="+78" swimtime="00:00:33.54" resultid="107717" heatid="110739" lane="5" entrytime="00:00:32.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="418" reactiontime="+80" swimtime="00:00:38.51" resultid="107718" heatid="110822" lane="4" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-15" firstname="Michal" gender="M" lastname="Jagiełło" nation="POL" athleteid="107719">
              <RESULTS>
                <RESULT eventid="98798" points="492" reactiontime="+91" swimtime="00:00:25.66" resultid="107720" heatid="110613" lane="1" entrytime="00:00:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="544" reactiontime="+62" swimtime="00:00:55.03" resultid="107721" heatid="110689" lane="6" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.03" />
                    <SPLIT distance="50" swimtime="00:00:25.89" />
                    <SPLIT distance="75" swimtime="00:00:40.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="505" reactiontime="+78" swimtime="00:00:27.36" resultid="107722" heatid="110750" lane="3" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-03" firstname="Wilhelm" gender="M" lastname="Gromisz" nation="POL" athleteid="107723">
              <RESULTS>
                <RESULT eventid="98798" points="465" swimtime="00:00:26.14" resultid="107724" heatid="110612" lane="9" entrytime="00:00:25.35">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="492" reactiontime="+76" swimtime="00:00:28.14" resultid="107725" heatid="110660" lane="3" entrytime="00:00:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="479" reactiontime="+100" swimtime="00:00:57.41" resultid="107726" heatid="110688" lane="2" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.38" />
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                    <SPLIT distance="75" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="510" reactiontime="+104" swimtime="00:00:27.28" resultid="107727" heatid="110751" lane="8" entrytime="00:00:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="482" reactiontime="+77" swimtime="00:01:02.37" resultid="107728" heatid="110763" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.54" />
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                    <SPLIT distance="75" swimtime="00:00:46.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="509" reactiontime="+108" swimtime="00:01:00.66" resultid="107729" heatid="110805" lane="1" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                    <SPLIT distance="75" swimtime="00:00:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="414" reactiontime="+84" swimtime="00:02:21.65" resultid="107730" heatid="110816" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.43" />
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="75" swimtime="00:00:49.16" />
                    <SPLIT distance="100" swimtime="00:01:06.90" />
                    <SPLIT distance="125" swimtime="00:01:25.03" />
                    <SPLIT distance="150" swimtime="00:01:43.94" />
                    <SPLIT distance="175" swimtime="00:02:02.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="438" reactiontime="+60" swimtime="00:01:48.75" resultid="107731" heatid="110632" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.60" />
                    <SPLIT distance="50" swimtime="00:00:25.48" />
                    <SPLIT distance="75" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:00:54.23" />
                    <SPLIT distance="125" swimtime="00:01:08.03" />
                    <SPLIT distance="150" swimtime="00:01:23.09" />
                    <SPLIT distance="175" swimtime="00:01:35.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107719" number="1" reactiontime="+60" status="DSQ" />
                    <RELAYPOSITION athleteid="107712" number="2" reactiontime="-66" status="DSQ" />
                    <RELAYPOSITION athleteid="107703" number="3" reactiontime="+24" status="DSQ" />
                    <RELAYPOSITION athleteid="107723" number="4" reactiontime="+41" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="393" swimtime="00:02:03.51" resultid="107732" heatid="110838" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                    <SPLIT distance="75" swimtime="00:00:46.29" />
                    <SPLIT distance="100" swimtime="00:01:07.27" />
                    <SPLIT distance="125" swimtime="00:01:19.19" />
                    <SPLIT distance="150" swimtime="00:01:34.33" />
                    <SPLIT distance="175" swimtime="00:01:48.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107723" number="1" />
                    <RELAYPOSITION athleteid="107712" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="107719" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="107703" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" nation="POL" region="MAL" clubid="107889" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Tomasz Doniec" phone="693703490" />
          <ATHLETES>
            <ATHLETE birthdate="1978-09-01" firstname="Grzegorz" gender="M" lastname="Grzybczyk" nation="POL" athleteid="107947">
              <RESULTS>
                <RESULT eventid="98798" points="149" reactiontime="+96" swimtime="00:00:38.15" resultid="107948" heatid="110598" lane="7" entrytime="00:00:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="78" reactiontime="+100" swimtime="00:04:15.78" resultid="107949" heatid="110619" lane="8">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.10" />
                    <SPLIT distance="50" swimtime="00:00:53.60" />
                    <SPLIT distance="75" swimtime="00:01:27.56" />
                    <SPLIT distance="100" swimtime="00:02:04.41" />
                    <SPLIT distance="125" swimtime="00:02:40.99" />
                    <SPLIT distance="150" swimtime="00:03:17.68" />
                    <SPLIT distance="175" swimtime="00:03:46.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="71" reactiontime="+88" swimtime="00:00:53.64" resultid="107950" heatid="110652" lane="8" entrytime="00:00:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="92" swimtime="00:04:26.31" resultid="107951" heatid="110666" lane="0" entrytime="00:04:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.53" />
                    <SPLIT distance="50" swimtime="00:00:58.00" />
                    <SPLIT distance="75" swimtime="00:01:29.88" />
                    <SPLIT distance="100" swimtime="00:02:05.61" />
                    <SPLIT distance="125" swimtime="00:02:40.19" />
                    <SPLIT distance="150" swimtime="00:03:16.52" />
                    <SPLIT distance="175" swimtime="00:03:51.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="102" reactiontime="+106" swimtime="00:01:58.71" resultid="107952" heatid="110727" lane="5" entrytime="00:01:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.01" />
                    <SPLIT distance="50" swimtime="00:00:56.60" />
                    <SPLIT distance="75" swimtime="00:01:27.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="65" reactiontime="+90" swimtime="00:02:01.61" resultid="107953" heatid="110757" lane="5" entrytime="00:02:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.81" />
                    <SPLIT distance="50" swimtime="00:00:56.98" />
                    <SPLIT distance="75" swimtime="00:01:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="55" reactiontime="+106" swimtime="00:04:36.91" resultid="107954" heatid="110810" lane="7">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.31" />
                    <SPLIT distance="50" swimtime="00:01:03.04" />
                    <SPLIT distance="75" swimtime="00:01:37.69" />
                    <SPLIT distance="100" swimtime="00:02:13.66" />
                    <SPLIT distance="125" swimtime="00:02:50.63" />
                    <SPLIT distance="150" swimtime="00:03:27.00" />
                    <SPLIT distance="175" swimtime="00:04:05.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="92" reactiontime="+128" swimtime="00:00:55.74" resultid="107955" heatid="110825" lane="1" entrytime="00:00:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-25" firstname="Jerzy" gender="M" lastname="Korba" nation="POL" athleteid="107929">
              <RESULTS>
                <RESULT eventid="98798" points="425" reactiontime="+73" swimtime="00:00:26.93" resultid="107930" heatid="110608" lane="2" entrytime="00:00:27.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="392" reactiontime="+87" swimtime="00:10:05.43" resultid="107931" heatid="110636" lane="5" entrytime="00:10:49.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.07" />
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="75" swimtime="00:00:49.67" />
                    <SPLIT distance="100" swimtime="00:01:07.63" />
                    <SPLIT distance="125" swimtime="00:01:26.10" />
                    <SPLIT distance="150" swimtime="00:01:44.81" />
                    <SPLIT distance="175" swimtime="00:02:03.73" />
                    <SPLIT distance="200" swimtime="00:02:22.70" />
                    <SPLIT distance="225" swimtime="00:02:41.61" />
                    <SPLIT distance="250" swimtime="00:03:00.63" />
                    <SPLIT distance="275" swimtime="00:03:19.71" />
                    <SPLIT distance="300" swimtime="00:03:38.82" />
                    <SPLIT distance="325" swimtime="00:03:58.03" />
                    <SPLIT distance="350" swimtime="00:04:17.36" />
                    <SPLIT distance="375" swimtime="00:04:36.74" />
                    <SPLIT distance="400" swimtime="00:04:56.31" />
                    <SPLIT distance="425" swimtime="00:05:15.68" />
                    <SPLIT distance="450" swimtime="00:05:35.02" />
                    <SPLIT distance="475" swimtime="00:05:54.33" />
                    <SPLIT distance="500" swimtime="00:06:13.68" />
                    <SPLIT distance="525" swimtime="00:06:32.97" />
                    <SPLIT distance="550" swimtime="00:06:52.38" />
                    <SPLIT distance="575" swimtime="00:07:11.82" />
                    <SPLIT distance="600" swimtime="00:07:31.24" />
                    <SPLIT distance="625" swimtime="00:08:29.26" />
                    <SPLIT distance="650" swimtime="00:08:09.92" />
                    <SPLIT distance="675" swimtime="00:09:08.43" />
                    <SPLIT distance="700" swimtime="00:08:48.96" />
                    <SPLIT distance="725" swimtime="00:09:47.48" />
                    <SPLIT distance="750" swimtime="00:09:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="339" reactiontime="+90" swimtime="00:02:52.72" resultid="107932" heatid="110668" lane="1" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.79" />
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="75" swimtime="00:00:59.63" />
                    <SPLIT distance="100" swimtime="00:01:22.07" />
                    <SPLIT distance="125" swimtime="00:01:44.77" />
                    <SPLIT distance="150" swimtime="00:02:07.95" />
                    <SPLIT distance="175" swimtime="00:02:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="447" reactiontime="+80" swimtime="00:00:58.75" resultid="107933" heatid="110687" lane="6" entrytime="00:00:59.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                    <SPLIT distance="75" swimtime="00:00:43.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="406" reactiontime="+80" swimtime="00:01:15.09" resultid="107934" heatid="110733" lane="1" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.80" />
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="75" swimtime="00:00:54.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="401" reactiontime="+79" swimtime="00:02:14.68" resultid="107935" heatid="110776" lane="2" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.70" />
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="75" swimtime="00:00:48.71" />
                    <SPLIT distance="100" swimtime="00:01:06.12" />
                    <SPLIT distance="125" swimtime="00:01:23.63" />
                    <SPLIT distance="150" swimtime="00:01:41.37" />
                    <SPLIT distance="175" swimtime="00:01:59.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="447" reactiontime="+77" swimtime="00:00:33.02" resultid="107936" heatid="110832" lane="7" entrytime="00:00:34.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="107937" heatid="110845" lane="8" entrytime="00:05:05.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-03-06" firstname="Ewa" gender="F" lastname="Rupp" nation="POL" athleteid="107901">
              <RESULTS>
                <RESULT eventid="98777" points="107" reactiontime="+137" swimtime="00:00:48.87" resultid="107902" heatid="110587" lane="0" entrytime="00:00:46.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="87" reactiontime="+107" swimtime="00:04:34.36" resultid="107903" heatid="110614" lane="6" entrytime="00:04:49.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.02" />
                    <SPLIT distance="50" swimtime="00:01:02.51" />
                    <SPLIT distance="75" swimtime="00:01:37.37" />
                    <SPLIT distance="100" swimtime="00:02:13.76" />
                    <SPLIT distance="125" swimtime="00:02:53.30" />
                    <SPLIT distance="150" swimtime="00:03:31.27" />
                    <SPLIT distance="175" swimtime="00:04:03.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="89" reactiontime="+72" swimtime="00:00:57.42" resultid="107904" heatid="110646" lane="6" entrytime="00:00:56.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="42" reactiontime="+114" swimtime="00:05:42.93" resultid="107905" heatid="110707" lane="7">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.72" />
                    <SPLIT distance="50" swimtime="00:01:03.69" />
                    <SPLIT distance="75" swimtime="00:01:43.14" />
                    <SPLIT distance="100" swimtime="00:02:28.34" />
                    <SPLIT distance="125" swimtime="00:03:18.54" />
                    <SPLIT distance="150" swimtime="00:04:07.88" />
                    <SPLIT distance="175" swimtime="00:04:58.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="61" reactiontime="+116" swimtime="00:01:01.85" resultid="107906" heatid="110736" lane="1" entrytime="00:00:58.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="75" reactiontime="+82" swimtime="00:02:10.17" resultid="107907" heatid="110753" lane="5" entrytime="00:02:03.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.88" />
                    <SPLIT distance="50" swimtime="00:01:01.98" />
                    <SPLIT distance="75" swimtime="00:01:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="68" reactiontime="+121" swimtime="00:02:13.19" resultid="107908" heatid="110793" lane="3" entrytime="00:02:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.56" />
                    <SPLIT distance="50" swimtime="00:01:03.05" />
                    <SPLIT distance="75" swimtime="00:01:38.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="84" reactiontime="+44" swimtime="00:04:32.13" resultid="107909" heatid="110806" lane="6" entrytime="00:04:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.44" />
                    <SPLIT distance="50" swimtime="00:01:02.64" />
                    <SPLIT distance="75" swimtime="00:01:38.02" />
                    <SPLIT distance="100" swimtime="00:02:13.56" />
                    <SPLIT distance="125" swimtime="00:02:50.50" />
                    <SPLIT distance="150" swimtime="00:03:26.22" />
                    <SPLIT distance="175" swimtime="00:04:00.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="107938">
              <RESULTS>
                <RESULT eventid="98777" points="593" reactiontime="+67" swimtime="00:00:27.66" resultid="107939" heatid="110593" lane="6" entrytime="00:00:27.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="602" reactiontime="+62" swimtime="00:02:24.27" resultid="107940" heatid="110618" lane="4" entrytime="00:02:25.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.08" />
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="75" swimtime="00:00:50.02" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="125" swimtime="00:01:29.16" />
                    <SPLIT distance="150" swimtime="00:01:50.10" />
                    <SPLIT distance="175" swimtime="00:02:07.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="627" reactiontime="+65" swimtime="00:00:59.45" resultid="107941" heatid="110676" lane="4" entrytime="00:00:59.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                    <SPLIT distance="75" swimtime="00:00:44.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="593" reactiontime="+58" swimtime="00:01:07.44" resultid="107942" heatid="110695" lane="4" entrytime="00:01:07.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                    <SPLIT distance="75" swimtime="00:00:51.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="595" reactiontime="+65" swimtime="00:01:14.13" resultid="107943" heatid="110725" lane="4" entrytime="00:01:14.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.96" />
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="75" swimtime="00:00:54.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="640" reactiontime="+66" swimtime="00:02:08.53" resultid="107944" heatid="110768" lane="4" entrytime="00:02:09.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.94" />
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                    <SPLIT distance="75" swimtime="00:00:45.20" />
                    <SPLIT distance="100" swimtime="00:01:01.67" />
                    <SPLIT distance="125" swimtime="00:01:18.06" />
                    <SPLIT distance="150" swimtime="00:01:34.90" />
                    <SPLIT distance="175" swimtime="00:01:52.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="518" reactiontime="+77" swimtime="00:01:07.97" resultid="107945" heatid="110796" lane="5" entrytime="00:01:09.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.55" />
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="75" swimtime="00:00:49.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="593" reactiontime="+72" swimtime="00:00:34.27" resultid="107946" heatid="110823" lane="4" entrytime="00:00:34.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-11-06" firstname="Małgorzata" gender="F" lastname="Wach" nation="POL" athleteid="107914">
              <RESULTS>
                <RESULT comment="O4" eventid="98777" reactiontime="+58" status="DSQ" swimtime="00:00:00.00" resultid="107915" heatid="110589" lane="1" entrytime="00:00:35.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="258" reactiontime="+66" swimtime="00:00:40.31" resultid="107916" heatid="110648" lane="5" entrytime="00:00:39.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4" eventid="98907" status="DSQ" swimtime="00:00:00.00" resultid="107917" heatid="110673" lane="6" entrytime="00:01:21.00" entrycourse="SCM" />
                <RESULT eventid="99314" points="250" reactiontime="+65" swimtime="00:01:27.29" resultid="107918" heatid="110755" lane="8" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.36" />
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                    <SPLIT distance="75" swimtime="00:01:06.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="221" swimtime="00:03:03.12" resultid="107919" heatid="110766" lane="0" entrytime="00:02:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.64" />
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                    <SPLIT distance="75" swimtime="00:01:03.03" />
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                    <SPLIT distance="125" swimtime="00:01:51.88" />
                    <SPLIT distance="150" swimtime="00:02:16.18" />
                    <SPLIT distance="175" swimtime="00:02:40.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="212" reactiontime="+72" swimtime="00:03:19.87" resultid="107920" heatid="110807" lane="4" entrytime="00:03:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.21" />
                    <SPLIT distance="50" swimtime="00:00:46.02" />
                    <SPLIT distance="75" swimtime="00:01:12.11" />
                    <SPLIT distance="100" swimtime="00:01:38.13" />
                    <SPLIT distance="125" swimtime="00:02:05.06" />
                    <SPLIT distance="150" swimtime="00:02:30.92" />
                    <SPLIT distance="175" swimtime="00:02:56.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="250" reactiontime="+93" swimtime="00:00:45.70" resultid="107921" heatid="110820" lane="8" entrytime="00:00:46.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-08-12" firstname="Konrad" gender="M" lastname="Plutecki" nation="POL" athleteid="107922">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="107923" heatid="110608" lane="0" entrytime="00:00:27.50" entrycourse="SCM" />
                <RESULT eventid="106277" points="469" reactiontime="+69" swimtime="00:00:57.83" resultid="107924" heatid="110687" lane="8" entrytime="00:00:59.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                    <SPLIT distance="75" swimtime="00:00:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="374" reactiontime="+69" swimtime="00:01:17.14" resultid="107925" heatid="110731" lane="5" entrytime="00:01:21.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.36" />
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="75" swimtime="00:00:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="411" reactiontime="+68" swimtime="00:02:13.62" resultid="107926" heatid="110775" lane="4" entrytime="00:02:19.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="75" swimtime="00:00:46.37" />
                    <SPLIT distance="100" swimtime="00:01:03.10" />
                    <SPLIT distance="125" swimtime="00:01:20.29" />
                    <SPLIT distance="150" swimtime="00:01:37.89" />
                    <SPLIT distance="175" swimtime="00:01:56.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="313" reactiontime="+71" swimtime="00:02:35.44" resultid="107927" heatid="110815" lane="8" entrytime="00:02:35.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.27" />
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                    <SPLIT distance="75" swimtime="00:00:56.20" />
                    <SPLIT distance="100" swimtime="00:01:15.93" />
                    <SPLIT distance="125" swimtime="00:01:35.77" />
                    <SPLIT distance="150" swimtime="00:01:55.97" />
                    <SPLIT distance="175" swimtime="00:02:15.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="107928" heatid="110845" lane="3" entrytime="00:04:59.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-19" firstname="Paulina" gender="F" lastname="Palka" nation="POL" athleteid="107910">
              <RESULTS>
                <RESULT eventid="106294" points="436" reactiontime="+55" swimtime="00:00:33.84" resultid="107911" heatid="110649" lane="5" entrytime="00:00:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="423" reactiontime="+63" swimtime="00:01:13.28" resultid="107912" heatid="110756" lane="7" entrytime="00:01:15.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.25" />
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="75" swimtime="00:00:54.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="389" reactiontime="+59" swimtime="00:02:43.30" resultid="107913" heatid="110809" lane="6" entrytime="00:02:50.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.66" />
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="75" swimtime="00:00:59.82" />
                    <SPLIT distance="100" swimtime="00:01:20.99" />
                    <SPLIT distance="125" swimtime="00:01:42.19" />
                    <SPLIT distance="150" swimtime="00:02:03.47" />
                    <SPLIT distance="175" swimtime="00:02:23.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Wisła Team 1" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="149" swimtime="00:02:35.66" resultid="107956" heatid="110630" lane="9" entrytime="00:02:45.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.32" />
                    <SPLIT distance="50" swimtime="00:00:50.16" />
                    <SPLIT distance="75" swimtime="00:01:03.93" />
                    <SPLIT distance="100" swimtime="00:01:18.23" />
                    <SPLIT distance="125" swimtime="00:01:35.67" />
                    <SPLIT distance="150" swimtime="00:01:55.73" />
                    <SPLIT distance="175" swimtime="00:02:13.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107901" number="1" />
                    <RELAYPOSITION athleteid="107929" number="2" />
                    <RELAYPOSITION athleteid="107914" number="3" />
                    <RELAYPOSITION athleteid="107947" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Wisła Team 2" number="2">
              <RESULTS>
                <RESULT eventid="99441" points="146" reactiontime="+59" swimtime="00:02:51.68" resultid="107957" heatid="110836" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.13" />
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="75" swimtime="00:00:58.35" />
                    <SPLIT distance="100" swimtime="00:01:26.85" />
                    <SPLIT distance="125" swimtime="00:01:52.02" />
                    <SPLIT distance="150" swimtime="00:02:24.50" />
                    <SPLIT distance="175" swimtime="00:02:37.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107910" number="1" reactiontime="+59" />
                    <RELAYPOSITION athleteid="107947" number="2" />
                    <RELAYPOSITION athleteid="107901" number="3" />
                    <RELAYPOSITION athleteid="107929" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="106964" name="MASTERS Zdzieszowice">
          <CONTACT city="Zdzieszowice" email="masters.zdzieszowice@gmail.com" name="Jajuga" phone="505127695" street="Dworcowa 4" zip="47-330" />
          <ATHLETES>
            <ATHLETE birthdate="1986-06-13" firstname="Magdalena" gender="F" lastname="Gorostiza" nation="POL" athleteid="106986">
              <RESULTS>
                <RESULT eventid="98814" points="260" swimtime="00:03:10.86" resultid="106987" heatid="110616" lane="9" entrytime="00:03:15.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.45" />
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="75" swimtime="00:01:07.92" />
                    <SPLIT distance="100" swimtime="00:01:33.46" />
                    <SPLIT distance="125" swimtime="00:01:58.98" />
                    <SPLIT distance="150" swimtime="00:02:25.49" />
                    <SPLIT distance="175" swimtime="00:02:49.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="288" reactiontime="+92" swimtime="00:03:23.61" resultid="106988" heatid="110663" lane="4" entrytime="00:03:15.78">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.59" />
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                    <SPLIT distance="75" swimtime="00:01:10.20" />
                    <SPLIT distance="100" swimtime="00:01:35.96" />
                    <SPLIT distance="125" swimtime="00:02:03.19" />
                    <SPLIT distance="150" swimtime="00:02:29.98" />
                    <SPLIT distance="175" swimtime="00:02:57.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="315" reactiontime="+91" swimtime="00:01:31.62" resultid="106989" heatid="110720" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.75" />
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                    <SPLIT distance="75" swimtime="00:01:07.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="302" reactiontime="+89" swimtime="00:00:36.31" resultid="106990" heatid="110738" lane="3" entrytime="00:00:37.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="229" reactiontime="+90" swimtime="00:01:29.20" resultid="106991" heatid="110794" lane="7" entrytime="00:01:40.96">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.64" />
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="75" swimtime="00:01:04.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="383" reactiontime="+97" swimtime="00:00:39.65" resultid="106992" heatid="110821" lane="3" entrytime="00:00:40.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-18" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="106981">
              <RESULTS>
                <RESULT eventid="98814" points="304" swimtime="00:03:01.18" resultid="106982" heatid="110617" lane="9" entrytime="00:03:03.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.18" />
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="75" swimtime="00:01:02.02" />
                    <SPLIT distance="100" swimtime="00:01:24.42" />
                    <SPLIT distance="125" swimtime="00:01:51.21" />
                    <SPLIT distance="150" swimtime="00:02:18.68" />
                    <SPLIT distance="175" swimtime="00:02:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="342" reactiontime="+100" swimtime="00:01:20.97" resultid="106983" heatid="110693" lane="3" entrytime="00:01:24.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="75" swimtime="00:01:01.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="318" reactiontime="+83" swimtime="00:01:20.57" resultid="106984" heatid="110755" lane="5" entrytime="00:01:24.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.65" />
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="75" swimtime="00:01:00.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="323" reactiontime="+77" swimtime="00:02:53.77" resultid="106985" heatid="110809" lane="0" entrytime="00:03:01.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.35" />
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="75" swimtime="00:01:03.34" />
                    <SPLIT distance="100" swimtime="00:01:25.17" />
                    <SPLIT distance="125" swimtime="00:01:47.68" />
                    <SPLIT distance="150" swimtime="00:02:10.28" />
                    <SPLIT distance="175" swimtime="00:02:32.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="106972">
              <RESULTS>
                <RESULT eventid="98830" points="497" reactiontime="+73" swimtime="00:02:18.32" resultid="106973" heatid="110628" lane="6" entrytime="00:02:18.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.83" />
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="75" swimtime="00:00:47.32" />
                    <SPLIT distance="100" swimtime="00:01:05.43" />
                    <SPLIT distance="125" swimtime="00:01:25.37" />
                    <SPLIT distance="150" swimtime="00:01:46.07" />
                    <SPLIT distance="175" swimtime="00:02:02.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="524" reactiontime="+82" swimtime="00:01:02.81" resultid="106975" heatid="110696" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.59" />
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                    <SPLIT distance="75" swimtime="00:00:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="432" reactiontime="+73" swimtime="00:02:23.50" resultid="106976" heatid="110713" lane="2" entrytime="00:02:20.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.51" />
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="75" swimtime="00:00:49.62" />
                    <SPLIT distance="100" swimtime="00:01:07.95" />
                    <SPLIT distance="125" swimtime="00:01:26.68" />
                    <SPLIT distance="150" swimtime="00:01:45.50" />
                    <SPLIT distance="175" swimtime="00:02:04.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="492" swimtime="00:02:05.81" resultid="106977" heatid="110778" lane="9" entrytime="00:02:05.66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:28.27" />
                    <SPLIT distance="75" swimtime="00:00:44.05" />
                    <SPLIT distance="100" swimtime="00:01:00.56" />
                    <SPLIT distance="125" swimtime="00:01:16.72" />
                    <SPLIT distance="150" swimtime="00:01:33.44" />
                    <SPLIT distance="175" swimtime="00:01:50.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="463" reactiontime="+84" swimtime="00:05:04.28" resultid="106978" heatid="110792" lane="3" entrytime="00:05:08.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.83" />
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="75" swimtime="00:00:48.32" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="125" swimtime="00:01:26.83" />
                    <SPLIT distance="150" swimtime="00:01:46.40" />
                    <SPLIT distance="175" swimtime="00:02:06.50" />
                    <SPLIT distance="200" swimtime="00:02:26.21" />
                    <SPLIT distance="225" swimtime="00:02:47.89" />
                    <SPLIT distance="250" swimtime="00:03:09.56" />
                    <SPLIT distance="275" swimtime="00:03:31.50" />
                    <SPLIT distance="300" swimtime="00:03:53.83" />
                    <SPLIT distance="325" swimtime="00:04:11.95" />
                    <SPLIT distance="350" swimtime="00:04:29.59" />
                    <SPLIT distance="375" swimtime="00:04:47.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="517" reactiontime="+77" swimtime="00:01:00.33" resultid="106979" heatid="110804" lane="4" entrytime="00:01:00.75">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="75" swimtime="00:00:43.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="444" swimtime="00:04:38.20" resultid="106980" heatid="110843" lane="0" entrytime="00:04:38.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.13" />
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="75" swimtime="00:00:49.61" />
                    <SPLIT distance="100" swimtime="00:01:07.34" />
                    <SPLIT distance="125" swimtime="00:01:25.00" />
                    <SPLIT distance="150" swimtime="00:01:42.53" />
                    <SPLIT distance="175" swimtime="00:02:00.27" />
                    <SPLIT distance="200" swimtime="00:02:18.38" />
                    <SPLIT distance="225" swimtime="00:02:36.01" />
                    <SPLIT distance="250" swimtime="00:02:53.88" />
                    <SPLIT distance="275" swimtime="00:03:11.57" />
                    <SPLIT distance="300" swimtime="00:03:29.40" />
                    <SPLIT distance="325" swimtime="00:03:47.15" />
                    <SPLIT distance="350" swimtime="00:04:05.08" />
                    <SPLIT distance="375" swimtime="00:04:22.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="347" reactiontime="+92" swimtime="00:20:06.56" resultid="110856" heatid="110642" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.87" />
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="75" swimtime="00:00:52.47" />
                    <SPLIT distance="100" swimtime="00:01:11.55" />
                    <SPLIT distance="125" swimtime="00:01:30.72" />
                    <SPLIT distance="150" swimtime="00:01:50.08" />
                    <SPLIT distance="175" swimtime="00:02:09.58" />
                    <SPLIT distance="200" swimtime="00:02:28.77" />
                    <SPLIT distance="225" swimtime="00:02:48.05" />
                    <SPLIT distance="250" swimtime="00:03:07.37" />
                    <SPLIT distance="275" swimtime="00:03:26.28" />
                    <SPLIT distance="300" swimtime="00:03:45.52" />
                    <SPLIT distance="325" swimtime="00:04:05.02" />
                    <SPLIT distance="350" swimtime="00:04:24.53" />
                    <SPLIT distance="375" swimtime="00:04:43.92" />
                    <SPLIT distance="400" swimtime="00:05:03.57" />
                    <SPLIT distance="425" swimtime="00:05:23.02" />
                    <SPLIT distance="450" swimtime="00:05:42.90" />
                    <SPLIT distance="475" swimtime="00:06:02.53" />
                    <SPLIT distance="500" swimtime="00:06:22.45" />
                    <SPLIT distance="525" swimtime="00:06:42.32" />
                    <SPLIT distance="550" swimtime="00:07:02.51" />
                    <SPLIT distance="575" swimtime="00:07:22.34" />
                    <SPLIT distance="600" swimtime="00:07:42.60" />
                    <SPLIT distance="625" swimtime="00:08:02.62" />
                    <SPLIT distance="650" swimtime="00:08:22.88" />
                    <SPLIT distance="675" swimtime="00:08:42.96" />
                    <SPLIT distance="700" swimtime="00:09:03.61" />
                    <SPLIT distance="725" swimtime="00:09:23.98" />
                    <SPLIT distance="750" swimtime="00:09:44.55" />
                    <SPLIT distance="775" swimtime="00:10:04.94" />
                    <SPLIT distance="800" swimtime="00:10:25.57" />
                    <SPLIT distance="825" swimtime="00:10:45.84" />
                    <SPLIT distance="850" swimtime="00:11:06.42" />
                    <SPLIT distance="875" swimtime="00:11:26.95" />
                    <SPLIT distance="900" swimtime="00:11:47.89" />
                    <SPLIT distance="925" swimtime="00:12:08.62" />
                    <SPLIT distance="950" swimtime="00:12:29.43" />
                    <SPLIT distance="975" swimtime="00:12:49.98" />
                    <SPLIT distance="1000" swimtime="00:13:10.74" />
                    <SPLIT distance="1025" swimtime="00:13:31.23" />
                    <SPLIT distance="1050" swimtime="00:13:52.05" />
                    <SPLIT distance="1075" swimtime="00:14:12.46" />
                    <SPLIT distance="1100" swimtime="00:14:33.40" />
                    <SPLIT distance="1125" swimtime="00:14:54.40" />
                    <SPLIT distance="1150" swimtime="00:15:15.32" />
                    <SPLIT distance="1175" swimtime="00:15:36.00" />
                    <SPLIT distance="1200" swimtime="00:15:57.07" />
                    <SPLIT distance="1225" swimtime="00:16:17.81" />
                    <SPLIT distance="1250" swimtime="00:16:38.67" />
                    <SPLIT distance="1275" swimtime="00:16:59.60" />
                    <SPLIT distance="1300" swimtime="00:17:20.77" />
                    <SPLIT distance="1325" swimtime="00:17:41.66" />
                    <SPLIT distance="1350" swimtime="00:18:02.74" />
                    <SPLIT distance="1375" swimtime="00:18:23.68" />
                    <SPLIT distance="1400" swimtime="00:18:44.77" />
                    <SPLIT distance="1425" swimtime="00:19:05.59" />
                    <SPLIT distance="1450" swimtime="00:19:26.77" />
                    <SPLIT distance="1475" swimtime="00:19:47.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-08" firstname="Przemysław" gender="M" lastname="Osiwała" nation="POL" athleteid="106965">
              <RESULTS>
                <RESULT eventid="98830" points="321" reactiontime="+91" swimtime="00:02:39.95" resultid="106966" heatid="110624" lane="3" entrytime="00:02:44.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.46" />
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="75" swimtime="00:00:55.65" />
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                    <SPLIT distance="125" swimtime="00:01:40.02" />
                    <SPLIT distance="150" swimtime="00:02:03.70" />
                    <SPLIT distance="175" swimtime="00:02:22.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="290" reactiontime="+95" swimtime="00:03:01.90" resultid="106967" heatid="110669" lane="3" entrytime="00:02:50.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.89" />
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                    <SPLIT distance="75" swimtime="00:01:03.47" />
                    <SPLIT distance="100" swimtime="00:01:26.63" />
                    <SPLIT distance="125" swimtime="00:01:50.21" />
                    <SPLIT distance="150" swimtime="00:02:14.25" />
                    <SPLIT distance="175" swimtime="00:02:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="324" swimtime="00:02:37.96" resultid="106968" heatid="110713" lane="0" entrytime="00:02:38.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.13" />
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="75" swimtime="00:00:55.59" />
                    <SPLIT distance="100" swimtime="00:01:16.06" />
                    <SPLIT distance="125" swimtime="00:01:36.49" />
                    <SPLIT distance="150" swimtime="00:01:57.03" />
                    <SPLIT distance="175" swimtime="00:02:17.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="358" reactiontime="+87" swimtime="00:00:30.70" resultid="106969" heatid="110746" lane="3" entrytime="00:00:31.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.18" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z2/G3" eventid="99282" reactiontime="+86" status="DSQ" swimtime="00:00:00.00" resultid="106970" heatid="110791" lane="7" entrytime="00:05:50.34" />
                <RESULT eventid="99361" points="345" swimtime="00:01:09.00" resultid="106971" heatid="110804" lane="9" entrytime="00:01:07.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="75" swimtime="00:00:49.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="253" reactiontime="+83" swimtime="00:02:10.57" resultid="106993" heatid="110630" lane="7" entrytime="00:02:22.22">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.27" />
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="75" swimtime="00:00:48.93" />
                    <SPLIT distance="100" swimtime="00:01:06.65" />
                    <SPLIT distance="125" swimtime="00:01:22.86" />
                    <SPLIT distance="150" swimtime="00:01:41.15" />
                    <SPLIT distance="175" swimtime="00:01:55.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106972" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="106981" number="2" reactiontime="+79" />
                    <RELAYPOSITION athleteid="106986" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="106965" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="317" reactiontime="+77" swimtime="00:02:12.73" resultid="106994" heatid="110837" lane="9" entrytime="00:02:22.22">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.74" />
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="75" swimtime="00:00:55.23" />
                    <SPLIT distance="100" swimtime="00:01:17.12" />
                    <SPLIT distance="125" swimtime="00:01:30.81" />
                    <SPLIT distance="150" swimtime="00:01:47.41" />
                    <SPLIT distance="175" swimtime="00:01:59.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106981" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="106986" number="2" />
                    <RELAYPOSITION athleteid="106965" number="3" />
                    <RELAYPOSITION athleteid="106972" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="107551" name="MASTERS Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos Rafał" phone="604184311" />
          <ATHLETES>
            <ATHLETE birthdate="1980-04-14" firstname="Damian" gender="M" lastname="Karkusiński" nation="POL" athleteid="107614">
              <RESULTS>
                <RESULT eventid="98798" points="307" reactiontime="+75" swimtime="00:00:30.01" resultid="107615" heatid="110603" lane="5" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="236" reactiontime="+64" swimtime="00:00:35.95" resultid="107616" heatid="110658" lane="9" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="251" swimtime="00:01:11.15" resultid="107617" heatid="110684" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.91" />
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="75" swimtime="00:00:50.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-11-02" firstname="Ksawery" gender="M" lastname="Wiaderek" nation="POL" athleteid="107628">
              <RESULTS>
                <RESULT eventid="98798" points="451" reactiontime="+85" swimtime="00:00:26.41" resultid="107629" heatid="110608" lane="8" entrytime="00:00:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="429" reactiontime="+95" swimtime="00:00:59.58" resultid="107630" heatid="110684" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="75" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="425" reactiontime="+88" swimtime="00:00:28.99" resultid="107631" heatid="110748" lane="7" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-11-12" firstname="Witold" gender="M" lastname="Pietrowski" nation="POL" athleteid="107624">
              <RESULTS>
                <RESULT eventid="98798" points="321" reactiontime="+82" swimtime="00:00:29.58" resultid="107625" heatid="110605" lane="7" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="238" reactiontime="+76" swimtime="00:00:35.84" resultid="107626" heatid="110656" lane="7" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="300" reactiontime="+95" swimtime="00:00:32.56" resultid="107627" heatid="110745" lane="2" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-18" firstname="Konrad" gender="M" lastname="Hasik" nation="POL" athleteid="107561">
              <RESULTS>
                <RESULT eventid="98830" points="407" reactiontime="+94" swimtime="00:02:27.85" resultid="107562" heatid="110627" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.65" />
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="75" swimtime="00:00:50.56" />
                    <SPLIT distance="100" swimtime="00:01:09.11" />
                    <SPLIT distance="125" swimtime="00:01:30.11" />
                    <SPLIT distance="150" swimtime="00:01:51.65" />
                    <SPLIT distance="175" swimtime="00:02:10.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="382" reactiontime="+74" swimtime="00:00:30.60" resultid="107563" heatid="110658" lane="2" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="260" reactiontime="+88" swimtime="00:02:50.08" resultid="107564" heatid="110712" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.90" />
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="75" swimtime="00:00:57.44" />
                    <SPLIT distance="100" swimtime="00:01:19.28" />
                    <SPLIT distance="125" swimtime="00:01:42.27" />
                    <SPLIT distance="150" swimtime="00:02:05.66" />
                    <SPLIT distance="175" swimtime="00:02:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="384" reactiontime="+84" swimtime="00:01:16.46" resultid="107565" heatid="110733" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.96" />
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="75" swimtime="00:00:56.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="400" reactiontime="+69" swimtime="00:01:06.38" resultid="107566" heatid="110763" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.31" />
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                    <SPLIT distance="75" swimtime="00:00:49.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="312" reactiontime="+69" swimtime="00:02:35.64" resultid="107567" heatid="110814" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.95" />
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="75" swimtime="00:00:57.14" />
                    <SPLIT distance="100" swimtime="00:01:17.79" />
                    <SPLIT distance="125" swimtime="00:01:38.95" />
                    <SPLIT distance="150" swimtime="00:01:59.25" />
                    <SPLIT distance="175" swimtime="00:02:18.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="433" reactiontime="+78" swimtime="00:00:33.36" resultid="107568" heatid="110831" lane="4" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-14" firstname="Jakub" gender="M" lastname="Gryczyński" nation="POL" athleteid="107574">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="107575" heatid="110602" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="107576" heatid="110698" lane="6" entrytime="00:01:25.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="107577" heatid="110729" lane="2" entrytime="00:01:35.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="107578" heatid="110827" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-10-05" firstname="Marcin" gender="M" lastname="Grabarczyk" nation="POL" athleteid="107588">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="107589" heatid="110609" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="98830" points="317" reactiontime="+81" swimtime="00:02:40.70" resultid="107590" heatid="110625" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.46" />
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                    <SPLIT distance="75" swimtime="00:00:53.04" />
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                    <SPLIT distance="125" swimtime="00:01:36.73" />
                    <SPLIT distance="150" swimtime="00:02:00.87" />
                    <SPLIT distance="175" swimtime="00:02:21.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="250" reactiontime="+94" swimtime="00:03:11.19" resultid="107591" heatid="110669" lane="2" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.81" />
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="75" swimtime="00:01:05.11" />
                    <SPLIT distance="100" swimtime="00:01:29.35" />
                    <SPLIT distance="125" swimtime="00:01:54.58" />
                    <SPLIT distance="150" swimtime="00:02:20.37" />
                    <SPLIT distance="175" swimtime="00:02:46.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="369" reactiontime="+78" swimtime="00:01:10.60" resultid="107592" heatid="110702" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.15" />
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="75" swimtime="00:00:53.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="308" reactiontime="+82" swimtime="00:01:22.28" resultid="107593" heatid="110731" lane="4" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.16" />
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="75" swimtime="00:00:59.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="107594" heatid="110776" lane="1" entrytime="00:02:17.00" />
                <RESULT eventid="99425" points="325" swimtime="00:00:36.71" resultid="107595" heatid="110829" lane="9" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="107596" heatid="110845" lane="5" entrytime="00:04:57.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-06-12" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" athleteid="107569">
              <RESULTS>
                <RESULT eventid="98798" points="443" reactiontime="+86" swimtime="00:00:26.56" resultid="107570" heatid="110610" lane="0" entrytime="00:00:26.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="446" reactiontime="+82" swimtime="00:00:58.79" resultid="107571" heatid="110686" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                    <SPLIT distance="75" swimtime="00:00:43.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="413" swimtime="00:00:29.26" resultid="107572" heatid="110749" lane="6" entrytime="00:00:28.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="389" swimtime="00:01:06.31" resultid="107573" heatid="110804" lane="0" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.87" />
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="75" swimtime="00:00:47.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-02" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="107597">
              <RESULTS>
                <RESULT eventid="98798" points="422" reactiontime="+102" swimtime="00:00:27.01" resultid="107598" heatid="110609" lane="3" entrytime="00:00:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="362" swimtime="00:01:03.03" resultid="107599" heatid="110684" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.77" />
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="75" swimtime="00:00:45.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="344" reactiontime="+77" swimtime="00:00:31.10" resultid="107600" heatid="110745" lane="5" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="367" reactiontime="+90" swimtime="00:00:35.25" resultid="107601" heatid="110831" lane="3" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-08-19" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" athleteid="107602">
              <RESULTS>
                <RESULT eventid="98798" points="308" swimtime="00:00:29.97" resultid="107603" heatid="110603" lane="9" entrytime="00:00:30.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="254" reactiontime="+75" swimtime="00:01:19.99" resultid="107604" heatid="110698" lane="5" entrytime="00:01:21.66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.47" />
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="75" swimtime="00:00:59.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="74" reactiontime="+88" swimtime="00:01:56.44" resultid="107605" heatid="110760" lane="1" entrytime="00:01:24.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.65" />
                    <SPLIT distance="50" swimtime="00:01:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="107606" heatid="110828" lane="8" entrytime="00:00:39.84" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-08" firstname="Marcin" gender="M" lastname="Babuchowski" nation="POL" athleteid="107618">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="107619" heatid="110613" lane="8" entrytime="00:00:24.00" />
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="107620" heatid="110689" lane="4" entrytime="00:00:52.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="107621" heatid="110751" lane="5" entrytime="00:00:24.60" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="107622" heatid="110778" lane="2" entrytime="00:01:58.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="107623" heatid="110805" lane="5" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-11" firstname="Przemysław" gender="M" lastname="Michniewski" nation="POL" athleteid="107607">
              <RESULTS>
                <RESULT eventid="98798" points="407" reactiontime="+79" swimtime="00:00:27.32" resultid="107608" heatid="110603" lane="6" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="330" reactiontime="+96" swimtime="00:02:38.58" resultid="107609" heatid="110627" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                    <SPLIT distance="75" swimtime="00:00:51.21" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="125" swimtime="00:01:33.94" />
                    <SPLIT distance="150" swimtime="00:01:57.11" />
                    <SPLIT distance="175" swimtime="00:02:18.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="393" reactiontime="+93" swimtime="00:01:09.12" resultid="107610" heatid="110702" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.70" />
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="75" swimtime="00:00:51.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="406" swimtime="00:01:15.07" resultid="107611" heatid="110732" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="75" swimtime="00:00:54.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="389" reactiontime="+89" swimtime="00:00:29.84" resultid="107612" heatid="110747" lane="2" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="420" reactiontime="+75" swimtime="00:00:33.71" resultid="107613" heatid="110833" lane="2" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="107579">
              <RESULTS>
                <RESULT eventid="98798" points="363" reactiontime="+91" swimtime="00:00:28.39" resultid="107580" heatid="110600" lane="1" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="241" reactiontime="+89" swimtime="00:02:56.00" resultid="107581" heatid="110621" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.31" />
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="75" swimtime="00:00:59.61" />
                    <SPLIT distance="100" swimtime="00:01:22.20" />
                    <SPLIT distance="125" swimtime="00:01:47.70" />
                    <SPLIT distance="150" swimtime="00:02:13.58" />
                    <SPLIT distance="175" swimtime="00:02:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="248" reactiontime="+100" swimtime="00:03:11.54" resultid="107582" heatid="110667" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.00" />
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="75" swimtime="00:01:05.01" />
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="125" swimtime="00:01:56.82" />
                    <SPLIT distance="150" swimtime="00:02:23.26" />
                    <SPLIT distance="175" swimtime="00:02:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="261" reactiontime="+93" swimtime="00:01:19.20" resultid="107583" heatid="110697" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.45" />
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                    <SPLIT distance="75" swimtime="00:01:00.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="252" reactiontime="+95" swimtime="00:01:28.00" resultid="107584" heatid="110729" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.43" />
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                    <SPLIT distance="75" swimtime="00:01:04.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="201" reactiontime="+75" swimtime="00:01:23.50" resultid="107585" heatid="110759" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="107586" heatid="110812" lane="4" entrytime="00:03:08.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="107587" heatid="110826" lane="7" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-28" firstname="Artur" gender="M" lastname="Frąckowiak" nation="POL" athleteid="107552">
              <RESULTS>
                <RESULT eventid="98798" points="456" reactiontime="+80" swimtime="00:00:26.32" resultid="107553" heatid="110609" lane="7" entrytime="00:00:26.86">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="386" reactiontime="+94" swimtime="00:10:08.95" resultid="107554" heatid="110635" lane="1" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.07" />
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="75" swimtime="00:00:49.02" />
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                    <SPLIT distance="125" swimtime="00:01:25.52" />
                    <SPLIT distance="150" swimtime="00:01:44.35" />
                    <SPLIT distance="175" swimtime="00:02:03.26" />
                    <SPLIT distance="200" swimtime="00:02:22.37" />
                    <SPLIT distance="225" swimtime="00:02:41.59" />
                    <SPLIT distance="250" swimtime="00:03:01.03" />
                    <SPLIT distance="275" swimtime="00:03:20.25" />
                    <SPLIT distance="300" swimtime="00:03:39.63" />
                    <SPLIT distance="325" swimtime="00:03:59.04" />
                    <SPLIT distance="350" swimtime="00:04:18.64" />
                    <SPLIT distance="375" swimtime="00:04:37.97" />
                    <SPLIT distance="400" swimtime="00:04:57.68" />
                    <SPLIT distance="425" swimtime="00:05:16.98" />
                    <SPLIT distance="450" swimtime="00:05:36.51" />
                    <SPLIT distance="475" swimtime="00:05:55.84" />
                    <SPLIT distance="500" swimtime="00:06:14.93" />
                    <SPLIT distance="525" swimtime="00:06:34.27" />
                    <SPLIT distance="550" swimtime="00:06:53.92" />
                    <SPLIT distance="575" swimtime="00:07:13.08" />
                    <SPLIT distance="600" swimtime="00:07:32.90" />
                    <SPLIT distance="625" swimtime="00:07:52.37" />
                    <SPLIT distance="650" swimtime="00:08:12.26" />
                    <SPLIT distance="675" swimtime="00:08:31.89" />
                    <SPLIT distance="700" swimtime="00:08:51.83" />
                    <SPLIT distance="725" swimtime="00:09:11.29" />
                    <SPLIT distance="750" swimtime="00:09:31.18" />
                    <SPLIT distance="775" swimtime="00:09:50.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="467" swimtime="00:00:57.89" resultid="107555" heatid="110688" lane="9" entrytime="00:00:58.84">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.47" />
                    <SPLIT distance="50" swimtime="00:00:28.01" />
                    <SPLIT distance="75" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="416" reactiontime="+94" swimtime="00:01:07.84" resultid="107556" heatid="110704" lane="3" entrytime="00:01:07.86">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="75" swimtime="00:00:52.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="424" swimtime="00:00:29.00" resultid="107557" heatid="110749" lane="9" entrytime="00:00:29.36">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="450" reactiontime="+79" swimtime="00:02:09.65" resultid="107558" heatid="110776" lane="4" entrytime="00:02:12.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                    <SPLIT distance="75" swimtime="00:00:44.53" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="125" swimtime="00:01:17.32" />
                    <SPLIT distance="150" swimtime="00:01:34.61" />
                    <SPLIT distance="175" swimtime="00:01:52.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="384" reactiontime="+83" swimtime="00:01:06.64" resultid="107559" heatid="110803" lane="7" entrytime="00:01:09.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.32" />
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="75" swimtime="00:00:48.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="395" swimtime="00:04:49.27" resultid="107560" heatid="110844" lane="9" entrytime="00:04:53.16">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.14" />
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="75" swimtime="00:00:49.43" />
                    <SPLIT distance="100" swimtime="00:01:07.27" />
                    <SPLIT distance="125" swimtime="00:01:25.39" />
                    <SPLIT distance="150" swimtime="00:01:43.47" />
                    <SPLIT distance="175" swimtime="00:02:02.07" />
                    <SPLIT distance="200" swimtime="00:02:21.00" />
                    <SPLIT distance="225" swimtime="00:02:39.57" />
                    <SPLIT distance="250" swimtime="00:02:58.43" />
                    <SPLIT distance="275" swimtime="00:03:17.29" />
                    <SPLIT distance="300" swimtime="00:03:36.16" />
                    <SPLIT distance="325" swimtime="00:03:55.01" />
                    <SPLIT distance="350" swimtime="00:04:13.75" />
                    <SPLIT distance="375" swimtime="00:04:32.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="429" reactiontime="+65" swimtime="00:01:59.97" resultid="107632" heatid="110719" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.39" />
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="75" swimtime="00:00:46.14" />
                    <SPLIT distance="100" swimtime="00:01:04.53" />
                    <SPLIT distance="125" swimtime="00:01:17.85" />
                    <SPLIT distance="150" swimtime="00:01:33.68" />
                    <SPLIT distance="175" swimtime="00:01:46.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107561" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="107607" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="107569" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="107552" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="324" reactiontime="+71" swimtime="00:02:11.72" resultid="107633" heatid="110718" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="75" swimtime="00:00:53.67" />
                    <SPLIT distance="100" swimtime="00:01:15.94" />
                    <SPLIT distance="125" swimtime="00:01:28.55" />
                    <SPLIT distance="150" swimtime="00:01:44.46" />
                    <SPLIT distance="175" swimtime="00:01:57.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107614" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="107624" number="2" />
                    <RELAYPOSITION athleteid="107628" number="3" />
                    <RELAYPOSITION athleteid="107597" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="99059" status="WDR" swimtime="00:00:00.00" resultid="107634" heatid="110717" lane="3" entrytime="00:02:16.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107614" number="1" />
                    <RELAYPOSITION athleteid="107574" number="2" />
                    <RELAYPOSITION athleteid="107628" number="3" />
                    <RELAYPOSITION athleteid="107579" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="99250" points="475" reactiontime="+94" swimtime="00:01:45.82" resultid="107635" heatid="110784" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.63" />
                    <SPLIT distance="50" swimtime="00:00:26.34" />
                    <SPLIT distance="75" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:00:53.18" />
                    <SPLIT distance="125" swimtime="00:01:05.67" />
                    <SPLIT distance="150" swimtime="00:01:19.19" />
                    <SPLIT distance="175" swimtime="00:01:32.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107628" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="107552" number="2" reactiontime="+14" />
                    <RELAYPOSITION athleteid="107569" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="107597" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="99250" points="415" reactiontime="+86" swimtime="00:01:50.71" resultid="107636" heatid="110783" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.17" />
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                    <SPLIT distance="75" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:00:53.75" />
                    <SPLIT distance="125" swimtime="00:01:06.85" />
                    <SPLIT distance="150" swimtime="00:01:21.08" />
                    <SPLIT distance="175" swimtime="00:01:34.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107607" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="107561" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="107588" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="107614" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="99250" status="WDR" swimtime="00:00:00.00" resultid="107637" heatid="110782" lane="6" entrytime="00:02:08.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107579" number="1" />
                    <RELAYPOSITION athleteid="107614" number="2" />
                    <RELAYPOSITION athleteid="107624" number="3" />
                    <RELAYPOSITION athleteid="107602" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MASTKRASNI" nation="POL" region="LU" clubid="108239" name="Masterskrasnik">
          <CONTACT city="Kraśnik" email="masterskrasnik@gmail.com" internet="www.masterskrasnik.za.pl" name="Michalczyk Jerzy" phone="601698977" state="LUB." street="Żwirki i Wigury 2" zip="23-203" />
          <ATHLETES>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="108240">
              <RESULTS>
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="108241" heatid="110653" lane="8" entrytime="00:00:49.20" />
                <RESULT eventid="98988" points="111" swimtime="00:01:45.22" resultid="108242" heatid="110697" lane="0" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.76" />
                    <SPLIT distance="50" swimtime="00:00:48.88" />
                    <SPLIT distance="75" swimtime="00:01:20.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="89" reactiontime="+88" swimtime="00:00:48.69" resultid="108243" heatid="110742" lane="7" entrytime="00:00:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="91" reactiontime="+99" swimtime="00:01:48.73" resultid="108244" heatid="110758" lane="3" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.65" />
                    <SPLIT distance="50" swimtime="00:00:52.60" />
                    <SPLIT distance="75" swimtime="00:01:22.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="94" reactiontime="+112" swimtime="00:03:52.16" resultid="108245" heatid="110811" lane="7" entrytime="00:04:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.85" />
                    <SPLIT distance="50" swimtime="00:00:54.54" />
                    <SPLIT distance="75" swimtime="00:01:24.30" />
                    <SPLIT distance="100" swimtime="00:01:55.41" />
                    <SPLIT distance="125" swimtime="00:02:25.97" />
                    <SPLIT distance="150" swimtime="00:02:56.50" />
                    <SPLIT distance="175" swimtime="00:03:26.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="108246" heatid="110825" lane="8" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="108258">
              <RESULTS>
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="108259" heatid="110652" lane="9" entrytime="00:00:57.00" />
                <RESULT eventid="106277" points="102" reactiontime="+94" swimtime="00:01:36.06" resultid="108260" heatid="110679" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.37" />
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                    <SPLIT distance="75" swimtime="00:01:10.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="112" reactiontime="+98" swimtime="00:01:55.31" resultid="108261" heatid="110727" lane="4" entrytime="00:01:57.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.22" />
                    <SPLIT distance="50" swimtime="00:00:55.07" />
                    <SPLIT distance="75" swimtime="00:01:25.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="92" reactiontime="+103" swimtime="00:00:48.29" resultid="108262" heatid="110742" lane="1" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="72" reactiontime="+98" swimtime="00:01:56.37" resultid="108263" heatid="110798" lane="5" entrytime="00:01:59.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.64" />
                    <SPLIT distance="50" swimtime="00:00:52.69" />
                    <SPLIT distance="75" swimtime="00:01:25.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-08-16" firstname="Andrzej" gender="M" lastname="Krawczyk" nation="POL" athleteid="108252">
              <RESULTS>
                <RESULT eventid="98798" points="88" reactiontime="+117" swimtime="00:00:45.51" resultid="108253" heatid="110596" lane="2" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="108254" heatid="110651" lane="4" entrytime="00:00:58.00" />
                <RESULT eventid="106277" points="76" swimtime="00:01:46.03" resultid="108255" heatid="110679" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.41" />
                    <SPLIT distance="50" swimtime="00:00:49.06" />
                    <SPLIT distance="75" swimtime="00:01:16.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="77" swimtime="00:02:10.24" resultid="108256" heatid="110727" lane="6" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.19" />
                    <SPLIT distance="50" swimtime="00:01:00.58" />
                    <SPLIT distance="75" swimtime="00:01:34.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="107" swimtime="00:00:53.03" resultid="108257" heatid="110825" lane="0" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-02-09" firstname="Marcin" gender="M" lastname="Mazurek" nation="POL" athleteid="108247">
              <RESULTS>
                <RESULT eventid="98798" points="198" reactiontime="+94" swimtime="00:00:34.71" resultid="108248" heatid="110602" lane="5" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" reactiontime="+110" status="DNS" swimtime="00:00:00.00" resultid="108249" heatid="110636" lane="1" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.76" />
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="75" swimtime="00:01:02.50" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="125" swimtime="00:01:50.60" />
                    <SPLIT distance="150" swimtime="00:02:15.05" />
                    <SPLIT distance="175" swimtime="00:02:40.18" />
                    <SPLIT distance="200" swimtime="00:03:05.79" />
                    <SPLIT distance="225" swimtime="00:03:31.43" />
                    <SPLIT distance="250" swimtime="00:03:57.44" />
                    <SPLIT distance="275" swimtime="00:04:23.76" />
                    <SPLIT distance="300" swimtime="00:04:50.06" />
                    <SPLIT distance="325" swimtime="00:05:17.10" />
                    <SPLIT distance="350" swimtime="00:05:44.24" />
                    <SPLIT distance="375" swimtime="00:06:11.31" />
                    <SPLIT distance="400" swimtime="00:06:38.02" />
                    <SPLIT distance="425" swimtime="00:07:05.58" />
                    <SPLIT distance="450" swimtime="00:07:33.35" />
                    <SPLIT distance="475" swimtime="00:08:00.85" />
                    <SPLIT distance="500" swimtime="00:08:28.72" />
                    <SPLIT distance="525" swimtime="00:08:56.73" />
                    <SPLIT distance="550" swimtime="00:09:24.70" />
                    <SPLIT distance="575" swimtime="00:09:52.86" />
                    <SPLIT distance="600" swimtime="00:10:20.73" />
                    <SPLIT distance="625" swimtime="00:10:49.15" />
                    <SPLIT distance="650" swimtime="00:11:17.33" />
                    <SPLIT distance="675" swimtime="00:11:46.30" />
                    <SPLIT distance="700" swimtime="00:12:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="170" reactiontime="+119" swimtime="00:02:59.20" resultid="108250" heatid="110772" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.41" />
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="75" swimtime="00:01:01.14" />
                    <SPLIT distance="100" swimtime="00:01:24.02" />
                    <SPLIT distance="125" swimtime="00:01:47.84" />
                    <SPLIT distance="150" swimtime="00:02:11.88" />
                    <SPLIT distance="175" swimtime="00:02:36.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="159" swimtime="00:06:31.73" resultid="108251" heatid="110850" lane="0" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.32" />
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="75" swimtime="00:01:05.77" />
                    <SPLIT distance="100" swimtime="00:01:29.30" />
                    <SPLIT distance="125" swimtime="00:01:52.95" />
                    <SPLIT distance="150" swimtime="00:02:17.47" />
                    <SPLIT distance="175" swimtime="00:02:42.34" />
                    <SPLIT distance="200" swimtime="00:03:07.14" />
                    <SPLIT distance="225" swimtime="00:03:31.91" />
                    <SPLIT distance="250" swimtime="00:03:57.40" />
                    <SPLIT distance="275" swimtime="00:04:23.39" />
                    <SPLIT distance="300" swimtime="00:04:49.28" />
                    <SPLIT distance="325" swimtime="00:05:15.16" />
                    <SPLIT distance="350" swimtime="00:05:40.86" />
                    <SPLIT distance="375" swimtime="00:06:07.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="109128" name="MCSiR Płońsk">
          <ATHLETES>
            <ATHLETE birthdate="1940-01-01" firstname="ALINA" gender="F" lastname="Wieczorkiewicz" nation="POL" athleteid="109129">
              <RESULTS>
                <RESULT eventid="98777" points="16" swimtime="00:01:30.46" resultid="109130" heatid="110585" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="21" reactiontime="+110" swimtime="00:01:32.47" resultid="109131" heatid="110646" lane="0" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:44.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="19" reactiontime="+150" swimtime="00:03:31.97" resultid="109132" heatid="110690" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:53.37" />
                    <SPLIT distance="50" swimtime="00:01:43.77" />
                    <SPLIT distance="75" swimtime="00:02:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="11" reactiontime="+114" swimtime="00:01:47.14" resultid="109133" heatid="110735" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="22" reactiontime="+98" swimtime="00:03:15.70" resultid="109134" heatid="110753" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:46.32" />
                    <SPLIT distance="50" swimtime="00:01:36.41" />
                    <SPLIT distance="75" swimtime="00:02:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="23" reactiontime="+106" swimtime="00:06:59.23" resultid="109135" heatid="110806" lane="7" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:47.15" />
                    <SPLIT distance="50" swimtime="00:01:37.34" />
                    <SPLIT distance="75" swimtime="00:02:27.44" />
                    <SPLIT distance="100" swimtime="00:03:21.42" />
                    <SPLIT distance="125" swimtime="00:04:15.95" />
                    <SPLIT distance="150" swimtime="00:05:11.69" />
                    <SPLIT distance="175" swimtime="00:06:05.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00308" nation="POL" region="PDK" clubid="107638" name="MKP Bobry Dębica">
          <CONTACT email="goben@interia.pl" name="GOGACZ" phone="506694816" />
          <ATHLETES>
            <ATHLETE birthdate="1991-10-29" firstname="Marcin" gender="M" lastname="Potoczny" nation="POL" athleteid="107676">
              <RESULTS>
                <RESULT eventid="98798" points="158" reactiontime="+86" swimtime="00:00:37.40" resultid="107677" heatid="110598" lane="8" entrytime="00:00:38.97">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="99" reactiontime="+90" swimtime="00:00:48.03" resultid="107678" heatid="110653" lane="1" entrytime="00:00:47.61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="138" swimtime="00:01:26.88" resultid="107679" heatid="110680" lane="9" entrytime="00:01:28.94">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.01" />
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                    <SPLIT distance="75" swimtime="00:01:04.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="100" reactiontime="+94" swimtime="00:01:45.20" resultid="107680" heatid="110757" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.76" />
                    <SPLIT distance="50" swimtime="00:00:51.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="131" reactiontime="+95" swimtime="00:03:15.31" resultid="107681" heatid="110770" lane="7" entrytime="00:03:23.41">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.62" />
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                    <SPLIT distance="75" swimtime="00:01:06.66" />
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                    <SPLIT distance="125" swimtime="00:01:58.00" />
                    <SPLIT distance="150" swimtime="00:02:23.98" />
                    <SPLIT distance="175" swimtime="00:02:49.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="118" reactiontime="+89" swimtime="00:07:12.16" resultid="107682" heatid="110851" lane="5" entrytime="00:07:18.62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.53" />
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                    <SPLIT distance="75" swimtime="00:01:09.05" />
                    <SPLIT distance="100" swimtime="00:01:35.57" />
                    <SPLIT distance="125" swimtime="00:02:02.95" />
                    <SPLIT distance="150" swimtime="00:02:30.51" />
                    <SPLIT distance="175" swimtime="00:02:58.24" />
                    <SPLIT distance="200" swimtime="00:03:26.68" />
                    <SPLIT distance="225" swimtime="00:03:54.96" />
                    <SPLIT distance="250" swimtime="00:04:23.36" />
                    <SPLIT distance="275" swimtime="00:04:51.66" />
                    <SPLIT distance="300" swimtime="00:05:20.32" />
                    <SPLIT distance="325" swimtime="00:05:48.94" />
                    <SPLIT distance="350" swimtime="00:06:17.11" />
                    <SPLIT distance="375" swimtime="00:06:45.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-12" firstname="Katarzyna" gender="F" lastname="Walkowicz" nation="POL" license="500308600144" athleteid="107671">
              <RESULTS>
                <RESULT eventid="98777" points="466" reactiontime="+77" swimtime="00:00:29.96" resultid="107672" heatid="110592" lane="7" entrytime="00:00:29.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="465" reactiontime="+83" swimtime="00:02:53.63" resultid="107673" heatid="110664" lane="4" entrytime="00:02:48.79">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.05" />
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="75" swimtime="00:01:00.32" />
                    <SPLIT distance="100" swimtime="00:01:22.66" />
                    <SPLIT distance="125" swimtime="00:01:45.29" />
                    <SPLIT distance="150" swimtime="00:02:08.27" />
                    <SPLIT distance="175" swimtime="00:02:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="498" reactiontime="+84" swimtime="00:01:18.66" resultid="107674" heatid="110725" lane="5" entrytime="00:01:19.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.11" />
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="75" swimtime="00:00:57.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="520" reactiontime="+82" swimtime="00:00:35.81" resultid="107675" heatid="110823" lane="1" entrytime="00:00:36.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-11" firstname="Przemysław" gender="M" lastname="Jurek" nation="POL" license="100308700118" athleteid="107662">
              <RESULTS>
                <RESULT eventid="98798" points="502" reactiontime="+92" swimtime="00:00:25.48" resultid="107663" heatid="110612" lane="2" entrytime="00:00:24.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="452" swimtime="00:02:22.79" resultid="107664" heatid="110628" lane="9" entrytime="00:02:23.46">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                    <SPLIT distance="75" swimtime="00:00:46.98" />
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                    <SPLIT distance="125" swimtime="00:01:26.53" />
                    <SPLIT distance="150" swimtime="00:01:48.94" />
                    <SPLIT distance="175" swimtime="00:02:06.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="551" reactiontime="+88" swimtime="00:00:54.79" resultid="107665" heatid="110689" lane="7" entrytime="00:00:55.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                    <SPLIT distance="75" swimtime="00:00:41.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="550" reactiontime="+86" swimtime="00:01:01.82" resultid="107666" heatid="110706" lane="7" entrytime="00:01:02.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.60" />
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                    <SPLIT distance="75" swimtime="00:00:46.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="499" swimtime="00:00:27.48" resultid="107667" heatid="110750" lane="0" entrytime="00:00:27.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="530" reactiontime="+92" swimtime="00:02:02.76" resultid="107668" heatid="110778" lane="1" entrytime="00:01:59.81">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.39" />
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                    <SPLIT distance="75" swimtime="00:00:44.04" />
                    <SPLIT distance="100" swimtime="00:00:59.69" />
                    <SPLIT distance="125" swimtime="00:01:15.41" />
                    <SPLIT distance="150" swimtime="00:01:31.47" />
                    <SPLIT distance="175" swimtime="00:01:47.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="507" swimtime="00:01:00.72" resultid="107669" heatid="110805" lane="0" entrytime="00:00:59.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.64" />
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                    <SPLIT distance="75" swimtime="00:00:44.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="451" swimtime="00:00:32.92" resultid="107670" heatid="110832" lane="2" entrytime="00:00:34.73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" region="ZAC" clubid="108190" name="MKP Szczecin">
          <CONTACT email="windmuhle@wp.pl" name="Kowalczyk Piotr" phone="509758055" />
          <ATHLETES>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="108195">
              <RESULTS>
                <RESULT eventid="106254" points="401" reactiontime="+85" swimtime="00:20:46.28" resultid="108196" heatid="110640" lane="4" entrytime="00:20:52.22">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.79" />
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="75" swimtime="00:00:54.65" />
                    <SPLIT distance="100" swimtime="00:01:14.45" />
                    <SPLIT distance="125" swimtime="00:01:34.62" />
                    <SPLIT distance="150" swimtime="00:01:54.93" />
                    <SPLIT distance="175" swimtime="00:02:15.36" />
                    <SPLIT distance="200" swimtime="00:02:35.89" />
                    <SPLIT distance="225" swimtime="00:02:56.40" />
                    <SPLIT distance="250" swimtime="00:03:17.05" />
                    <SPLIT distance="275" swimtime="00:03:37.70" />
                    <SPLIT distance="300" swimtime="00:03:58.38" />
                    <SPLIT distance="325" swimtime="00:04:19.23" />
                    <SPLIT distance="350" swimtime="00:04:40.01" />
                    <SPLIT distance="375" swimtime="00:05:00.85" />
                    <SPLIT distance="400" swimtime="00:05:21.65" />
                    <SPLIT distance="425" swimtime="00:05:42.50" />
                    <SPLIT distance="450" swimtime="00:06:03.11" />
                    <SPLIT distance="475" swimtime="00:06:23.78" />
                    <SPLIT distance="500" swimtime="00:06:44.39" />
                    <SPLIT distance="525" swimtime="00:07:05.12" />
                    <SPLIT distance="550" swimtime="00:07:25.88" />
                    <SPLIT distance="575" swimtime="00:07:46.73" />
                    <SPLIT distance="600" swimtime="00:08:07.51" />
                    <SPLIT distance="625" swimtime="00:08:28.30" />
                    <SPLIT distance="650" swimtime="00:08:49.03" />
                    <SPLIT distance="675" swimtime="00:09:09.77" />
                    <SPLIT distance="700" swimtime="00:09:30.59" />
                    <SPLIT distance="725" swimtime="00:09:51.43" />
                    <SPLIT distance="750" swimtime="00:10:12.22" />
                    <SPLIT distance="775" swimtime="00:10:33.18" />
                    <SPLIT distance="800" swimtime="00:10:54.16" />
                    <SPLIT distance="825" swimtime="00:11:15.00" />
                    <SPLIT distance="850" swimtime="00:11:35.98" />
                    <SPLIT distance="875" swimtime="00:11:56.97" />
                    <SPLIT distance="900" swimtime="00:12:18.07" />
                    <SPLIT distance="925" swimtime="00:12:39.30" />
                    <SPLIT distance="950" swimtime="00:13:00.35" />
                    <SPLIT distance="975" swimtime="00:13:21.45" />
                    <SPLIT distance="1000" swimtime="00:13:42.52" />
                    <SPLIT distance="1025" swimtime="00:14:03.73" />
                    <SPLIT distance="1050" swimtime="00:14:24.71" />
                    <SPLIT distance="1075" swimtime="00:14:45.90" />
                    <SPLIT distance="1100" swimtime="00:15:07.16" />
                    <SPLIT distance="1125" swimtime="00:15:28.41" />
                    <SPLIT distance="1150" swimtime="00:15:49.54" />
                    <SPLIT distance="1175" swimtime="00:16:10.72" />
                    <SPLIT distance="1200" swimtime="00:16:31.81" />
                    <SPLIT distance="1225" swimtime="00:16:53.04" />
                    <SPLIT distance="1250" swimtime="00:17:14.21" />
                    <SPLIT distance="1275" swimtime="00:17:35.66" />
                    <SPLIT distance="1300" swimtime="00:17:56.92" />
                    <SPLIT distance="1325" swimtime="00:18:18.31" />
                    <SPLIT distance="1350" swimtime="00:18:39.53" />
                    <SPLIT distance="1375" swimtime="00:19:00.96" />
                    <SPLIT distance="1400" swimtime="00:19:22.25" />
                    <SPLIT distance="1425" swimtime="00:19:43.50" />
                    <SPLIT distance="1450" swimtime="00:20:04.66" />
                    <SPLIT distance="1475" swimtime="00:20:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="394" swimtime="00:02:31.04" resultid="108197" heatid="110768" lane="9" entrytime="00:02:29.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.42" />
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="75" swimtime="00:00:53.74" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="125" swimtime="00:01:33.08" />
                    <SPLIT distance="150" swimtime="00:01:52.74" />
                    <SPLIT distance="175" swimtime="00:02:12.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="326" reactiontime="+95" swimtime="00:02:53.12" resultid="108198" heatid="110809" lane="2" entrytime="00:02:51.05">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.37" />
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="75" swimtime="00:01:03.46" />
                    <SPLIT distance="100" swimtime="00:01:25.38" />
                    <SPLIT distance="125" swimtime="00:01:47.38" />
                    <SPLIT distance="150" swimtime="00:02:09.78" />
                    <SPLIT distance="175" swimtime="00:02:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="399" reactiontime="+90" swimtime="00:05:18.53" resultid="108199" heatid="110839" lane="1" entrytime="00:05:13.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.84" />
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="75" swimtime="00:00:55.09" />
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                    <SPLIT distance="125" swimtime="00:01:35.03" />
                    <SPLIT distance="150" swimtime="00:01:55.21" />
                    <SPLIT distance="175" swimtime="00:02:15.35" />
                    <SPLIT distance="200" swimtime="00:02:35.60" />
                    <SPLIT distance="225" swimtime="00:02:55.89" />
                    <SPLIT distance="250" swimtime="00:03:16.54" />
                    <SPLIT distance="275" swimtime="00:03:37.00" />
                    <SPLIT distance="300" swimtime="00:03:57.57" />
                    <SPLIT distance="325" swimtime="00:04:17.83" />
                    <SPLIT distance="350" swimtime="00:04:38.48" />
                    <SPLIT distance="375" swimtime="00:04:58.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="108200">
              <RESULTS>
                <RESULT eventid="98830" points="177" reactiontime="+103" swimtime="00:03:15.20" resultid="108201" heatid="110621" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.52" />
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="75" swimtime="00:01:06.57" />
                    <SPLIT distance="100" swimtime="00:01:31.82" />
                    <SPLIT distance="125" swimtime="00:01:58.72" />
                    <SPLIT distance="150" swimtime="00:02:26.53" />
                    <SPLIT distance="175" swimtime="00:02:52.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="197" reactiontime="+92" swimtime="00:03:26.76" resultid="108202" heatid="110666" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.42" />
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                    <SPLIT distance="75" swimtime="00:01:13.29" />
                    <SPLIT distance="100" swimtime="00:01:40.35" />
                    <SPLIT distance="125" swimtime="00:02:06.93" />
                    <SPLIT distance="150" swimtime="00:02:33.70" />
                    <SPLIT distance="175" swimtime="00:03:00.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="228" reactiontime="+81" swimtime="00:01:31.01" resultid="108203" heatid="110729" lane="5" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.56" />
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="75" swimtime="00:01:06.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="262" reactiontime="+68" swimtime="00:00:39.42" resultid="108204" heatid="110827" lane="7" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-07-26" firstname="Marcin" gender="M" lastname="Gargas" nation="POL" athleteid="108211">
              <RESULTS>
                <RESULT eventid="98798" points="194" reactiontime="+93" swimtime="00:00:34.95" resultid="108212" heatid="110599" lane="2" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-06" firstname="Lech" gender="M" lastname="Orecki" nation="POL" athleteid="108205">
              <RESULTS>
                <RESULT eventid="98798" points="301" reactiontime="+96" swimtime="00:00:30.21" resultid="108206" heatid="110602" lane="4" entrytime="00:00:30.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="265" reactiontime="+110" swimtime="00:11:29.90" resultid="108207" heatid="110637" lane="3" entrytime="00:11:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.02" />
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="75" swimtime="00:00:57.24" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="125" swimtime="00:01:39.34" />
                    <SPLIT distance="150" swimtime="00:02:01.48" />
                    <SPLIT distance="175" swimtime="00:02:23.79" />
                    <SPLIT distance="200" swimtime="00:02:46.33" />
                    <SPLIT distance="225" swimtime="00:03:08.22" />
                    <SPLIT distance="250" swimtime="00:03:30.65" />
                    <SPLIT distance="275" swimtime="00:03:53.03" />
                    <SPLIT distance="300" swimtime="00:04:15.18" />
                    <SPLIT distance="325" swimtime="00:04:37.33" />
                    <SPLIT distance="350" swimtime="00:04:59.48" />
                    <SPLIT distance="375" swimtime="00:05:21.40" />
                    <SPLIT distance="400" swimtime="00:05:42.65" />
                    <SPLIT distance="425" swimtime="00:06:04.54" />
                    <SPLIT distance="450" swimtime="00:06:26.68" />
                    <SPLIT distance="475" swimtime="00:06:48.49" />
                    <SPLIT distance="500" swimtime="00:07:10.49" />
                    <SPLIT distance="525" swimtime="00:07:31.98" />
                    <SPLIT distance="550" swimtime="00:07:53.77" />
                    <SPLIT distance="575" swimtime="00:08:15.48" />
                    <SPLIT distance="600" swimtime="00:08:37.45" />
                    <SPLIT distance="625" swimtime="00:08:58.98" />
                    <SPLIT distance="650" swimtime="00:09:21.82" />
                    <SPLIT distance="675" swimtime="00:09:44.08" />
                    <SPLIT distance="700" swimtime="00:10:06.13" />
                    <SPLIT distance="725" swimtime="00:10:28.04" />
                    <SPLIT distance="750" swimtime="00:10:50.09" />
                    <SPLIT distance="775" swimtime="00:11:10.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="299" reactiontime="+105" swimtime="00:01:07.15" resultid="108208" heatid="110682" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.49" />
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="75" swimtime="00:00:50.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="297" reactiontime="+101" swimtime="00:02:28.83" resultid="108209" heatid="110772" lane="3" entrytime="00:02:41.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.45" />
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="75" swimtime="00:00:52.23" />
                    <SPLIT distance="100" swimtime="00:01:11.41" />
                    <SPLIT distance="125" swimtime="00:01:31.32" />
                    <SPLIT distance="150" swimtime="00:01:51.23" />
                    <SPLIT distance="175" swimtime="00:02:10.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="275" swimtime="00:05:26.19" resultid="108210" heatid="110848" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.50" />
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="75" swimtime="00:00:55.87" />
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                    <SPLIT distance="125" swimtime="00:01:37.59" />
                    <SPLIT distance="150" swimtime="00:01:59.25" />
                    <SPLIT distance="175" swimtime="00:02:20.36" />
                    <SPLIT distance="200" swimtime="00:02:41.69" />
                    <SPLIT distance="225" swimtime="00:03:02.83" />
                    <SPLIT distance="250" swimtime="00:03:24.24" />
                    <SPLIT distance="275" swimtime="00:03:45.49" />
                    <SPLIT distance="300" swimtime="00:04:07.10" />
                    <SPLIT distance="325" swimtime="00:04:27.96" />
                    <SPLIT distance="350" swimtime="00:04:48.58" />
                    <SPLIT distance="375" swimtime="00:05:08.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-08-21" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="108191">
              <RESULTS>
                <RESULT eventid="98940" points="90" swimtime="00:04:59.68" resultid="108192" heatid="110661" lane="6" entrytime="00:04:58.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.83" />
                    <SPLIT distance="50" swimtime="00:01:10.82" />
                    <SPLIT distance="75" swimtime="00:01:48.33" />
                    <SPLIT distance="100" swimtime="00:02:26.84" />
                    <SPLIT distance="125" swimtime="00:03:05.74" />
                    <SPLIT distance="150" swimtime="00:03:45.41" />
                    <SPLIT distance="175" swimtime="00:04:23.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="86" swimtime="00:02:20.95" resultid="108193" heatid="110721" lane="7" entrytime="00:02:20.46">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.62" />
                    <SPLIT distance="50" swimtime="00:01:09.02" />
                    <SPLIT distance="75" swimtime="00:01:44.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="81" swimtime="00:01:06.50" resultid="108194" heatid="110817" lane="4" entrytime="00:01:08.85">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00816" nation="POL" region="SZ" clubid="107526" name="MKS Neptun Stargard">
          <CONTACT city="Stargard" email="prezes@mksneptun.pl" internet="www.mksneptun.pl" name="Miedzyszkolny Klub Sportowy &quot;Neptun&quot;" phone="602731410" state="ZACHO" street="Os. Zachód B 15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1994-09-30" firstname="Mateusz" gender="M" lastname="Drozd" nation="POL" athleteid="107540">
              <RESULTS>
                <RESULT eventid="98798" points="561" reactiontime="+80" swimtime="00:00:24.56" resultid="107541" heatid="110613" lane="3" entrytime="00:00:23.82">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="565" reactiontime="+78" swimtime="00:02:12.61" resultid="107542" heatid="110628" lane="5" entrytime="00:02:12.41">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.58" />
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                    <SPLIT distance="75" swimtime="00:00:46.46" />
                    <SPLIT distance="100" swimtime="00:01:03.96" />
                    <SPLIT distance="125" swimtime="00:01:23.18" />
                    <SPLIT distance="150" swimtime="00:01:42.28" />
                    <SPLIT distance="175" swimtime="00:01:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="592" reactiontime="+73" swimtime="00:01:00.33" resultid="107543" heatid="110706" lane="5" entrytime="00:01:00.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.06" />
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                    <SPLIT distance="75" swimtime="00:00:45.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="560" swimtime="00:00:26.44" resultid="107544" heatid="110751" lane="9" entrytime="00:00:26.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="614" swimtime="00:01:56.90" resultid="107545" heatid="110778" lane="6" entrytime="00:01:57.42">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                    <SPLIT distance="75" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:00:56.74" />
                    <SPLIT distance="125" swimtime="00:01:11.92" />
                    <SPLIT distance="150" swimtime="00:01:27.20" />
                    <SPLIT distance="175" swimtime="00:01:42.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="471" reactiontime="+83" swimtime="00:02:15.67" resultid="107546" heatid="110816" lane="4" entrytime="00:02:04.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.61" />
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="75" swimtime="00:00:46.91" />
                    <SPLIT distance="100" swimtime="00:01:03.94" />
                    <SPLIT distance="125" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:01:39.77" />
                    <SPLIT distance="175" swimtime="00:01:57.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-08-18" firstname="Ireneusz" gender="M" lastname="Drozd" nation="POL" athleteid="107547">
              <RESULTS>
                <RESULT eventid="98924" points="287" reactiontime="+91" swimtime="00:00:33.65" resultid="107548" heatid="110656" lane="4" entrytime="00:00:34.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="380" reactiontime="+66" swimtime="00:00:30.08" resultid="107549" heatid="110748" lane="2" entrytime="00:00:29.65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="209" reactiontime="+87" swimtime="00:02:57.93" resultid="107550" heatid="110814" lane="1" entrytime="00:02:44.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.27" />
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="75" swimtime="00:00:58.91" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="125" swimtime="00:01:42.54" />
                    <SPLIT distance="150" swimtime="00:02:06.50" />
                    <SPLIT distance="175" swimtime="00:02:33.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWDOL" nation="POL" region="DOL" clubid="108213" name="MKS Swim Academy Termy Jakuba Oława" shortname="MKS Swim Academy Termy Jakuba ">
          <CONTACT city="Oława" email="biuro@swim-academy.pl" internet="www.swim-academy.pl" name="Grzegorz Fidala / Jacek Bereżnicki" phone="601316031 / 69643365" state="DOL" street="1 Maja 33a" zip="55-200" />
          <ATHLETES>
            <ATHLETE birthdate="1991-07-06" firstname="Agnieszka" gender="F" lastname="Burdelak" nation="POL" license="5045016000019" athleteid="108214">
              <RESULTS>
                <RESULT eventid="98777" points="522" reactiontime="+79" swimtime="00:00:28.85" resultid="108215" heatid="110592" lane="4" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="460" swimtime="00:02:37.84" resultid="108216" heatid="110618" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.94" />
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="75" swimtime="00:00:55.29" />
                    <SPLIT distance="100" swimtime="00:01:16.60" />
                    <SPLIT distance="125" swimtime="00:01:38.83" />
                    <SPLIT distance="150" swimtime="00:02:01.15" />
                    <SPLIT distance="175" swimtime="00:02:19.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="464" reactiontime="+70" swimtime="00:02:53.74" resultid="108217" heatid="110664" lane="5" entrytime="00:02:52.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.76" />
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="75" swimtime="00:01:01.24" />
                    <SPLIT distance="100" swimtime="00:01:23.29" />
                    <SPLIT distance="125" swimtime="00:01:45.74" />
                    <SPLIT distance="150" swimtime="00:02:08.48" />
                    <SPLIT distance="175" swimtime="00:02:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="488" reactiontime="+69" swimtime="00:01:11.98" resultid="108218" heatid="110695" lane="6" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.63" />
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="75" swimtime="00:00:54.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="488" reactiontime="+60" swimtime="00:01:19.18" resultid="108219" heatid="110725" lane="2" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.29" />
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="75" swimtime="00:00:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="435" reactiontime="+63" swimtime="00:01:12.62" resultid="108220" heatid="110756" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.09" />
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="75" swimtime="00:00:53.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="386" reactiontime="+77" swimtime="00:01:14.97" resultid="108221" heatid="110796" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.56" />
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="75" swimtime="00:00:53.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="501" swimtime="00:00:36.24" resultid="108222" heatid="110823" lane="2" entrytime="00:00:36.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="107769" name="MOSiR KSZO Ostrowiec Św.">
          <CONTACT name="Różalski Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" athleteid="107770">
              <RESULTS>
                <RESULT eventid="98798" points="234" reactiontime="+85" swimtime="00:00:32.87" resultid="107771" heatid="110599" lane="8" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="143" reactiontime="+105" swimtime="00:03:29.56" resultid="107772" heatid="110620" lane="1" entrytime="00:03:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.26" />
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                    <SPLIT distance="75" swimtime="00:01:14.29" />
                    <SPLIT distance="100" swimtime="00:01:44.44" />
                    <SPLIT distance="125" swimtime="00:02:15.06" />
                    <SPLIT distance="150" swimtime="00:02:45.74" />
                    <SPLIT distance="175" swimtime="00:03:08.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="144" reactiontime="+101" swimtime="00:03:49.68" resultid="107773" heatid="110666" lane="1" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.62" />
                    <SPLIT distance="50" swimtime="00:00:49.92" />
                    <SPLIT distance="75" swimtime="00:01:17.72" />
                    <SPLIT distance="100" swimtime="00:01:46.28" />
                    <SPLIT distance="125" swimtime="00:02:16.34" />
                    <SPLIT distance="150" swimtime="00:02:47.58" />
                    <SPLIT distance="175" swimtime="00:03:18.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="170" reactiontime="+101" swimtime="00:01:31.36" resultid="107774" heatid="110697" lane="2" entrytime="00:01:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.52" />
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                    <SPLIT distance="75" swimtime="00:01:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="171" reactiontime="+94" swimtime="00:01:40.16" resultid="107775" heatid="110728" lane="7" entrytime="00:01:45.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.45" />
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                    <SPLIT distance="75" swimtime="00:01:13.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="194" swimtime="00:00:37.64" resultid="107776" heatid="110743" lane="0" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="114" reactiontime="+125" swimtime="00:01:39.77" resultid="107777" heatid="110799" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.18" />
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                    <SPLIT distance="75" swimtime="00:01:12.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="161" reactiontime="+104" swimtime="00:00:46.39" resultid="107778" heatid="110825" lane="3" entrytime="00:00:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="106396" name="MOSIR MIELEC">
          <ATHLETES>
            <ATHLETE birthdate="1988-01-01" firstname="DANIEL" gender="M" lastname="PADUCH " nation="POL" athleteid="106397">
              <RESULTS>
                <RESULT eventid="106256" points="470" reactiontime="+74" swimtime="00:18:10.27" resultid="106398" heatid="110641" lane="5" entrytime="00:18:21.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.60" />
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="75" swimtime="00:00:48.66" />
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                    <SPLIT distance="125" swimtime="00:01:24.11" />
                    <SPLIT distance="150" swimtime="00:01:41.80" />
                    <SPLIT distance="175" swimtime="00:01:59.82" />
                    <SPLIT distance="200" swimtime="00:02:17.63" />
                    <SPLIT distance="225" swimtime="00:02:35.63" />
                    <SPLIT distance="250" swimtime="00:02:53.69" />
                    <SPLIT distance="275" swimtime="00:03:11.83" />
                    <SPLIT distance="300" swimtime="00:03:30.09" />
                    <SPLIT distance="325" swimtime="00:03:48.28" />
                    <SPLIT distance="350" swimtime="00:04:06.38" />
                    <SPLIT distance="375" swimtime="00:04:24.52" />
                    <SPLIT distance="400" swimtime="00:04:43.42" />
                    <SPLIT distance="425" swimtime="00:05:01.68" />
                    <SPLIT distance="450" swimtime="00:05:19.77" />
                    <SPLIT distance="475" swimtime="00:05:38.45" />
                    <SPLIT distance="500" swimtime="00:05:56.90" />
                    <SPLIT distance="525" swimtime="00:06:15.39" />
                    <SPLIT distance="550" swimtime="00:06:33.72" />
                    <SPLIT distance="575" swimtime="00:06:51.90" />
                    <SPLIT distance="600" swimtime="00:07:10.92" />
                    <SPLIT distance="625" swimtime="00:07:29.05" />
                    <SPLIT distance="650" swimtime="00:07:47.35" />
                    <SPLIT distance="675" swimtime="00:08:05.85" />
                    <SPLIT distance="700" swimtime="00:08:24.39" />
                    <SPLIT distance="725" swimtime="00:08:43.47" />
                    <SPLIT distance="750" swimtime="00:09:02.47" />
                    <SPLIT distance="775" swimtime="00:09:21.26" />
                    <SPLIT distance="800" swimtime="00:09:39.85" />
                    <SPLIT distance="825" swimtime="00:09:58.30" />
                    <SPLIT distance="850" swimtime="00:10:16.88" />
                    <SPLIT distance="875" swimtime="00:10:35.51" />
                    <SPLIT distance="900" swimtime="00:10:53.74" />
                    <SPLIT distance="925" swimtime="00:11:12.26" />
                    <SPLIT distance="950" swimtime="00:11:30.81" />
                    <SPLIT distance="975" swimtime="00:11:49.28" />
                    <SPLIT distance="1000" swimtime="00:12:08.13" />
                    <SPLIT distance="1025" swimtime="00:12:26.49" />
                    <SPLIT distance="1050" swimtime="00:12:45.09" />
                    <SPLIT distance="1075" swimtime="00:13:03.29" />
                    <SPLIT distance="1100" swimtime="00:13:22.05" />
                    <SPLIT distance="1125" swimtime="00:13:40.34" />
                    <SPLIT distance="1150" swimtime="00:13:58.33" />
                    <SPLIT distance="1175" swimtime="00:14:16.25" />
                    <SPLIT distance="1200" swimtime="00:14:34.14" />
                    <SPLIT distance="1225" swimtime="00:14:52.31" />
                    <SPLIT distance="1250" swimtime="00:15:10.53" />
                    <SPLIT distance="1275" swimtime="00:15:28.75" />
                    <SPLIT distance="1300" swimtime="00:15:47.20" />
                    <SPLIT distance="1325" swimtime="00:16:05.01" />
                    <SPLIT distance="1350" swimtime="00:16:23.65" />
                    <SPLIT distance="1375" swimtime="00:16:42.20" />
                    <SPLIT distance="1400" swimtime="00:17:00.29" />
                    <SPLIT distance="1425" swimtime="00:17:17.84" />
                    <SPLIT distance="1450" swimtime="00:17:35.70" />
                    <SPLIT distance="1475" swimtime="00:17:53.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="507" reactiontime="+70" swimtime="00:02:16.06" resultid="106399" heatid="110713" lane="6" entrytime="00:02:16.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.87" />
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="75" swimtime="00:00:47.76" />
                    <SPLIT distance="100" swimtime="00:01:06.50" />
                    <SPLIT distance="125" swimtime="00:01:22.83" />
                    <SPLIT distance="150" swimtime="00:01:40.95" />
                    <SPLIT distance="175" swimtime="00:01:58.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="463" reactiontime="+55" swimtime="00:02:08.43" resultid="106400" heatid="110777" lane="2" entrytime="00:02:09.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.96" />
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="75" swimtime="00:00:46.19" />
                    <SPLIT distance="100" swimtime="00:01:02.95" />
                    <SPLIT distance="125" swimtime="00:01:19.45" />
                    <SPLIT distance="150" swimtime="00:01:36.30" />
                    <SPLIT distance="175" swimtime="00:01:52.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="106401" heatid="110792" lane="6" entrytime="00:05:09.98" />
                <RESULT eventid="99473" points="455" swimtime="00:04:35.78" resultid="106402" heatid="110843" lane="6" entrytime="00:04:29.78">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.29" />
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="75" swimtime="00:00:47.67" />
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="125" swimtime="00:01:22.55" />
                    <SPLIT distance="150" swimtime="00:01:40.07" />
                    <SPLIT distance="175" swimtime="00:01:57.55" />
                    <SPLIT distance="200" swimtime="00:02:15.25" />
                    <SPLIT distance="225" swimtime="00:02:32.58" />
                    <SPLIT distance="250" swimtime="00:02:50.38" />
                    <SPLIT distance="275" swimtime="00:03:08.04" />
                    <SPLIT distance="300" swimtime="00:03:25.70" />
                    <SPLIT distance="325" swimtime="00:03:43.71" />
                    <SPLIT distance="350" swimtime="00:04:00.99" />
                    <SPLIT distance="375" swimtime="00:04:18.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" clubid="108396" name="MOTYL-SENIOR MOSiR Stalowa Wola" shortname="MOTYL-SENIOR MOSiR St. Wola">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Niedbałowski Jarosław" state="PODK" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="108430">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="108431" heatid="110589" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="98814" points="265" reactiontime="+109" swimtime="00:03:09.60" resultid="108432" heatid="110616" lane="1" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.60" />
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="75" swimtime="00:01:06.02" />
                    <SPLIT distance="100" swimtime="00:01:31.01" />
                    <SPLIT distance="125" swimtime="00:01:57.53" />
                    <SPLIT distance="150" swimtime="00:02:25.26" />
                    <SPLIT distance="175" swimtime="00:02:47.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="256" reactiontime="+80" swimtime="00:03:31.77" resultid="108433" heatid="110662" lane="4" entrytime="00:03:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.53" />
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                    <SPLIT distance="75" swimtime="00:01:15.63" />
                    <SPLIT distance="100" swimtime="00:01:43.45" />
                    <SPLIT distance="125" swimtime="00:02:11.61" />
                    <SPLIT distance="150" swimtime="00:02:39.49" />
                    <SPLIT distance="175" swimtime="00:03:06.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="279" swimtime="00:01:26.72" resultid="108434" heatid="110692" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.40" />
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="75" swimtime="00:01:06.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="250" swimtime="00:01:38.93" resultid="108435" heatid="110723" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.29" />
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                    <SPLIT distance="75" swimtime="00:01:12.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="251" swimtime="00:00:38.62" resultid="108436" heatid="110738" lane="0" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="194" swimtime="00:01:34.23" resultid="108437" heatid="110794" lane="3" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.37" />
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="75" swimtime="00:01:09.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="274" swimtime="00:00:44.34" resultid="108438" heatid="110820" lane="6" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-12" firstname="Adam" gender="M" lastname="Przybylski" nation="POL" athleteid="108422">
              <RESULTS>
                <RESULT eventid="98798" points="398" reactiontime="+85" swimtime="00:00:27.53" resultid="108423" heatid="110608" lane="7" entrytime="00:00:27.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="246" reactiontime="+70" swimtime="00:00:35.45" resultid="108424" heatid="110656" lane="3" entrytime="00:00:34.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="108425" heatid="110712" lane="0" entrytime="00:03:01.48" />
                <RESULT comment="o4" eventid="99170" status="DSQ" swimtime="00:00:00.00" resultid="108426" heatid="110748" lane="9" entrytime="00:00:30.99" />
                <RESULT eventid="99186" points="248" reactiontime="+90" swimtime="00:01:17.80" resultid="108427" heatid="110761" lane="1" entrytime="00:01:15.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.26" />
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                    <SPLIT distance="75" swimtime="00:00:57.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="108428" heatid="110802" lane="0" entrytime="00:01:14.48" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="108429" heatid="110814" lane="9" entrytime="00:02:48.48" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="108406">
              <RESULTS>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="108407" heatid="110625" lane="9" entrytime="00:02:42.83" />
                <RESULT eventid="106256" points="287" reactiontime="+85" swimtime="00:21:24.80" resultid="108408" heatid="110642" lane="5" entrytime="00:21:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.64" />
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="75" swimtime="00:00:54.28" />
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="125" swimtime="00:01:33.50" />
                    <SPLIT distance="150" swimtime="00:01:53.62" />
                    <SPLIT distance="175" swimtime="00:02:13.92" />
                    <SPLIT distance="200" swimtime="00:02:34.21" />
                    <SPLIT distance="225" swimtime="00:02:54.58" />
                    <SPLIT distance="250" swimtime="00:03:15.05" />
                    <SPLIT distance="275" swimtime="00:03:35.89" />
                    <SPLIT distance="300" swimtime="00:03:56.55" />
                    <SPLIT distance="325" swimtime="00:04:17.57" />
                    <SPLIT distance="350" swimtime="00:04:38.59" />
                    <SPLIT distance="375" swimtime="00:04:59.99" />
                    <SPLIT distance="400" swimtime="00:05:21.12" />
                    <SPLIT distance="425" swimtime="00:05:42.67" />
                    <SPLIT distance="450" swimtime="00:06:04.20" />
                    <SPLIT distance="475" swimtime="00:06:25.76" />
                    <SPLIT distance="500" swimtime="00:06:47.04" />
                    <SPLIT distance="525" swimtime="00:07:08.74" />
                    <SPLIT distance="550" swimtime="00:07:30.09" />
                    <SPLIT distance="575" swimtime="00:07:51.94" />
                    <SPLIT distance="600" swimtime="00:08:13.83" />
                    <SPLIT distance="625" swimtime="00:08:35.66" />
                    <SPLIT distance="650" swimtime="00:08:57.52" />
                    <SPLIT distance="675" swimtime="00:09:19.68" />
                    <SPLIT distance="700" swimtime="00:09:41.46" />
                    <SPLIT distance="725" swimtime="00:10:03.16" />
                    <SPLIT distance="750" swimtime="00:10:24.64" />
                    <SPLIT distance="775" swimtime="00:10:46.77" />
                    <SPLIT distance="800" swimtime="00:11:08.61" />
                    <SPLIT distance="825" swimtime="00:11:29.97" />
                    <SPLIT distance="850" swimtime="00:11:51.41" />
                    <SPLIT distance="875" swimtime="00:12:13.18" />
                    <SPLIT distance="900" swimtime="00:12:35.28" />
                    <SPLIT distance="925" swimtime="00:12:57.33" />
                    <SPLIT distance="950" swimtime="00:13:19.37" />
                    <SPLIT distance="975" swimtime="00:13:41.39" />
                    <SPLIT distance="1000" swimtime="00:14:03.44" />
                    <SPLIT distance="1025" swimtime="00:14:25.56" />
                    <SPLIT distance="1050" swimtime="00:14:47.89" />
                    <SPLIT distance="1075" swimtime="00:15:10.01" />
                    <SPLIT distance="1100" swimtime="00:15:31.97" />
                    <SPLIT distance="1125" swimtime="00:15:53.84" />
                    <SPLIT distance="1150" swimtime="00:16:15.91" />
                    <SPLIT distance="1175" swimtime="00:16:37.99" />
                    <SPLIT distance="1200" swimtime="00:16:59.93" />
                    <SPLIT distance="1225" swimtime="00:17:21.94" />
                    <SPLIT distance="1250" swimtime="00:17:43.93" />
                    <SPLIT distance="1275" swimtime="00:18:05.80" />
                    <SPLIT distance="1300" swimtime="00:18:27.57" />
                    <SPLIT distance="1325" swimtime="00:18:49.73" />
                    <SPLIT distance="1350" swimtime="00:19:11.76" />
                    <SPLIT distance="1375" swimtime="00:19:33.50" />
                    <SPLIT distance="1400" swimtime="00:19:55.74" />
                    <SPLIT distance="1425" swimtime="00:20:18.17" />
                    <SPLIT distance="1450" swimtime="00:20:40.38" />
                    <SPLIT distance="1475" swimtime="00:21:02.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="325" reactiontime="+74" swimtime="00:02:55.16" resultid="108409" heatid="110669" lane="7" entrytime="00:02:57.93">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.30" />
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="75" swimtime="00:01:00.26" />
                    <SPLIT distance="100" swimtime="00:01:22.71" />
                    <SPLIT distance="125" swimtime="00:01:45.33" />
                    <SPLIT distance="150" swimtime="00:02:08.46" />
                    <SPLIT distance="175" swimtime="00:02:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="108410" heatid="110711" lane="4" entrytime="00:03:07.56" />
                <RESULT eventid="99091" points="331" reactiontime="+82" swimtime="00:01:20.36" resultid="108411" heatid="110732" lane="1" entrytime="00:01:20.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.44" />
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="75" swimtime="00:00:59.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="108412" heatid="110790" lane="5" entrytime="00:06:03.57" />
                <RESULT eventid="99393" points="280" reactiontime="+76" swimtime="00:02:41.44" resultid="108413" heatid="110814" lane="4" entrytime="00:02:38.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.17" />
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="75" swimtime="00:00:58.64" />
                    <SPLIT distance="100" swimtime="00:01:18.99" />
                    <SPLIT distance="125" swimtime="00:01:39.67" />
                    <SPLIT distance="150" swimtime="00:02:00.72" />
                    <SPLIT distance="175" swimtime="00:02:21.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="108414" heatid="110846" lane="8" entrytime="00:05:16.93" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="108397">
              <RESULTS>
                <RESULT eventid="98798" points="443" swimtime="00:00:26.57" resultid="108398" heatid="110610" lane="9" entrytime="00:00:26.47">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="400" reactiontime="+85" swimtime="00:02:28.75" resultid="108399" heatid="110627" lane="6" entrytime="00:02:29.96">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.53" />
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="75" swimtime="00:00:50.53" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="125" swimtime="00:01:31.45" />
                    <SPLIT distance="150" swimtime="00:01:54.16" />
                    <SPLIT distance="175" swimtime="00:02:12.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="414" reactiontime="+78" swimtime="00:00:29.80" resultid="108400" heatid="110660" lane="0" entrytime="00:00:29.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="448" swimtime="00:00:58.73" resultid="108401" heatid="110688" lane="0" entrytime="00:00:58.82">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="75" swimtime="00:00:43.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="394" reactiontime="+84" swimtime="00:00:29.72" resultid="108402" heatid="110742" lane="4" entrytime="00:00:45.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="416" reactiontime="+81" swimtime="00:01:05.51" resultid="108403" heatid="110763" lane="7" entrytime="00:01:04.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.44" />
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="75" swimtime="00:00:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="373" reactiontime="+75" swimtime="00:02:26.65" resultid="108404" heatid="110816" lane="9" entrytime="00:02:25.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.96" />
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="75" swimtime="00:00:51.39" />
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                    <SPLIT distance="125" swimtime="00:01:28.65" />
                    <SPLIT distance="150" swimtime="00:01:47.81" />
                    <SPLIT distance="175" swimtime="00:02:07.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="108405" heatid="110830" lane="5" entrytime="00:00:36.27" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="108439">
              <RESULTS>
                <RESULT eventid="98798" points="293" reactiontime="+82" swimtime="00:00:30.48" resultid="108440" heatid="110603" lane="0" entrytime="00:00:30.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="256" reactiontime="+94" swimtime="00:02:52.47" resultid="108441" heatid="110623" lane="2" entrytime="00:02:54.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.02" />
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="75" swimtime="00:00:59.14" />
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                    <SPLIT distance="125" swimtime="00:01:46.41" />
                    <SPLIT distance="150" swimtime="00:02:13.28" />
                    <SPLIT distance="175" swimtime="00:02:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="228" reactiontime="+76" swimtime="00:00:36.34" resultid="108442" heatid="110656" lane="9" entrytime="00:00:35.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="304" reactiontime="+91" swimtime="00:01:06.82" resultid="108443" heatid="110682" lane="5" entrytime="00:01:08.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.95" />
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="75" swimtime="00:00:49.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="233" reactiontime="+79" swimtime="00:01:19.46" resultid="108444" heatid="110760" lane="3" entrytime="00:01:19.72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.48" />
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                    <SPLIT distance="75" swimtime="00:00:58.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="244" reactiontime="+82" swimtime="00:06:16.87" resultid="108445" heatid="110790" lane="2" entrytime="00:06:14.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.39" />
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="75" swimtime="00:01:01.90" />
                    <SPLIT distance="100" swimtime="00:01:26.85" />
                    <SPLIT distance="125" swimtime="00:01:50.18" />
                    <SPLIT distance="150" swimtime="00:02:12.63" />
                    <SPLIT distance="175" swimtime="00:02:35.47" />
                    <SPLIT distance="200" swimtime="00:02:58.44" />
                    <SPLIT distance="225" swimtime="00:03:27.16" />
                    <SPLIT distance="250" swimtime="00:03:55.55" />
                    <SPLIT distance="275" swimtime="00:04:23.36" />
                    <SPLIT distance="300" swimtime="00:04:51.21" />
                    <SPLIT distance="325" swimtime="00:05:12.81" />
                    <SPLIT distance="350" swimtime="00:05:34.39" />
                    <SPLIT distance="375" swimtime="00:05:56.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="222" reactiontime="+96" swimtime="00:02:54.28" resultid="108446" heatid="110813" lane="6" entrytime="00:02:55.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.97" />
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="75" swimtime="00:01:02.81" />
                    <SPLIT distance="100" swimtime="00:01:25.05" />
                    <SPLIT distance="125" swimtime="00:01:47.60" />
                    <SPLIT distance="150" swimtime="00:02:10.32" />
                    <SPLIT distance="175" swimtime="00:02:33.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="108447" heatid="110848" lane="7" entrytime="00:05:50.91" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-15" firstname="Michał" gender="M" lastname="Skrok" nation="POL" athleteid="108415">
              <RESULTS>
                <RESULT eventid="98798" points="392" reactiontime="+58" swimtime="00:00:27.67" resultid="108416" heatid="110605" lane="4" entrytime="00:00:28.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="430" reactiontime="+69" swimtime="00:02:25.18" resultid="108417" heatid="110626" lane="6" entrytime="00:02:32.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.76" />
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="75" swimtime="00:00:51.93" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="125" swimtime="00:01:30.89" />
                    <SPLIT distance="150" swimtime="00:01:50.73" />
                    <SPLIT distance="175" swimtime="00:02:08.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="433" swimtime="00:02:39.24" resultid="108418" heatid="110670" lane="9" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.41" />
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="75" swimtime="00:00:56.08" />
                    <SPLIT distance="100" swimtime="00:01:16.87" />
                    <SPLIT distance="125" swimtime="00:01:37.66" />
                    <SPLIT distance="150" swimtime="00:01:58.22" />
                    <SPLIT distance="175" swimtime="00:02:18.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="434" reactiontime="+69" swimtime="00:01:06.88" resultid="108419" heatid="110703" lane="6" entrytime="00:01:09.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="75" swimtime="00:00:50.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="464" swimtime="00:01:11.81" resultid="108420" heatid="110733" lane="6" entrytime="00:01:14.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.60" />
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="75" swimtime="00:00:52.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="475" swimtime="00:00:32.35" resultid="108421" heatid="110833" lane="0" entrytime="00:00:34.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="424" reactiontime="+91" swimtime="00:02:00.47" resultid="108448" heatid="110719" lane="0" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.11" />
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="75" swimtime="00:00:44.94" />
                    <SPLIT distance="100" swimtime="00:01:02.00" />
                    <SPLIT distance="125" swimtime="00:01:15.38" />
                    <SPLIT distance="150" swimtime="00:01:32.19" />
                    <SPLIT distance="175" swimtime="00:01:45.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108397" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="108415" number="2" />
                    <RELAYPOSITION athleteid="108422" number="3" />
                    <RELAYPOSITION athleteid="108406" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="ZAC" clubid="108346" name="Mswim Szczecin">
          <CONTACT city="Szczecin" email="jadwiga.w@wp.pl" name="WEBER JADWIGA" phone="601855955" state="ZACH" street="Boguchwały 1 B m 6" zip="71-531" />
          <ATHLETES>
            <ATHLETE birthdate="1960-01-12" firstname="Zbigniew" gender="M" lastname="Szozda" nation="POL" license="G" athleteid="108351">
              <RESULTS>
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="108352" heatid="110667" lane="3" entrytime="00:03:18.00" entrycourse="SCM" />
                <RESULT eventid="98988" points="256" reactiontime="+84" swimtime="00:01:19.70" resultid="108353" heatid="110699" lane="6" entrytime="00:01:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.87" />
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="75" swimtime="00:00:59.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="249" swimtime="00:01:28.34" resultid="108354" heatid="110730" lane="6" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.91" />
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                    <SPLIT distance="75" swimtime="00:01:04.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="203" reactiontime="+84" swimtime="00:01:23.12" resultid="108355" heatid="110760" lane="2" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.30" />
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="75" swimtime="00:01:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="108356" heatid="110812" lane="3" entrytime="00:03:10.00" entrycourse="SCM" />
                <RESULT eventid="99425" points="257" reactiontime="+107" swimtime="00:00:39.67" resultid="108357" heatid="110828" lane="5" entrytime="00:00:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" license="G" athleteid="108347">
              <RESULTS>
                <RESULT eventid="106294" points="232" reactiontime="+90" swimtime="00:00:41.74" resultid="108348" heatid="110648" lane="8" entrytime="00:00:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="242" reactiontime="+90" swimtime="00:01:28.21" resultid="108349" heatid="110755" lane="0" entrytime="00:01:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.75" />
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                    <SPLIT distance="75" swimtime="00:01:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="247" reactiontime="+102" swimtime="00:03:09.95" resultid="108350" heatid="110808" lane="1" entrytime="00:03:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.79" />
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                    <SPLIT distance="75" swimtime="00:01:08.74" />
                    <SPLIT distance="100" swimtime="00:01:32.91" />
                    <SPLIT distance="125" swimtime="00:01:57.05" />
                    <SPLIT distance="150" swimtime="00:02:21.32" />
                    <SPLIT distance="175" swimtime="00:02:46.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NABAIJI" nation="POL" clubid="107102" name="Nabaiji Team Decathlon">
          <CONTACT city="Toruń" email="filip.wojciechowski@decathlon.com" internet="http://www.decathlon.pl" name="Filip Wojciechowski" phone="503414875" street="Decathlon Toruń Copernicus" street2="ul. Żółkiewskiego 15" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1994-01-06" firstname="Paweł" gender="M" lastname="Bednarczyk" nation="POL" athleteid="107110">
              <RESULTS>
                <RESULT eventid="98798" points="629" reactiontime="+68" swimtime="00:00:23.64" resultid="107111" heatid="110613" lane="7" entrytime="00:00:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="662" reactiontime="+75" swimtime="00:00:51.56" resultid="107112" heatid="110689" lane="3" entrytime="00:00:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:25.13" />
                    <SPLIT distance="75" swimtime="00:00:38.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="633" reactiontime="+82" swimtime="00:00:58.98" resultid="107113" heatid="110706" lane="2" entrytime="00:01:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="75" swimtime="00:00:45.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="684" reactiontime="+72" swimtime="00:00:24.74" resultid="107114" heatid="110751" lane="3" entrytime="00:00:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="650" swimtime="00:00:55.91" resultid="107115" heatid="110805" lane="6" entrytime="00:00:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.01" />
                    <SPLIT distance="50" swimtime="00:00:26.37" />
                    <SPLIT distance="75" swimtime="00:00:41.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-04-06" firstname="Martyna" gender="F" lastname="Górajewska" nation="POL" athleteid="107121">
              <RESULTS>
                <RESULT eventid="98777" points="400" swimtime="00:00:31.52" resultid="107122" heatid="110592" lane="9" entrytime="00:00:30.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="341" reactiontime="+78" swimtime="00:01:21.07" resultid="107123" heatid="110694" lane="5" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.21" />
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="75" swimtime="00:01:01.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="359" reactiontime="+76" swimtime="00:00:40.50" resultid="107124" heatid="110822" lane="7" entrytime="00:00:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-04" firstname="Filip" gender="M" lastname="Wojciechowski" nation="POL" athleteid="107103">
              <RESULTS>
                <RESULT eventid="98798" points="520" reactiontime="+71" swimtime="00:00:25.18" resultid="107104" heatid="110612" lane="7" entrytime="00:00:24.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="560" reactiontime="+78" swimtime="00:00:54.52" resultid="107105" heatid="110689" lane="2" entrytime="00:00:54.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.17" />
                    <SPLIT distance="50" swimtime="00:00:25.58" />
                    <SPLIT distance="75" swimtime="00:00:39.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="447" swimtime="00:01:06.22" resultid="107106" heatid="110705" lane="2" entrytime="00:01:05.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.12" />
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="75" swimtime="00:00:51.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="513" reactiontime="+81" swimtime="00:00:27.23" resultid="107107" heatid="110750" lane="2" entrytime="00:00:27.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="531" reactiontime="+71" swimtime="00:02:02.69" resultid="107108" heatid="110778" lane="8" entrytime="00:02:00.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.69" />
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                    <SPLIT distance="75" swimtime="00:00:42.39" />
                    <SPLIT distance="100" swimtime="00:00:58.08" />
                    <SPLIT distance="125" swimtime="00:01:14.11" />
                    <SPLIT distance="150" swimtime="00:01:30.72" />
                    <SPLIT distance="175" swimtime="00:01:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="494" reactiontime="+61" swimtime="00:04:28.39" resultid="107109" heatid="110843" lane="5" entrytime="00:04:18.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                    <SPLIT distance="75" swimtime="00:00:44.16" />
                    <SPLIT distance="100" swimtime="00:01:00.51" />
                    <SPLIT distance="125" swimtime="00:01:17.33" />
                    <SPLIT distance="150" swimtime="00:01:34.45" />
                    <SPLIT distance="175" swimtime="00:01:51.76" />
                    <SPLIT distance="200" swimtime="00:02:09.07" />
                    <SPLIT distance="225" swimtime="00:02:26.46" />
                    <SPLIT distance="250" swimtime="00:02:44.13" />
                    <SPLIT distance="275" swimtime="00:03:01.78" />
                    <SPLIT distance="300" swimtime="00:03:19.87" />
                    <SPLIT distance="325" swimtime="00:03:37.41" />
                    <SPLIT distance="350" swimtime="00:03:54.86" />
                    <SPLIT distance="375" swimtime="00:04:12.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-20" firstname="Rafał" gender="M" lastname="Liszewski" nation="POL" athleteid="107116">
              <RESULTS>
                <RESULT eventid="98798" points="470" reactiontime="+83" swimtime="00:00:26.05" resultid="107117" heatid="110609" lane="2" entrytime="00:00:26.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="383" reactiontime="+76" swimtime="00:00:30.58" resultid="107118" heatid="110658" lane="5" entrytime="00:00:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="431" reactiontime="+79" swimtime="00:01:07.06" resultid="107119" heatid="110703" lane="7" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.78" />
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="75" swimtime="00:00:50.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="517" reactiontime="+72" swimtime="00:00:31.45" resultid="107120" heatid="110833" lane="4" entrytime="00:00:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" region="WA" clubid="106442" name="NENDRE KLAIPEDA">
          <CONTACT state="MAZ" />
          <ATHLETES>
            <ATHLETE birthdate="1962-08-02" firstname=" AIDA" gender="F" nameprefix="VILIMIENE " nation="LTU" athleteid="108922">
              <RESULTS>
                <RESULT eventid="106254" points="353" reactiontime="+96" swimtime="00:21:40.98" resultid="108923" heatid="110640" lane="3" entrytime="00:21:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.39" />
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="75" swimtime="00:00:56.36" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="125" swimtime="00:01:37.37" />
                    <SPLIT distance="150" swimtime="00:01:58.55" />
                    <SPLIT distance="175" swimtime="00:02:19.91" />
                    <SPLIT distance="200" swimtime="00:02:41.40" />
                    <SPLIT distance="225" swimtime="00:03:03.12" />
                    <SPLIT distance="250" swimtime="00:03:24.88" />
                    <SPLIT distance="275" swimtime="00:03:46.55" />
                    <SPLIT distance="300" swimtime="00:04:08.27" />
                    <SPLIT distance="325" swimtime="00:04:30.16" />
                    <SPLIT distance="350" swimtime="00:04:52.13" />
                    <SPLIT distance="375" swimtime="00:05:13.90" />
                    <SPLIT distance="400" swimtime="00:05:35.63" />
                    <SPLIT distance="425" swimtime="00:05:57.46" />
                    <SPLIT distance="450" swimtime="00:06:19.43" />
                    <SPLIT distance="475" swimtime="00:06:41.26" />
                    <SPLIT distance="500" swimtime="00:07:03.07" />
                    <SPLIT distance="525" swimtime="00:07:24.91" />
                    <SPLIT distance="550" swimtime="00:07:47.01" />
                    <SPLIT distance="575" swimtime="00:08:09.21" />
                    <SPLIT distance="600" swimtime="00:08:31.33" />
                    <SPLIT distance="625" swimtime="00:08:53.19" />
                    <SPLIT distance="650" swimtime="00:09:15.31" />
                    <SPLIT distance="675" swimtime="00:09:37.40" />
                    <SPLIT distance="700" swimtime="00:09:59.48" />
                    <SPLIT distance="725" swimtime="00:10:21.46" />
                    <SPLIT distance="750" swimtime="00:10:43.52" />
                    <SPLIT distance="775" swimtime="00:11:05.39" />
                    <SPLIT distance="800" swimtime="00:11:27.30" />
                    <SPLIT distance="825" swimtime="00:11:49.35" />
                    <SPLIT distance="850" swimtime="00:12:11.16" />
                    <SPLIT distance="875" swimtime="00:12:33.13" />
                    <SPLIT distance="900" swimtime="00:12:55.09" />
                    <SPLIT distance="925" swimtime="00:13:17.03" />
                    <SPLIT distance="950" swimtime="00:13:38.92" />
                    <SPLIT distance="975" swimtime="00:14:01.02" />
                    <SPLIT distance="1000" swimtime="00:14:23.12" />
                    <SPLIT distance="1025" swimtime="00:14:45.17" />
                    <SPLIT distance="1050" swimtime="00:15:07.22" />
                    <SPLIT distance="1075" swimtime="00:15:29.28" />
                    <SPLIT distance="1100" swimtime="00:15:51.11" />
                    <SPLIT distance="1125" swimtime="00:16:13.05" />
                    <SPLIT distance="1150" swimtime="00:16:35.07" />
                    <SPLIT distance="1175" swimtime="00:16:57.56" />
                    <SPLIT distance="1200" swimtime="00:17:19.53" />
                    <SPLIT distance="1225" swimtime="00:17:41.59" />
                    <SPLIT distance="1250" swimtime="00:18:03.47" />
                    <SPLIT distance="1275" swimtime="00:18:25.43" />
                    <SPLIT distance="1300" swimtime="00:18:47.37" />
                    <SPLIT distance="1325" swimtime="00:19:09.22" />
                    <SPLIT distance="1350" swimtime="00:19:31.02" />
                    <SPLIT distance="1375" swimtime="00:19:52.88" />
                    <SPLIT distance="1400" swimtime="00:20:14.94" />
                    <SPLIT distance="1425" swimtime="00:20:36.79" />
                    <SPLIT distance="1450" swimtime="00:20:58.72" />
                    <SPLIT distance="1475" swimtime="00:21:20.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="344" reactiontime="+82" swimtime="00:01:12.64" resultid="108924" heatid="110675" lane="8" entrytime="00:01:12.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.38" />
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="75" swimtime="00:00:54.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="310" swimtime="00:06:23.28" resultid="108925" heatid="110787" lane="0" entrytime="00:06:31.28">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.44" />
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="75" swimtime="00:01:05.18" />
                    <SPLIT distance="100" swimtime="00:01:29.97" />
                    <SPLIT distance="125" swimtime="00:01:56.15" />
                    <SPLIT distance="150" swimtime="00:02:21.30" />
                    <SPLIT distance="175" swimtime="00:02:45.97" />
                    <SPLIT distance="200" swimtime="00:03:10.81" />
                    <SPLIT distance="225" swimtime="00:03:37.47" />
                    <SPLIT distance="250" swimtime="00:04:04.45" />
                    <SPLIT distance="275" swimtime="00:04:31.21" />
                    <SPLIT distance="300" swimtime="00:04:58.32" />
                    <SPLIT distance="325" swimtime="00:05:20.75" />
                    <SPLIT distance="350" swimtime="00:05:41.98" />
                    <SPLIT distance="375" swimtime="00:06:03.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="370" swimtime="00:05:26.49" resultid="108926" heatid="110839" lane="0" entrytime="00:05:29.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.19" />
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="75" swimtime="00:00:56.26" />
                    <SPLIT distance="100" swimtime="00:01:16.65" />
                    <SPLIT distance="125" swimtime="00:01:37.19" />
                    <SPLIT distance="150" swimtime="00:01:57.92" />
                    <SPLIT distance="175" swimtime="00:02:18.74" />
                    <SPLIT distance="200" swimtime="00:02:39.86" />
                    <SPLIT distance="225" swimtime="00:03:00.57" />
                    <SPLIT distance="250" swimtime="00:03:22.02" />
                    <SPLIT distance="275" swimtime="00:03:42.62" />
                    <SPLIT distance="300" swimtime="00:04:03.53" />
                    <SPLIT distance="325" swimtime="00:04:24.42" />
                    <SPLIT distance="350" swimtime="00:04:45.54" />
                    <SPLIT distance="375" swimtime="00:05:05.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" status="DNS" swimtime="00:00:00.00" resultid="106494" heatid="110718" lane="7" entrytime="00:02:08.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" status="DNS" swimtime="00:00:00.00" resultid="106495" heatid="110783" lane="2" entrytime="00:01:56.00" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" status="DNS" swimtime="00:00:00.00" resultid="106492" heatid="110631" lane="0" entrytime="00:02:08.00" />
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="106493" heatid="110837" lane="3" entrytime="00:02:15.00" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="107740" name="One Man Team">
          <CONTACT city="Daszewice" email="gmo@o2.pl" internet="open-water.pl" name="Grzegorz Monczak" phone="608639696" state="WLKP" street="ul. Przy Lesie 17" zip="61-160" />
          <ATHLETES>
            <ATHLETE birthdate="1973-05-25" firstname="Grzegorz" gender="M" lastname="Monczak" nation="POL" athleteid="107741">
              <RESULTS>
                <RESULT eventid="98830" points="352" reactiontime="+70" swimtime="00:02:35.22" resultid="107742" heatid="110625" lane="6" entrytime="00:02:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.21" />
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                    <SPLIT distance="75" swimtime="00:00:55.20" />
                    <SPLIT distance="100" swimtime="00:01:15.05" />
                    <SPLIT distance="125" swimtime="00:01:37.89" />
                    <SPLIT distance="150" swimtime="00:02:01.29" />
                    <SPLIT distance="175" swimtime="00:02:19.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="423" reactiontime="+97" swimtime="00:18:49.51" resultid="107743" heatid="110641" lane="3" entrytime="00:18:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.26" />
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="75" swimtime="00:00:52.25" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="125" swimtime="00:01:29.07" />
                    <SPLIT distance="150" swimtime="00:01:47.73" />
                    <SPLIT distance="175" swimtime="00:02:06.19" />
                    <SPLIT distance="200" swimtime="00:02:24.81" />
                    <SPLIT distance="225" swimtime="00:02:43.49" />
                    <SPLIT distance="250" swimtime="00:03:02.20" />
                    <SPLIT distance="275" swimtime="00:03:20.94" />
                    <SPLIT distance="300" swimtime="00:03:39.57" />
                    <SPLIT distance="325" swimtime="00:03:58.15" />
                    <SPLIT distance="350" swimtime="00:04:16.91" />
                    <SPLIT distance="375" swimtime="00:04:35.49" />
                    <SPLIT distance="400" swimtime="00:04:55.06" />
                    <SPLIT distance="425" swimtime="00:05:13.95" />
                    <SPLIT distance="450" swimtime="00:05:32.73" />
                    <SPLIT distance="475" swimtime="00:05:51.48" />
                    <SPLIT distance="500" swimtime="00:06:10.29" />
                    <SPLIT distance="525" swimtime="00:06:29.68" />
                    <SPLIT distance="550" swimtime="00:06:48.82" />
                    <SPLIT distance="575" swimtime="00:07:07.82" />
                    <SPLIT distance="600" swimtime="00:07:26.67" />
                    <SPLIT distance="625" swimtime="00:07:45.50" />
                    <SPLIT distance="650" swimtime="00:08:04.20" />
                    <SPLIT distance="675" swimtime="00:08:23.03" />
                    <SPLIT distance="700" swimtime="00:08:41.86" />
                    <SPLIT distance="725" swimtime="00:09:00.77" />
                    <SPLIT distance="750" swimtime="00:09:19.50" />
                    <SPLIT distance="775" swimtime="00:09:38.34" />
                    <SPLIT distance="800" swimtime="00:09:57.23" />
                    <SPLIT distance="825" swimtime="00:10:16.03" />
                    <SPLIT distance="850" swimtime="00:10:35.03" />
                    <SPLIT distance="875" swimtime="00:10:53.91" />
                    <SPLIT distance="900" swimtime="00:11:12.94" />
                    <SPLIT distance="925" swimtime="00:11:32.08" />
                    <SPLIT distance="950" swimtime="00:11:51.14" />
                    <SPLIT distance="975" swimtime="00:12:10.16" />
                    <SPLIT distance="1000" swimtime="00:12:29.07" />
                    <SPLIT distance="1025" swimtime="00:12:48.33" />
                    <SPLIT distance="1050" swimtime="00:13:07.31" />
                    <SPLIT distance="1075" swimtime="00:13:26.32" />
                    <SPLIT distance="1100" swimtime="00:13:45.20" />
                    <SPLIT distance="1125" swimtime="00:14:04.58" />
                    <SPLIT distance="1150" swimtime="00:14:24.24" />
                    <SPLIT distance="1175" swimtime="00:14:43.21" />
                    <SPLIT distance="1200" swimtime="00:15:02.55" />
                    <SPLIT distance="1225" swimtime="00:15:21.41" />
                    <SPLIT distance="1250" swimtime="00:15:40.42" />
                    <SPLIT distance="1275" swimtime="00:15:59.45" />
                    <SPLIT distance="1300" swimtime="00:16:18.48" />
                    <SPLIT distance="1325" swimtime="00:16:37.54" />
                    <SPLIT distance="1350" swimtime="00:16:56.24" />
                    <SPLIT distance="1375" swimtime="00:17:15.44" />
                    <SPLIT distance="1400" swimtime="00:17:34.53" />
                    <SPLIT distance="1425" swimtime="00:17:53.39" />
                    <SPLIT distance="1450" swimtime="00:18:12.37" />
                    <SPLIT distance="1475" swimtime="00:18:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="408" reactiontime="+87" swimtime="00:01:00.59" resultid="107744" heatid="110687" lane="1" entrytime="00:00:59.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.23" />
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="75" swimtime="00:00:45.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="322" reactiontime="+56" swimtime="00:01:13.86" resultid="107745" heatid="110702" lane="6" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.38" />
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="75" swimtime="00:00:56.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="268" reactiontime="+84" swimtime="00:01:26.21" resultid="107746" heatid="110730" lane="4" entrytime="00:01:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.13" />
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="75" swimtime="00:01:03.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="435" reactiontime="+98" swimtime="00:02:11.08" resultid="107747" heatid="110777" lane="1" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.59" />
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="75" swimtime="00:00:48.78" />
                    <SPLIT distance="100" swimtime="00:01:05.38" />
                    <SPLIT distance="125" swimtime="00:01:21.91" />
                    <SPLIT distance="150" swimtime="00:01:38.53" />
                    <SPLIT distance="175" swimtime="00:01:54.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="250" reactiontime="+84" swimtime="00:01:16.88" resultid="107748" heatid="110801" lane="4" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.61" />
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="75" swimtime="00:00:56.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="438" reactiontime="+101" swimtime="00:04:39.42" resultid="107749" heatid="110843" lane="1" entrytime="00:04:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.87" />
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="75" swimtime="00:00:50.23" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="125" swimtime="00:01:25.25" />
                    <SPLIT distance="150" swimtime="00:01:42.82" />
                    <SPLIT distance="175" swimtime="00:02:00.50" />
                    <SPLIT distance="200" swimtime="00:02:18.49" />
                    <SPLIT distance="225" swimtime="00:02:36.46" />
                    <SPLIT distance="250" swimtime="00:02:54.12" />
                    <SPLIT distance="275" swimtime="00:03:11.85" />
                    <SPLIT distance="300" swimtime="00:03:29.56" />
                    <SPLIT distance="325" swimtime="00:03:47.24" />
                    <SPLIT distance="350" swimtime="00:04:04.76" />
                    <SPLIT distance="375" swimtime="00:04:22.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORSOPOLE" nation="POL" region="OPO" clubid="108887" name="ORS Opole">
          <CONTACT name="Kania" />
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="108903">
              <RESULTS>
                <RESULT eventid="98814" points="388" reactiontime="+76" swimtime="00:02:46.96" resultid="108904" heatid="110617" lane="4" entrytime="00:02:46.39">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.93" />
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="75" swimtime="00:00:58.03" />
                    <SPLIT distance="100" swimtime="00:01:20.57" />
                    <SPLIT distance="125" swimtime="00:01:44.51" />
                    <SPLIT distance="150" swimtime="00:02:09.05" />
                    <SPLIT distance="175" swimtime="00:02:29.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="359" reactiontime="+95" swimtime="00:11:14.40" resultid="108905" heatid="110633" lane="5" entrytime="00:11:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.70" />
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="75" swimtime="00:00:58.09" />
                    <SPLIT distance="100" swimtime="00:01:18.97" />
                    <SPLIT distance="125" swimtime="00:01:39.73" />
                    <SPLIT distance="150" swimtime="00:02:01.07" />
                    <SPLIT distance="175" swimtime="00:02:22.41" />
                    <SPLIT distance="200" swimtime="00:02:43.68" />
                    <SPLIT distance="225" swimtime="00:03:04.99" />
                    <SPLIT distance="250" swimtime="00:03:26.59" />
                    <SPLIT distance="275" swimtime="00:03:48.00" />
                    <SPLIT distance="300" swimtime="00:04:09.43" />
                    <SPLIT distance="325" swimtime="00:04:31.28" />
                    <SPLIT distance="350" swimtime="00:04:52.73" />
                    <SPLIT distance="375" swimtime="00:05:14.50" />
                    <SPLIT distance="400" swimtime="00:05:35.83" />
                    <SPLIT distance="425" swimtime="00:05:57.58" />
                    <SPLIT distance="450" swimtime="00:06:18.89" />
                    <SPLIT distance="475" swimtime="00:06:40.74" />
                    <SPLIT distance="500" swimtime="00:07:02.09" />
                    <SPLIT distance="525" swimtime="00:07:24.18" />
                    <SPLIT distance="550" swimtime="00:07:45.90" />
                    <SPLIT distance="575" swimtime="00:08:07.56" />
                    <SPLIT distance="600" swimtime="00:08:29.12" />
                    <SPLIT distance="625" swimtime="00:08:50.72" />
                    <SPLIT distance="650" swimtime="00:09:11.93" />
                    <SPLIT distance="675" swimtime="00:09:33.72" />
                    <SPLIT distance="700" swimtime="00:09:55.02" />
                    <SPLIT distance="725" swimtime="00:10:16.63" />
                    <SPLIT distance="750" swimtime="00:10:37.10" />
                    <SPLIT distance="775" swimtime="00:10:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="401" swimtime="00:05:51.57" resultid="108906" heatid="110787" lane="6" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.59" />
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="75" swimtime="00:01:02.61" />
                    <SPLIT distance="100" swimtime="00:01:26.51" />
                    <SPLIT distance="125" swimtime="00:01:49.35" />
                    <SPLIT distance="150" swimtime="00:02:11.28" />
                    <SPLIT distance="175" swimtime="00:02:33.32" />
                    <SPLIT distance="200" swimtime="00:02:56.01" />
                    <SPLIT distance="225" swimtime="00:03:20.50" />
                    <SPLIT distance="250" swimtime="00:03:45.57" />
                    <SPLIT distance="275" swimtime="00:04:10.29" />
                    <SPLIT distance="300" swimtime="00:04:35.10" />
                    <SPLIT distance="325" swimtime="00:04:55.99" />
                    <SPLIT distance="350" swimtime="00:05:15.16" />
                    <SPLIT distance="375" swimtime="00:05:34.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="374" swimtime="00:01:15.77" resultid="108907" heatid="110796" lane="9" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.67" />
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="75" swimtime="00:00:55.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="386" reactiontime="+90" swimtime="00:05:22.02" resultid="108908" heatid="110839" lane="8" entrytime="00:05:20.07">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.87" />
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                    <SPLIT distance="75" swimtime="00:00:55.62" />
                    <SPLIT distance="100" swimtime="00:01:16.09" />
                    <SPLIT distance="125" swimtime="00:01:36.70" />
                    <SPLIT distance="150" swimtime="00:01:57.35" />
                    <SPLIT distance="175" swimtime="00:02:18.23" />
                    <SPLIT distance="200" swimtime="00:02:39.04" />
                    <SPLIT distance="225" swimtime="00:02:59.86" />
                    <SPLIT distance="250" swimtime="00:03:20.87" />
                    <SPLIT distance="275" swimtime="00:03:42.01" />
                    <SPLIT distance="300" swimtime="00:04:03.17" />
                    <SPLIT distance="325" swimtime="00:04:24.00" />
                    <SPLIT distance="350" swimtime="00:04:44.38" />
                    <SPLIT distance="375" swimtime="00:05:04.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" clubid="110209" name="OSIR Inowrocław">
          <ATHLETES>
            <ATHLETE birthdate="1937-09-19" firstname="ZYGMUNT" gender="M" lastname="LEWANDOWSKI" nation="POL" athleteid="106347">
              <RESULTS>
                <RESULT eventid="98891" points="98" reactiontime="+100" swimtime="00:16:00.36" resultid="106348" heatid="110638" lane="2" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.44" />
                    <SPLIT distance="50" swimtime="00:00:51.03" />
                    <SPLIT distance="75" swimtime="00:01:18.67" />
                    <SPLIT distance="100" swimtime="00:01:47.01" />
                    <SPLIT distance="125" swimtime="00:02:15.80" />
                    <SPLIT distance="150" swimtime="00:02:45.60" />
                    <SPLIT distance="175" swimtime="00:03:14.81" />
                    <SPLIT distance="200" swimtime="00:03:44.20" />
                    <SPLIT distance="225" swimtime="00:04:13.50" />
                    <SPLIT distance="250" swimtime="00:04:43.33" />
                    <SPLIT distance="275" swimtime="00:05:12.80" />
                    <SPLIT distance="300" swimtime="00:05:42.71" />
                    <SPLIT distance="325" swimtime="00:06:12.43" />
                    <SPLIT distance="350" swimtime="00:06:42.90" />
                    <SPLIT distance="375" swimtime="00:07:13.08" />
                    <SPLIT distance="400" swimtime="00:07:44.24" />
                    <SPLIT distance="425" swimtime="00:08:15.02" />
                    <SPLIT distance="450" swimtime="00:08:46.52" />
                    <SPLIT distance="475" swimtime="00:09:17.02" />
                    <SPLIT distance="500" swimtime="00:09:48.55" />
                    <SPLIT distance="525" swimtime="00:10:19.08" />
                    <SPLIT distance="550" swimtime="00:10:50.83" />
                    <SPLIT distance="575" swimtime="00:11:21.44" />
                    <SPLIT distance="600" swimtime="00:11:52.92" />
                    <SPLIT distance="625" swimtime="00:12:23.22" />
                    <SPLIT distance="650" swimtime="00:12:54.14" />
                    <SPLIT distance="675" swimtime="00:13:24.84" />
                    <SPLIT distance="700" swimtime="00:13:55.96" />
                    <SPLIT distance="725" swimtime="00:14:26.61" />
                    <SPLIT distance="750" swimtime="00:14:58.40" />
                    <SPLIT distance="775" swimtime="00:15:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="102" swimtime="00:01:35.99" resultid="106349" heatid="110679" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.04" />
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                    <SPLIT distance="75" swimtime="00:01:10.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="100" reactiontime="+106" swimtime="00:03:33.79" resultid="106350" heatid="110769" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.69" />
                    <SPLIT distance="50" swimtime="00:00:49.58" />
                    <SPLIT distance="75" swimtime="00:01:16.61" />
                    <SPLIT distance="100" swimtime="00:01:44.67" />
                    <SPLIT distance="125" swimtime="00:02:12.02" />
                    <SPLIT distance="150" swimtime="00:02:40.42" />
                    <SPLIT distance="175" swimtime="00:03:08.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="97" reactiontime="+106" swimtime="00:07:40.66" resultid="106351" heatid="110851" lane="1" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.98" />
                    <SPLIT distance="50" swimtime="00:00:52.86" />
                    <SPLIT distance="75" swimtime="00:01:21.07" />
                    <SPLIT distance="100" swimtime="00:01:50.30" />
                    <SPLIT distance="125" swimtime="00:02:19.63" />
                    <SPLIT distance="150" swimtime="00:02:48.73" />
                    <SPLIT distance="175" swimtime="00:03:18.83" />
                    <SPLIT distance="200" swimtime="00:03:48.83" />
                    <SPLIT distance="225" swimtime="00:04:18.49" />
                    <SPLIT distance="250" swimtime="00:04:48.23" />
                    <SPLIT distance="275" swimtime="00:05:17.33" />
                    <SPLIT distance="300" swimtime="00:05:46.81" />
                    <SPLIT distance="325" swimtime="00:06:15.85" />
                    <SPLIT distance="350" swimtime="00:06:45.39" />
                    <SPLIT distance="375" swimtime="00:07:13.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PAKA" nation="POL" region="SLA" clubid="107047" name="Pałac Katowice">
          <CONTACT name="Bucholz" phone="606 135 860" />
          <ATHLETES>
            <ATHLETE birthdate="1972-02-13" firstname="Damian" gender="M" lastname="Hostyński" nation="POL" athleteid="107052" />
            <ATHLETE birthdate="1972-09-12" firstname="Mateusz" gender="M" lastname="Matusiewicz" nation="POL" athleteid="107054" />
            <ATHLETE birthdate="1973-08-30" firstname="Jacek" gender="M" lastname="Kobylczak" nation="POL" athleteid="107053" />
            <ATHLETE birthdate="1972-01-26" firstname="Tomasz" gender="M" lastname="Bucholz" nation="POL" athleteid="107048">
              <RESULTS>
                <RESULT eventid="98891" points="337" reactiontime="+106" swimtime="00:10:37.03" resultid="107049" heatid="110635" lane="2" entrytime="00:09:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.01" />
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="75" swimtime="00:00:52.06" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="125" swimtime="00:01:30.21" />
                    <SPLIT distance="150" swimtime="00:01:49.73" />
                    <SPLIT distance="175" swimtime="00:02:09.32" />
                    <SPLIT distance="200" swimtime="00:02:29.34" />
                    <SPLIT distance="225" swimtime="00:02:48.88" />
                    <SPLIT distance="250" swimtime="00:03:08.43" />
                    <SPLIT distance="275" swimtime="00:03:28.97" />
                    <SPLIT distance="300" swimtime="00:03:49.17" />
                    <SPLIT distance="325" swimtime="00:04:09.80" />
                    <SPLIT distance="350" swimtime="00:04:30.34" />
                    <SPLIT distance="375" swimtime="00:04:50.68" />
                    <SPLIT distance="400" swimtime="00:05:11.43" />
                    <SPLIT distance="425" swimtime="00:05:32.43" />
                    <SPLIT distance="450" swimtime="00:05:52.84" />
                    <SPLIT distance="475" swimtime="00:06:13.55" />
                    <SPLIT distance="500" swimtime="00:06:34.18" />
                    <SPLIT distance="525" swimtime="00:06:54.75" />
                    <SPLIT distance="550" swimtime="00:07:15.35" />
                    <SPLIT distance="575" swimtime="00:07:35.93" />
                    <SPLIT distance="600" swimtime="00:07:56.18" />
                    <SPLIT distance="625" swimtime="00:08:16.63" />
                    <SPLIT distance="650" swimtime="00:08:37.13" />
                    <SPLIT distance="675" swimtime="00:08:57.12" />
                    <SPLIT distance="700" swimtime="00:09:17.66" />
                    <SPLIT distance="725" swimtime="00:09:38.25" />
                    <SPLIT distance="750" swimtime="00:09:58.58" />
                    <SPLIT distance="775" swimtime="00:10:18.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="286" reactiontime="+93" swimtime="00:01:16.85" resultid="107050" heatid="110699" lane="5" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.96" />
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="75" swimtime="00:00:59.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="107051" heatid="110791" lane="1" entrytime="00:05:51.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="250" reactiontime="+95" swimtime="00:02:23.55" resultid="107055" heatid="110717" lane="7" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.16" />
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                    <SPLIT distance="75" swimtime="00:00:55.16" />
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="125" swimtime="00:01:32.78" />
                    <SPLIT distance="150" swimtime="00:01:51.62" />
                    <SPLIT distance="175" swimtime="00:02:07.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107053" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="107052" number="2" reactiontime="+83" />
                    <RELAYPOSITION athleteid="107048" number="3" reactiontime="+91" />
                    <RELAYPOSITION athleteid="107054" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="311" reactiontime="+92" swimtime="00:02:01.85" resultid="107056" heatid="110782" lane="5" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.46" />
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="75" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:03.43" />
                    <SPLIT distance="125" swimtime="00:01:17.56" />
                    <SPLIT distance="150" swimtime="00:01:33.03" />
                    <SPLIT distance="175" swimtime="00:01:46.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107052" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="107054" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="107053" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="107048" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="109163" name="Plavecký klub Stráž pod Ralskem " shortname="PK SpR">
          <ATHLETES>
            <ATHLETE birthdate="1964-01-01" firstname="Jiří" gender="M" lastname="Janovský" nation="CZE" athleteid="109164">
              <RESULTS>
                <RESULT eventid="106256" points="314" swimtime="00:20:47.12" resultid="109165" heatid="110641" lane="9" entrytime="00:21:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.92" />
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="75" swimtime="00:00:55.55" />
                    <SPLIT distance="100" swimtime="00:01:15.85" />
                    <SPLIT distance="125" swimtime="00:01:35.96" />
                    <SPLIT distance="150" swimtime="00:01:56.32" />
                    <SPLIT distance="175" swimtime="00:02:16.01" />
                    <SPLIT distance="200" swimtime="00:02:36.96" />
                    <SPLIT distance="225" swimtime="00:02:56.59" />
                    <SPLIT distance="250" swimtime="00:03:17.41" />
                    <SPLIT distance="275" swimtime="00:03:37.87" />
                    <SPLIT distance="300" swimtime="00:03:58.50" />
                    <SPLIT distance="325" swimtime="00:04:18.92" />
                    <SPLIT distance="350" swimtime="00:05:21.38" />
                    <SPLIT distance="375" swimtime="00:05:00.66" />
                    <SPLIT distance="400" swimtime="00:06:03.42" />
                    <SPLIT distance="425" swimtime="00:05:42.55" />
                    <SPLIT distance="450" swimtime="00:06:45.07" />
                    <SPLIT distance="475" swimtime="00:06:23.75" />
                    <SPLIT distance="525" swimtime="00:07:05.87" />
                    <SPLIT distance="550" swimtime="00:07:27.22" />
                    <SPLIT distance="575" swimtime="00:07:47.98" />
                    <SPLIT distance="600" swimtime="00:08:09.28" />
                    <SPLIT distance="625" swimtime="00:08:30.03" />
                    <SPLIT distance="650" swimtime="00:08:51.12" />
                    <SPLIT distance="675" swimtime="00:09:12.07" />
                    <SPLIT distance="700" swimtime="00:09:33.58" />
                    <SPLIT distance="725" swimtime="00:09:54.74" />
                    <SPLIT distance="750" swimtime="00:10:58.42" />
                    <SPLIT distance="775" swimtime="00:10:36.93" />
                    <SPLIT distance="825" swimtime="00:11:19.19" />
                    <SPLIT distance="875" swimtime="00:12:01.81" />
                    <SPLIT distance="900" swimtime="00:12:22.53" />
                    <SPLIT distance="925" swimtime="00:12:43.49" />
                    <SPLIT distance="975" swimtime="00:13:25.91" />
                    <SPLIT distance="1000" swimtime="00:13:46.87" />
                    <SPLIT distance="1025" swimtime="00:14:07.88" />
                    <SPLIT distance="1050" swimtime="00:14:29.23" />
                    <SPLIT distance="1075" swimtime="00:14:50.36" />
                    <SPLIT distance="1100" swimtime="00:15:11.16" />
                    <SPLIT distance="1125" swimtime="00:15:32.43" />
                    <SPLIT distance="1150" swimtime="00:15:53.90" />
                    <SPLIT distance="1175" swimtime="00:16:15.21" />
                    <SPLIT distance="1200" swimtime="00:16:36.35" />
                    <SPLIT distance="1225" swimtime="00:16:56.81" />
                    <SPLIT distance="1250" swimtime="00:17:18.63" />
                    <SPLIT distance="1275" swimtime="00:17:39.72" />
                    <SPLIT distance="1300" swimtime="00:18:00.90" />
                    <SPLIT distance="1325" swimtime="00:18:21.52" />
                    <SPLIT distance="1350" swimtime="00:18:42.69" />
                    <SPLIT distance="1375" swimtime="00:19:03.52" />
                    <SPLIT distance="1400" swimtime="00:19:24.74" />
                    <SPLIT distance="1425" swimtime="00:19:45.67" />
                    <SPLIT distance="1450" swimtime="00:20:06.38" />
                    <SPLIT distance="1475" swimtime="00:20:26.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="293" reactiontime="+117" swimtime="00:01:07.62" resultid="109166" heatid="110682" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.72" />
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="75" swimtime="00:00:50.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="260" reactiontime="+113" swimtime="00:06:08.86" resultid="109167" heatid="110790" lane="1" entrytime="00:06:18.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.97" />
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="75" swimtime="00:00:59.52" />
                    <SPLIT distance="100" swimtime="00:01:22.28" />
                    <SPLIT distance="125" swimtime="00:01:46.51" />
                    <SPLIT distance="150" swimtime="00:02:09.08" />
                    <SPLIT distance="175" swimtime="00:02:32.00" />
                    <SPLIT distance="200" swimtime="00:02:55.21" />
                    <SPLIT distance="225" swimtime="00:03:22.56" />
                    <SPLIT distance="250" swimtime="00:03:50.26" />
                    <SPLIT distance="275" swimtime="00:04:18.29" />
                    <SPLIT distance="300" swimtime="00:04:47.03" />
                    <SPLIT distance="325" swimtime="00:05:08.18" />
                    <SPLIT distance="350" swimtime="00:05:29.12" />
                    <SPLIT distance="375" swimtime="00:05:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="330" swimtime="00:05:07.05" resultid="109168" heatid="110846" lane="0" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.51" />
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="75" swimtime="00:00:54.29" />
                    <SPLIT distance="100" swimtime="00:01:13.34" />
                    <SPLIT distance="125" swimtime="00:01:32.50" />
                    <SPLIT distance="150" swimtime="00:01:51.92" />
                    <SPLIT distance="175" swimtime="00:02:11.23" />
                    <SPLIT distance="200" swimtime="00:02:30.63" />
                    <SPLIT distance="225" swimtime="00:02:49.90" />
                    <SPLIT distance="250" swimtime="00:03:09.78" />
                    <SPLIT distance="275" swimtime="00:03:29.19" />
                    <SPLIT distance="300" swimtime="00:03:49.14" />
                    <SPLIT distance="325" swimtime="00:04:08.80" />
                    <SPLIT distance="350" swimtime="00:04:28.98" />
                    <SPLIT distance="375" swimtime="00:04:48.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="109136" name="Polish Extreme Ice Swimming">
          <ATHLETES>
            <ATHLETE birthdate="1975-03-01" firstname="PIOTR" gender="M" lastname="BIANKOWSKI " nation="POL" athleteid="109137">
              <RESULTS>
                <RESULT eventid="98798" points="277" reactiontime="+68" swimtime="00:00:31.05" resultid="109138" heatid="110599" lane="7" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="261" reactiontime="+110" swimtime="00:22:06.38" resultid="109139" heatid="110642" lane="3" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.29" />
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="75" swimtime="00:00:59.46" />
                    <SPLIT distance="100" swimtime="00:01:20.51" />
                    <SPLIT distance="125" swimtime="00:01:41.90" />
                    <SPLIT distance="150" swimtime="00:02:03.23" />
                    <SPLIT distance="175" swimtime="00:02:25.08" />
                    <SPLIT distance="200" swimtime="00:02:46.74" />
                    <SPLIT distance="225" swimtime="00:03:08.26" />
                    <SPLIT distance="250" swimtime="00:03:29.85" />
                    <SPLIT distance="275" swimtime="00:03:51.70" />
                    <SPLIT distance="300" swimtime="00:04:13.64" />
                    <SPLIT distance="325" swimtime="00:04:35.76" />
                    <SPLIT distance="350" swimtime="00:04:57.52" />
                    <SPLIT distance="375" swimtime="00:05:19.55" />
                    <SPLIT distance="400" swimtime="00:05:41.63" />
                    <SPLIT distance="425" swimtime="00:06:03.93" />
                    <SPLIT distance="450" swimtime="00:06:26.03" />
                    <SPLIT distance="475" swimtime="00:06:48.25" />
                    <SPLIT distance="500" swimtime="00:07:10.40" />
                    <SPLIT distance="525" swimtime="00:07:32.72" />
                    <SPLIT distance="550" swimtime="00:07:54.87" />
                    <SPLIT distance="575" swimtime="00:08:17.00" />
                    <SPLIT distance="600" swimtime="00:08:39.23" />
                    <SPLIT distance="625" swimtime="00:09:01.67" />
                    <SPLIT distance="650" swimtime="00:09:23.89" />
                    <SPLIT distance="675" swimtime="00:09:46.53" />
                    <SPLIT distance="700" swimtime="00:10:08.72" />
                    <SPLIT distance="725" swimtime="00:10:31.41" />
                    <SPLIT distance="750" swimtime="00:10:53.59" />
                    <SPLIT distance="775" swimtime="00:11:16.22" />
                    <SPLIT distance="800" swimtime="00:11:38.64" />
                    <SPLIT distance="825" swimtime="00:12:00.99" />
                    <SPLIT distance="850" swimtime="00:12:23.36" />
                    <SPLIT distance="875" swimtime="00:12:45.88" />
                    <SPLIT distance="900" swimtime="00:13:08.17" />
                    <SPLIT distance="925" swimtime="00:13:30.53" />
                    <SPLIT distance="950" swimtime="00:13:52.89" />
                    <SPLIT distance="975" swimtime="00:14:15.43" />
                    <SPLIT distance="1000" swimtime="00:14:38.18" />
                    <SPLIT distance="1025" swimtime="00:15:01.08" />
                    <SPLIT distance="1050" swimtime="00:15:23.42" />
                    <SPLIT distance="1075" swimtime="00:15:46.23" />
                    <SPLIT distance="1100" swimtime="00:16:08.59" />
                    <SPLIT distance="1125" swimtime="00:16:31.29" />
                    <SPLIT distance="1150" swimtime="00:16:53.59" />
                    <SPLIT distance="1175" swimtime="00:17:16.74" />
                    <SPLIT distance="1200" swimtime="00:17:39.11" />
                    <SPLIT distance="1225" swimtime="00:18:01.66" />
                    <SPLIT distance="1250" swimtime="00:18:24.20" />
                    <SPLIT distance="1275" swimtime="00:18:46.93" />
                    <SPLIT distance="1300" swimtime="00:19:09.44" />
                    <SPLIT distance="1325" swimtime="00:19:32.26" />
                    <SPLIT distance="1350" swimtime="00:19:55.00" />
                    <SPLIT distance="1375" swimtime="00:20:17.86" />
                    <SPLIT distance="1400" swimtime="00:20:40.36" />
                    <SPLIT distance="1425" swimtime="00:21:02.63" />
                    <SPLIT distance="1450" swimtime="00:21:24.53" />
                    <SPLIT distance="1475" swimtime="00:21:46.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="225" reactiontime="+55" swimtime="00:02:58.44" resultid="109140" heatid="110711" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.33" />
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                    <SPLIT distance="75" swimtime="00:00:59.85" />
                    <SPLIT distance="100" swimtime="00:01:22.44" />
                    <SPLIT distance="125" swimtime="00:01:45.69" />
                    <SPLIT distance="150" swimtime="00:02:09.39" />
                    <SPLIT distance="175" swimtime="00:02:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="263" reactiontime="+90" swimtime="00:00:34.02" resultid="109141" heatid="110743" lane="1" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="283" swimtime="00:02:31.26" resultid="109142" heatid="110772" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.29" />
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="75" swimtime="00:00:54.40" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="125" swimtime="00:01:33.99" />
                    <SPLIT distance="150" swimtime="00:01:54.34" />
                    <SPLIT distance="175" swimtime="00:02:14.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="234" swimtime="00:01:18.59" resultid="109143" heatid="110799" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.01" />
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="75" swimtime="00:00:58.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="265" reactiontime="+54" swimtime="00:05:30.13" resultid="109144" heatid="110850" lane="7" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.65" />
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="75" swimtime="00:00:57.07" />
                    <SPLIT distance="100" swimtime="00:01:18.22" />
                    <SPLIT distance="125" swimtime="00:01:39.67" />
                    <SPLIT distance="150" swimtime="00:02:00.77" />
                    <SPLIT distance="175" swimtime="00:02:22.29" />
                    <SPLIT distance="200" swimtime="00:02:43.61" />
                    <SPLIT distance="225" swimtime="00:03:05.07" />
                    <SPLIT distance="250" swimtime="00:03:26.38" />
                    <SPLIT distance="275" swimtime="00:03:47.81" />
                    <SPLIT distance="300" swimtime="00:04:09.11" />
                    <SPLIT distance="325" swimtime="00:04:30.63" />
                    <SPLIT distance="350" swimtime="00:04:51.86" />
                    <SPLIT distance="375" swimtime="00:05:11.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="106730" name="Pregel">
          <CONTACT email="alkonter@gmail.com" name="Liubavin Viktor" />
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Viktor" gender="M" lastname="Liubavin" nation="RUS" athleteid="106861">
              <RESULTS>
                <RESULT eventid="98798" points="377" reactiontime="+80" swimtime="00:00:28.03" resultid="106862" heatid="110606" lane="7" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="291" reactiontime="+96" swimtime="00:11:08.72" resultid="106863" heatid="110636" lane="7" entrytime="00:10:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="75" swimtime="00:00:57.62" />
                    <SPLIT distance="100" swimtime="00:01:18.14" />
                    <SPLIT distance="125" swimtime="00:01:38.49" />
                    <SPLIT distance="150" swimtime="00:01:59.47" />
                    <SPLIT distance="175" swimtime="00:02:20.69" />
                    <SPLIT distance="200" swimtime="00:02:41.94" />
                    <SPLIT distance="225" swimtime="00:03:02.39" />
                    <SPLIT distance="250" swimtime="00:03:23.64" />
                    <SPLIT distance="275" swimtime="00:03:44.64" />
                    <SPLIT distance="300" swimtime="00:04:06.24" />
                    <SPLIT distance="325" swimtime="00:04:26.84" />
                    <SPLIT distance="350" swimtime="00:04:48.08" />
                    <SPLIT distance="375" swimtime="00:05:08.98" />
                    <SPLIT distance="400" swimtime="00:05:29.99" />
                    <SPLIT distance="425" swimtime="00:05:51.54" />
                    <SPLIT distance="450" swimtime="00:06:12.66" />
                    <SPLIT distance="475" swimtime="00:06:33.67" />
                    <SPLIT distance="500" swimtime="00:06:55.08" />
                    <SPLIT distance="525" swimtime="00:07:16.45" />
                    <SPLIT distance="550" swimtime="00:07:37.62" />
                    <SPLIT distance="575" swimtime="00:07:58.71" />
                    <SPLIT distance="600" swimtime="00:08:19.94" />
                    <SPLIT distance="625" swimtime="00:08:41.29" />
                    <SPLIT distance="650" swimtime="00:09:02.90" />
                    <SPLIT distance="675" swimtime="00:09:24.64" />
                    <SPLIT distance="700" swimtime="00:09:45.91" />
                    <SPLIT distance="725" swimtime="00:10:07.03" />
                    <SPLIT distance="750" swimtime="00:10:28.10" />
                    <SPLIT distance="775" swimtime="00:10:49.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="328" reactiontime="+86" swimtime="00:02:54.67" resultid="106864" heatid="110668" lane="5" entrytime="00:03:03.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.60" />
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                    <SPLIT distance="75" swimtime="00:01:01.57" />
                    <SPLIT distance="100" swimtime="00:01:24.60" />
                    <SPLIT distance="125" swimtime="00:01:46.81" />
                    <SPLIT distance="150" swimtime="00:02:09.69" />
                    <SPLIT distance="175" swimtime="00:02:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="383" reactiontime="+84" swimtime="00:01:01.86" resultid="106865" heatid="110685" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.66" />
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="75" swimtime="00:00:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="364" reactiontime="+82" swimtime="00:01:17.84" resultid="106866" heatid="110732" lane="8" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.93" />
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="75" swimtime="00:00:57.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="334" reactiontime="+88" swimtime="00:02:23.10" resultid="106867" heatid="110775" lane="1" entrytime="00:02:22.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.82" />
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="75" swimtime="00:00:51.28" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="125" swimtime="00:01:28.63" />
                    <SPLIT distance="150" swimtime="00:01:47.51" />
                    <SPLIT distance="175" swimtime="00:02:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="198" swimtime="00:01:23.03" resultid="106868" heatid="110801" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.52" />
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="75" swimtime="00:00:59.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="379" swimtime="00:00:34.88" resultid="106869" heatid="110830" lane="6" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Vadim" gender="M" lastname="Ezhkov" nation="RUS" athleteid="106855">
              <RESULTS>
                <RESULT eventid="98988" points="270" swimtime="00:01:18.35" resultid="106856" heatid="110700" lane="9" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.68" />
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="75" swimtime="00:00:59.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="322" swimtime="00:01:21.10" resultid="106857" heatid="110731" lane="6" entrytime="00:01:21.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.00" />
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="75" swimtime="00:00:58.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="282" reactiontime="+74" swimtime="00:02:31.39" resultid="106858" heatid="110774" lane="8" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.95" />
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="75" swimtime="00:00:52.40" />
                    <SPLIT distance="100" swimtime="00:01:11.73" />
                    <SPLIT distance="125" swimtime="00:01:31.40" />
                    <SPLIT distance="150" swimtime="00:01:51.44" />
                    <SPLIT distance="175" swimtime="00:02:11.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="343" reactiontime="+54" swimtime="00:00:36.07" resultid="106859" heatid="110830" lane="7" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="267" swimtime="00:05:29.26" resultid="106860" heatid="110846" lane="9" entrytime="00:05:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.63" />
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="75" swimtime="00:00:56.02" />
                    <SPLIT distance="100" swimtime="00:01:16.35" />
                    <SPLIT distance="125" swimtime="00:01:36.78" />
                    <SPLIT distance="150" swimtime="00:01:57.77" />
                    <SPLIT distance="175" swimtime="00:02:18.70" />
                    <SPLIT distance="200" swimtime="00:02:39.97" />
                    <SPLIT distance="225" swimtime="00:03:01.16" />
                    <SPLIT distance="250" swimtime="00:03:22.61" />
                    <SPLIT distance="275" swimtime="00:03:44.12" />
                    <SPLIT distance="300" swimtime="00:04:05.74" />
                    <SPLIT distance="325" swimtime="00:04:26.82" />
                    <SPLIT distance="350" swimtime="00:04:48.34" />
                    <SPLIT distance="375" swimtime="00:05:09.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Vitalii" gender="M" lastname="Avdeev" nation="RUS" athleteid="106805">
              <RESULTS>
                <RESULT eventid="98798" points="176" swimtime="00:00:36.12" resultid="106806" heatid="110599" lane="9" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="141" reactiontime="+99" swimtime="00:03:30.24" resultid="106807" heatid="110620" lane="5" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.92" />
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                    <SPLIT distance="75" swimtime="00:01:13.90" />
                    <SPLIT distance="100" swimtime="00:01:45.83" />
                    <SPLIT distance="125" swimtime="00:02:15.33" />
                    <SPLIT distance="150" swimtime="00:02:45.72" />
                    <SPLIT distance="175" swimtime="00:03:08.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="186" reactiontime="+97" swimtime="00:01:18.62" resultid="106808" heatid="110680" lane="5" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.35" />
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="75" swimtime="00:00:59.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="118" reactiontime="+104" swimtime="00:03:41.19" resultid="106809" heatid="110711" lane="1" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.34" />
                    <SPLIT distance="50" swimtime="00:00:47.51" />
                    <SPLIT distance="75" swimtime="00:01:15.55" />
                    <SPLIT distance="100" swimtime="00:01:44.89" />
                    <SPLIT distance="125" swimtime="00:02:14.89" />
                    <SPLIT distance="150" swimtime="00:02:45.02" />
                    <SPLIT distance="175" swimtime="00:03:14.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="201" reactiontime="+97" swimtime="00:00:37.17" resultid="106810" heatid="110743" lane="7" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="151" reactiontime="+109" swimtime="00:01:30.78" resultid="106811" heatid="110799" lane="5" entrytime="00:01:37.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.83" />
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="75" swimtime="00:01:03.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Grigorii" gender="M" lastname="Lopin" nation="RUS" athleteid="106843">
              <RESULTS>
                <RESULT eventid="98798" points="305" reactiontime="+87" swimtime="00:00:30.07" resultid="106844" heatid="110602" lane="8" entrytime="00:00:31.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="252" reactiontime="+102" swimtime="00:11:41.57" resultid="106845" heatid="110637" lane="2" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.31" />
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="75" swimtime="00:00:58.27" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="125" swimtime="00:01:40.24" />
                    <SPLIT distance="150" swimtime="00:02:01.83" />
                    <SPLIT distance="175" swimtime="00:02:24.15" />
                    <SPLIT distance="200" swimtime="00:02:46.40" />
                    <SPLIT distance="225" swimtime="00:03:08.86" />
                    <SPLIT distance="250" swimtime="00:03:31.25" />
                    <SPLIT distance="275" swimtime="00:03:53.59" />
                    <SPLIT distance="300" swimtime="00:04:15.74" />
                    <SPLIT distance="325" swimtime="00:04:38.18" />
                    <SPLIT distance="350" swimtime="00:05:00.00" />
                    <SPLIT distance="375" swimtime="00:05:22.28" />
                    <SPLIT distance="400" swimtime="00:05:44.56" />
                    <SPLIT distance="425" swimtime="00:06:06.56" />
                    <SPLIT distance="450" swimtime="00:06:29.01" />
                    <SPLIT distance="475" swimtime="00:06:51.36" />
                    <SPLIT distance="500" swimtime="00:07:13.89" />
                    <SPLIT distance="525" swimtime="00:07:36.78" />
                    <SPLIT distance="550" swimtime="00:07:59.25" />
                    <SPLIT distance="575" swimtime="00:08:21.67" />
                    <SPLIT distance="600" swimtime="00:08:44.85" />
                    <SPLIT distance="625" swimtime="00:09:06.99" />
                    <SPLIT distance="650" swimtime="00:09:28.91" />
                    <SPLIT distance="675" swimtime="00:09:51.15" />
                    <SPLIT distance="700" swimtime="00:10:14.25" />
                    <SPLIT distance="725" swimtime="00:10:36.77" />
                    <SPLIT distance="750" swimtime="00:10:59.36" />
                    <SPLIT distance="775" swimtime="00:11:21.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="266" reactiontime="+96" swimtime="00:03:07.13" resultid="106846" heatid="110667" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.44" />
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="75" swimtime="00:01:05.84" />
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                    <SPLIT distance="125" swimtime="00:01:54.07" />
                    <SPLIT distance="150" swimtime="00:02:18.86" />
                    <SPLIT distance="175" swimtime="00:02:43.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="285" reactiontime="+83" swimtime="00:01:24.48" resultid="106847" heatid="110730" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.04" />
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                    <SPLIT distance="75" swimtime="00:01:02.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="220" reactiontime="+95" swimtime="00:06:29.67" resultid="106848" heatid="110789" lane="4" entrytime="00:06:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.35" />
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                    <SPLIT distance="75" swimtime="00:01:11.68" />
                    <SPLIT distance="100" swimtime="00:01:37.27" />
                    <SPLIT distance="125" swimtime="00:02:03.79" />
                    <SPLIT distance="150" swimtime="00:02:29.93" />
                    <SPLIT distance="175" swimtime="00:02:55.43" />
                    <SPLIT distance="200" swimtime="00:03:20.62" />
                    <SPLIT distance="225" swimtime="00:03:45.77" />
                    <SPLIT distance="250" swimtime="00:04:11.57" />
                    <SPLIT distance="275" swimtime="00:04:36.84" />
                    <SPLIT distance="300" swimtime="00:05:03.54" />
                    <SPLIT distance="325" swimtime="00:05:25.40" />
                    <SPLIT distance="350" swimtime="00:05:48.37" />
                    <SPLIT distance="375" swimtime="00:06:08.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="300" swimtime="00:00:37.69" resultid="106849" heatid="110828" lane="6" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="250" reactiontime="+95" swimtime="00:05:36.48" resultid="106850" heatid="110848" lane="4" entrytime="00:05:44.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:56.50" />
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="75" swimtime="00:01:38.73" />
                    <SPLIT distance="100" swimtime="00:01:17.32" />
                    <SPLIT distance="150" swimtime="00:02:00.56" />
                    <SPLIT distance="175" swimtime="00:02:21.84" />
                    <SPLIT distance="200" swimtime="00:02:43.99" />
                    <SPLIT distance="225" swimtime="00:03:05.78" />
                    <SPLIT distance="250" swimtime="00:03:27.86" />
                    <SPLIT distance="275" swimtime="00:03:49.66" />
                    <SPLIT distance="300" swimtime="00:04:11.71" />
                    <SPLIT distance="325" swimtime="00:04:33.24" />
                    <SPLIT distance="350" swimtime="00:04:55.66" />
                    <SPLIT distance="375" swimtime="00:05:17.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Olga" gender="F" lastname="Tikhomirova" nation="RUS" athleteid="106757">
              <RESULTS>
                <RESULT eventid="98814" status="WDR" swimtime="00:00:00.00" resultid="106758" entrytime="00:03:39.00" />
                <RESULT eventid="106294" status="WDR" swimtime="00:00:00.00" resultid="106759" entrytime="00:00:44.50" />
                <RESULT eventid="98972" status="WDR" swimtime="00:00:00.00" resultid="106760" entrytime="00:01:35.50" />
                <RESULT eventid="99314" status="WDR" swimtime="00:00:00.00" resultid="106761" entrytime="00:01:39.00" />
                <RESULT eventid="99266" status="WDR" swimtime="00:00:00.00" resultid="106762" entrytime="00:07:59.00" />
                <RESULT eventid="99344" status="WDR" swimtime="00:00:00.00" resultid="106763" entrytime="00:01:39.50" />
                <RESULT eventid="99409" status="WDR" swimtime="00:00:00.00" resultid="106764" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Tatiana" gender="F" lastname="Logvinova" nation="RUS" athleteid="106765">
              <RESULTS>
                <RESULT eventid="106294" status="DNS" swimtime="00:00:00.00" resultid="106766" heatid="110647" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="98972" points="215" swimtime="00:01:34.47" resultid="106767" heatid="110692" lane="9" entrytime="00:01:34.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.52" />
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                    <SPLIT distance="75" swimtime="00:01:12.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="245" reactiontime="+87" swimtime="00:01:39.60" resultid="106768" heatid="110722" lane="4" entrytime="00:01:41.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.65" />
                    <SPLIT distance="50" swimtime="00:00:47.48" />
                    <SPLIT distance="75" swimtime="00:01:13.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="157" swimtime="00:00:45.17" resultid="106769" heatid="110737" lane="0" entrytime="00:00:44.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="106" swimtime="00:01:55.29" resultid="106770" heatid="110794" lane="6" entrytime="00:01:39.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.89" />
                    <SPLIT distance="50" swimtime="00:00:53.55" />
                    <SPLIT distance="75" swimtime="00:01:23.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="263" reactiontime="+113" swimtime="00:00:44.93" resultid="106771" heatid="110819" lane="3" entrytime="00:00:46.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Sergei" gender="M" lastname="Mikhaylov" nation="RUS" athleteid="106829">
              <RESULTS>
                <RESULT eventid="98798" points="117" swimtime="00:00:41.42" resultid="106830" heatid="110598" lane="9" entrytime="00:00:39.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="155" reactiontime="+105" swimtime="00:26:17.97" resultid="106831" heatid="110643" lane="7" entrytime="00:26:37.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.20" />
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                    <SPLIT distance="75" swimtime="00:01:10.23" />
                    <SPLIT distance="100" swimtime="00:01:35.44" />
                    <SPLIT distance="125" swimtime="00:02:01.56" />
                    <SPLIT distance="150" swimtime="00:02:27.33" />
                    <SPLIT distance="175" swimtime="00:02:53.72" />
                    <SPLIT distance="200" swimtime="00:03:20.23" />
                    <SPLIT distance="225" swimtime="00:03:45.73" />
                    <SPLIT distance="250" swimtime="00:04:11.77" />
                    <SPLIT distance="275" swimtime="00:04:37.87" />
                    <SPLIT distance="300" swimtime="00:05:04.10" />
                    <SPLIT distance="325" swimtime="00:05:30.58" />
                    <SPLIT distance="350" swimtime="00:05:56.80" />
                    <SPLIT distance="375" swimtime="00:06:23.46" />
                    <SPLIT distance="400" swimtime="00:06:48.88" />
                    <SPLIT distance="425" swimtime="00:07:15.91" />
                    <SPLIT distance="450" swimtime="00:07:42.15" />
                    <SPLIT distance="475" swimtime="00:08:08.46" />
                    <SPLIT distance="500" swimtime="00:08:35.02" />
                    <SPLIT distance="525" swimtime="00:09:00.21" />
                    <SPLIT distance="550" swimtime="00:09:27.01" />
                    <SPLIT distance="575" swimtime="00:09:52.72" />
                    <SPLIT distance="600" swimtime="00:10:19.48" />
                    <SPLIT distance="625" swimtime="00:10:45.90" />
                    <SPLIT distance="650" swimtime="00:11:12.63" />
                    <SPLIT distance="675" swimtime="00:11:38.65" />
                    <SPLIT distance="700" swimtime="00:12:05.69" />
                    <SPLIT distance="725" swimtime="00:12:32.13" />
                    <SPLIT distance="750" swimtime="00:12:58.97" />
                    <SPLIT distance="775" swimtime="00:13:24.86" />
                    <SPLIT distance="800" swimtime="00:13:51.66" />
                    <SPLIT distance="825" swimtime="00:14:18.50" />
                    <SPLIT distance="850" swimtime="00:14:45.21" />
                    <SPLIT distance="875" swimtime="00:15:11.47" />
                    <SPLIT distance="900" swimtime="00:15:38.12" />
                    <SPLIT distance="925" swimtime="00:16:04.94" />
                    <SPLIT distance="950" swimtime="00:16:31.80" />
                    <SPLIT distance="975" swimtime="00:16:57.79" />
                    <SPLIT distance="1000" swimtime="00:17:24.77" />
                    <SPLIT distance="1025" swimtime="00:17:52.34" />
                    <SPLIT distance="1050" swimtime="00:18:19.49" />
                    <SPLIT distance="1075" swimtime="00:18:46.14" />
                    <SPLIT distance="1100" swimtime="00:19:12.38" />
                    <SPLIT distance="1125" swimtime="00:19:38.97" />
                    <SPLIT distance="1150" swimtime="00:20:05.92" />
                    <SPLIT distance="1175" swimtime="00:20:32.59" />
                    <SPLIT distance="1200" swimtime="00:20:59.83" />
                    <SPLIT distance="1225" swimtime="00:21:27.11" />
                    <SPLIT distance="1250" swimtime="00:21:52.85" />
                    <SPLIT distance="1275" swimtime="00:22:19.67" />
                    <SPLIT distance="1300" swimtime="00:22:46.73" />
                    <SPLIT distance="1325" swimtime="00:23:13.78" />
                    <SPLIT distance="1350" swimtime="00:23:40.28" />
                    <SPLIT distance="1375" swimtime="00:24:06.97" />
                    <SPLIT distance="1400" swimtime="00:24:33.94" />
                    <SPLIT distance="1425" swimtime="00:25:00.35" />
                    <SPLIT distance="1450" swimtime="00:25:27.07" />
                    <SPLIT distance="1475" swimtime="00:25:53.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="119" swimtime="00:01:31.15" resultid="106832" heatid="110680" lane="0" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.23" />
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="75" swimtime="00:01:07.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="146" reactiontime="+103" swimtime="00:03:08.49" resultid="106833" heatid="110770" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.84" />
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                    <SPLIT distance="75" swimtime="00:01:06.91" />
                    <SPLIT distance="100" swimtime="00:01:31.71" />
                    <SPLIT distance="125" swimtime="00:01:56.83" />
                    <SPLIT distance="150" swimtime="00:02:22.44" />
                    <SPLIT distance="175" swimtime="00:02:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4" eventid="99473" reactiontime="+107" status="DSQ" swimtime="00:00:00.00" resultid="106834" heatid="110850" lane="8" entrytime="00:06:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Elena" gender="F" lastname="Mekhteleva" nation="RUS" athleteid="106784">
              <RESULTS>
                <RESULT eventid="98940" points="455" reactiontime="+98" swimtime="00:02:54.95" resultid="106785" heatid="110664" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.37" />
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="75" swimtime="00:01:01.38" />
                    <SPLIT distance="100" swimtime="00:01:23.64" />
                    <SPLIT distance="125" swimtime="00:01:46.19" />
                    <SPLIT distance="150" swimtime="00:02:09.07" />
                    <SPLIT distance="175" swimtime="00:02:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="501" reactiontime="+91" swimtime="00:01:18.50" resultid="106786" heatid="110725" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.29" />
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="75" swimtime="00:00:57.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="403" swimtime="00:00:32.98" resultid="106787" heatid="110739" lane="6" entrytime="00:00:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="502" reactiontime="+78" swimtime="00:00:36.23" resultid="106788" heatid="110823" lane="8" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Aleksandr" gender="M" lastname="Smirnov" nation="RUS" athleteid="106876">
              <RESULTS>
                <RESULT eventid="106256" points="391" reactiontime="+81" swimtime="00:19:19.07" resultid="106877" heatid="110641" lane="7" entrytime="00:19:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.88" />
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="75" swimtime="00:00:52.74" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="125" swimtime="00:01:30.80" />
                    <SPLIT distance="150" swimtime="00:01:50.07" />
                    <SPLIT distance="175" swimtime="00:02:09.39" />
                    <SPLIT distance="200" swimtime="00:02:28.64" />
                    <SPLIT distance="225" swimtime="00:02:48.02" />
                    <SPLIT distance="250" swimtime="00:03:07.47" />
                    <SPLIT distance="275" swimtime="00:03:27.03" />
                    <SPLIT distance="300" swimtime="00:03:46.31" />
                    <SPLIT distance="325" swimtime="00:04:05.46" />
                    <SPLIT distance="350" swimtime="00:04:24.78" />
                    <SPLIT distance="375" swimtime="00:04:44.02" />
                    <SPLIT distance="400" swimtime="00:05:03.44" />
                    <SPLIT distance="425" swimtime="00:05:23.05" />
                    <SPLIT distance="450" swimtime="00:05:42.45" />
                    <SPLIT distance="475" swimtime="00:06:01.77" />
                    <SPLIT distance="500" swimtime="00:06:21.18" />
                    <SPLIT distance="525" swimtime="00:06:40.63" />
                    <SPLIT distance="550" swimtime="00:07:00.08" />
                    <SPLIT distance="575" swimtime="00:07:19.41" />
                    <SPLIT distance="600" swimtime="00:07:38.87" />
                    <SPLIT distance="625" swimtime="00:07:58.45" />
                    <SPLIT distance="650" swimtime="00:08:18.18" />
                    <SPLIT distance="675" swimtime="00:08:37.62" />
                    <SPLIT distance="700" swimtime="00:08:57.27" />
                    <SPLIT distance="725" swimtime="00:09:16.81" />
                    <SPLIT distance="750" swimtime="00:09:36.54" />
                    <SPLIT distance="775" swimtime="00:09:55.89" />
                    <SPLIT distance="800" swimtime="00:10:15.73" />
                    <SPLIT distance="825" swimtime="00:10:35.51" />
                    <SPLIT distance="850" swimtime="00:10:55.31" />
                    <SPLIT distance="875" swimtime="00:11:14.80" />
                    <SPLIT distance="900" swimtime="00:11:34.32" />
                    <SPLIT distance="925" swimtime="00:11:53.88" />
                    <SPLIT distance="950" swimtime="00:12:13.47" />
                    <SPLIT distance="975" swimtime="00:12:33.17" />
                    <SPLIT distance="1000" swimtime="00:12:52.77" />
                    <SPLIT distance="1025" swimtime="00:13:12.22" />
                    <SPLIT distance="1050" swimtime="00:13:31.86" />
                    <SPLIT distance="1075" swimtime="00:13:51.46" />
                    <SPLIT distance="1100" swimtime="00:14:11.05" />
                    <SPLIT distance="1125" swimtime="00:14:30.70" />
                    <SPLIT distance="1150" swimtime="00:14:50.26" />
                    <SPLIT distance="1175" swimtime="00:15:09.88" />
                    <SPLIT distance="1200" swimtime="00:15:29.74" />
                    <SPLIT distance="1225" swimtime="00:15:49.42" />
                    <SPLIT distance="1250" swimtime="00:16:08.80" />
                    <SPLIT distance="1275" swimtime="00:16:28.18" />
                    <SPLIT distance="1300" swimtime="00:16:47.39" />
                    <SPLIT distance="1325" swimtime="00:17:06.56" />
                    <SPLIT distance="1350" swimtime="00:17:25.66" />
                    <SPLIT distance="1375" swimtime="00:17:44.83" />
                    <SPLIT distance="1400" swimtime="00:18:04.25" />
                    <SPLIT distance="1425" swimtime="00:18:23.85" />
                    <SPLIT distance="1450" swimtime="00:18:42.90" />
                    <SPLIT distance="1475" swimtime="00:19:01.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="379" reactiontime="+86" swimtime="00:01:02.07" resultid="106878" heatid="110686" lane="8" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.12" />
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="75" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="380" swimtime="00:02:17.09" resultid="106879" heatid="110776" lane="9" entrytime="00:02:18.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.07" />
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="75" swimtime="00:00:49.49" />
                    <SPLIT distance="100" swimtime="00:01:07.43" />
                    <SPLIT distance="125" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:01:42.90" />
                    <SPLIT distance="175" swimtime="00:02:00.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="106880" heatid="110830" lane="2" entrytime="00:00:36.50" />
                <RESULT eventid="99473" points="393" swimtime="00:04:49.65" resultid="106881" heatid="110844" lane="0" entrytime="00:04:52.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.78" />
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="75" swimtime="00:00:51.46" />
                    <SPLIT distance="100" swimtime="00:01:10.13" />
                    <SPLIT distance="125" swimtime="00:01:28.71" />
                    <SPLIT distance="150" swimtime="00:01:47.55" />
                    <SPLIT distance="175" swimtime="00:02:05.87" />
                    <SPLIT distance="200" swimtime="00:02:24.39" />
                    <SPLIT distance="225" swimtime="00:02:42.65" />
                    <SPLIT distance="250" swimtime="00:03:01.23" />
                    <SPLIT distance="275" swimtime="00:03:19.34" />
                    <SPLIT distance="300" swimtime="00:03:37.89" />
                    <SPLIT distance="325" swimtime="00:03:56.25" />
                    <SPLIT distance="350" swimtime="00:04:14.58" />
                    <SPLIT distance="375" swimtime="00:04:32.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Yuri" gender="M" lastname="Yakovenko" nation="RUS" athleteid="106818">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="106819" heatid="110599" lane="0" entrytime="00:00:36.50" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="106820" heatid="110653" lane="7" entrytime="00:00:46.50" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="106821" heatid="110728" lane="6" entrytime="00:01:44.50" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="106822" heatid="110828" lane="1" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Elena" gender="F" lastname="Kolyadina" nation="RUS" athleteid="106745">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="106746" heatid="110589" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="106747" heatid="110615" lane="6" entrytime="00:03:25.00" />
                <RESULT eventid="98940" status="DNS" swimtime="00:00:00.00" resultid="106748" heatid="110662" lane="3" entrytime="00:03:35.00" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="106749" heatid="110673" lane="2" entrytime="00:01:22.00" />
                <RESULT eventid="99089" status="DNS" swimtime="00:00:00.00" resultid="106750" heatid="110723" lane="6" entrytime="00:01:36.50" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="106751" heatid="110821" lane="9" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Olga" gender="F" lastname="Sulimova" nation="RUS" athleteid="106772">
              <RESULTS>
                <RESULT eventid="98777" points="221" reactiontime="+106" swimtime="00:00:38.40" resultid="106773" heatid="110588" lane="8" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="190" reactiontime="+111" swimtime="00:01:28.48" resultid="106774" heatid="110672" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.12" />
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="75" swimtime="00:01:04.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="125" reactiontime="+104" swimtime="00:00:48.67" resultid="106775" heatid="110736" lane="4" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="179" reactiontime="+102" swimtime="00:03:16.39" resultid="106776" heatid="110765" lane="6" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.12" />
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                    <SPLIT distance="75" swimtime="00:01:08.58" />
                    <SPLIT distance="100" swimtime="00:01:34.20" />
                    <SPLIT distance="125" swimtime="00:02:00.14" />
                    <SPLIT distance="150" swimtime="00:02:26.38" />
                    <SPLIT distance="175" swimtime="00:02:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="167" swimtime="00:00:52.21" resultid="106777" heatid="110819" lane="9" entrytime="00:00:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Sergei" gender="M" lastname="Karakchiev" nation="RUS" athleteid="106882">
              <RESULTS>
                <RESULT eventid="98830" points="354" reactiontime="+83" swimtime="00:02:34.86" resultid="106883" heatid="110625" lane="3" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.78" />
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="75" swimtime="00:00:51.40" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="125" swimtime="00:01:32.91" />
                    <SPLIT distance="150" swimtime="00:01:56.08" />
                    <SPLIT distance="175" swimtime="00:02:16.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="334" reactiontime="+75" swimtime="00:00:32.02" resultid="106884" heatid="110657" lane="6" entrytime="00:00:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="402" reactiontime="+70" swimtime="00:01:08.60" resultid="106885" heatid="110703" lane="2" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.37" />
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="75" swimtime="00:00:51.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="347" reactiontime="+79" swimtime="00:01:09.61" resultid="106886" heatid="110762" lane="0" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.29" />
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="75" swimtime="00:00:51.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="333" reactiontime="+78" swimtime="00:02:32.28" resultid="106887" heatid="110814" lane="7" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.80" />
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="75" swimtime="00:00:54.27" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="125" swimtime="00:01:33.83" />
                    <SPLIT distance="150" swimtime="00:01:53.64" />
                    <SPLIT distance="175" swimtime="00:02:13.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Igor" gender="M" lastname="Geyt" nation="RUS" athleteid="106870">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="106871" heatid="110602" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="98956" points="273" reactiontime="+84" swimtime="00:03:05.65" resultid="106872" heatid="110667" lane="5" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.42" />
                    <SPLIT distance="50" swimtime="00:00:42.70" />
                    <SPLIT distance="75" swimtime="00:01:06.52" />
                    <SPLIT distance="100" swimtime="00:01:31.08" />
                    <SPLIT distance="125" swimtime="00:01:54.91" />
                    <SPLIT distance="150" swimtime="00:02:18.89" />
                    <SPLIT distance="175" swimtime="00:02:42.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="259" reactiontime="+112" swimtime="00:01:19.46" resultid="106873" heatid="110699" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="75" swimtime="00:01:01.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="284" reactiontime="+88" swimtime="00:01:24.53" resultid="106874" heatid="110730" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.82" />
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="75" swimtime="00:01:01.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="283" reactiontime="+69" swimtime="00:00:38.43" resultid="106875" heatid="110828" lane="4" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Elena" gender="F" lastname="Dautova" nation="RUS" athleteid="106778">
              <RESULTS>
                <RESULT eventid="98777" points="395" reactiontime="+95" swimtime="00:00:31.66" resultid="106779" heatid="110591" lane="0" entrytime="00:00:32.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="323" reactiontime="+81" swimtime="00:00:37.39" resultid="106780" heatid="110649" lane="1" entrytime="00:00:38.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="357" swimtime="00:01:11.73" resultid="106781" heatid="110674" lane="4" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.28" />
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="75" swimtime="00:00:53.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="252" reactiontime="+62" swimtime="00:01:27.04" resultid="106782" heatid="110755" lane="6" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.01" />
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                    <SPLIT distance="75" swimtime="00:01:05.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="234" reactiontime="+75" swimtime="00:03:13.32" resultid="106783" heatid="110807" lane="5" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.84" />
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                    <SPLIT distance="75" swimtime="00:01:09.22" />
                    <SPLIT distance="100" swimtime="00:01:33.41" />
                    <SPLIT distance="125" swimtime="00:01:59.02" />
                    <SPLIT distance="150" swimtime="00:02:24.35" />
                    <SPLIT distance="175" swimtime="00:02:49.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-01-01" firstname="Luiza" gender="F" lastname="Shcherbich" nation="RUS" athleteid="106740">
              <RESULTS>
                <RESULT eventid="98777" points="51" reactiontime="+113" swimtime="00:01:02.31" resultid="106741" heatid="110586" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="39" reactiontime="+133" swimtime="00:02:29.44" resultid="106742" heatid="110671" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.37" />
                    <SPLIT distance="50" swimtime="00:01:07.40" />
                    <SPLIT distance="75" swimtime="00:01:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="58" reactiontime="+119" swimtime="00:02:40.69" resultid="106743" heatid="110720" lane="5" entrytime="00:05:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.22" />
                    <SPLIT distance="50" swimtime="00:01:16.27" />
                    <SPLIT distance="75" swimtime="00:01:58.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="68" reactiontime="+119" swimtime="00:01:10.48" resultid="106744" heatid="110817" lane="5" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Liudmila" gender="F" lastname="Kokhan" nation="RUS" athleteid="106789">
              <RESULTS>
                <RESULT eventid="98777" points="353" swimtime="00:00:32.86" resultid="106790" heatid="110591" lane="9" entrytime="00:00:32.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="208" swimtime="00:03:47.10" resultid="106791" heatid="110662" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.62" />
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                    <SPLIT distance="75" swimtime="00:01:16.88" />
                    <SPLIT distance="100" swimtime="00:01:45.91" />
                    <SPLIT distance="125" swimtime="00:02:15.44" />
                    <SPLIT distance="150" swimtime="00:02:45.27" />
                    <SPLIT distance="175" swimtime="00:03:15.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="229" reactiontime="+87" swimtime="00:01:32.52" resultid="106792" heatid="110692" lane="8" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.46" />
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="75" swimtime="00:01:11.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="229" swimtime="00:01:41.80" resultid="106793" heatid="110723" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.90" />
                    <SPLIT distance="50" swimtime="00:00:47.71" />
                    <SPLIT distance="75" swimtime="00:01:14.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="200" reactiontime="+95" swimtime="00:00:41.64" resultid="106794" heatid="110737" lane="2" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="106795" heatid="110819" lane="2" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Regina" gender="F" lastname="Sych" nation="RUS" athleteid="106796">
              <RESULTS>
                <RESULT eventid="98777" points="649" reactiontime="+86" swimtime="00:00:26.84" resultid="106797" heatid="110593" lane="1" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="106798" heatid="110618" lane="2" entrytime="00:02:40.00" />
                <RESULT eventid="106294" points="488" reactiontime="+75" swimtime="00:00:32.59" resultid="106799" heatid="110650" lane="9" entrytime="00:00:34.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="647" reactiontime="+60" swimtime="00:00:58.86" resultid="106800" heatid="110676" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.89" />
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="75" swimtime="00:00:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="573" reactiontime="+75" swimtime="00:00:29.35" resultid="106801" heatid="110740" lane="8" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="106802" heatid="110768" lane="6" entrytime="00:02:19.00" />
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="106803" heatid="110796" lane="7" entrytime="00:01:13.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="106804" heatid="110823" lane="0" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Sergei" gender="M" lastname="Ryabov" nation="RUS" athleteid="106835">
              <RESULTS>
                <RESULT eventid="98798" status="WDR" swimtime="00:00:00.00" resultid="106836" entrytime="00:00:31.50" />
                <RESULT eventid="106256" status="WDR" swimtime="00:00:00.00" resultid="106837" entrytime="00:23:39.50" />
                <RESULT eventid="106277" status="WDR" swimtime="00:00:00.00" resultid="106838" entrytime="00:01:10.50" />
                <RESULT eventid="99170" status="WDR" swimtime="00:00:00.00" resultid="106839" entrytime="00:00:34.50" />
                <RESULT eventid="99218" status="WDR" swimtime="00:00:00.00" resultid="106840" entrytime="00:02:42.50" />
                <RESULT eventid="99425" status="WDR" swimtime="00:00:00.00" resultid="106841" entrytime="00:00:41.30" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="106842" entrytime="00:05:39.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Aleksandr" gender="M" lastname="Zelenov" nation="RUS" athleteid="106812">
              <RESULTS>
                <RESULT eventid="98798" points="99" reactiontime="+127" swimtime="00:00:43.69" resultid="106813" heatid="110596" lane="7" entrytime="00:00:42.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="102" reactiontime="+108" swimtime="00:15:47.01" resultid="106814" heatid="110638" lane="7" entrytime="00:15:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.15" />
                    <SPLIT distance="50" swimtime="00:00:49.65" />
                    <SPLIT distance="75" swimtime="00:01:18.13" />
                    <SPLIT distance="100" swimtime="00:01:47.84" />
                    <SPLIT distance="125" swimtime="00:02:17.31" />
                    <SPLIT distance="150" swimtime="00:02:47.40" />
                    <SPLIT distance="175" swimtime="00:03:17.63" />
                    <SPLIT distance="200" swimtime="00:03:47.50" />
                    <SPLIT distance="225" swimtime="00:04:17.76" />
                    <SPLIT distance="250" swimtime="00:04:47.92" />
                    <SPLIT distance="275" swimtime="00:05:17.68" />
                    <SPLIT distance="300" swimtime="00:05:47.83" />
                    <SPLIT distance="325" swimtime="00:06:18.19" />
                    <SPLIT distance="350" swimtime="00:06:48.38" />
                    <SPLIT distance="375" swimtime="00:07:18.71" />
                    <SPLIT distance="400" swimtime="00:07:48.93" />
                    <SPLIT distance="425" swimtime="00:08:18.93" />
                    <SPLIT distance="450" swimtime="00:08:49.19" />
                    <SPLIT distance="475" swimtime="00:09:19.60" />
                    <SPLIT distance="500" swimtime="00:09:50.04" />
                    <SPLIT distance="525" swimtime="00:10:20.01" />
                    <SPLIT distance="550" swimtime="00:10:50.95" />
                    <SPLIT distance="575" swimtime="00:11:20.89" />
                    <SPLIT distance="600" swimtime="00:11:51.25" />
                    <SPLIT distance="625" swimtime="00:12:20.83" />
                    <SPLIT distance="650" swimtime="00:12:50.97" />
                    <SPLIT distance="675" swimtime="00:13:20.68" />
                    <SPLIT distance="700" swimtime="00:13:50.28" />
                    <SPLIT distance="725" swimtime="00:14:20.11" />
                    <SPLIT distance="750" swimtime="00:14:49.95" />
                    <SPLIT distance="775" swimtime="00:15:18.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="91" reactiontime="+123" swimtime="00:01:39.65" resultid="106815" heatid="110679" lane="1" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.32" />
                    <SPLIT distance="50" swimtime="00:00:45.77" />
                    <SPLIT distance="75" swimtime="00:01:12.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="87" swimtime="00:03:43.62" resultid="106816" heatid="110769" lane="4" entrytime="00:03:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.86" />
                    <SPLIT distance="50" swimtime="00:00:47.42" />
                    <SPLIT distance="75" swimtime="00:01:15.44" />
                    <SPLIT distance="100" swimtime="00:01:45.53" />
                    <SPLIT distance="125" swimtime="00:02:15.55" />
                    <SPLIT distance="150" swimtime="00:02:45.62" />
                    <SPLIT distance="175" swimtime="00:03:15.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="99" reactiontime="+121" swimtime="00:07:38.55" resultid="106817" heatid="110851" lane="7" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.46" />
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                    <SPLIT distance="75" swimtime="00:01:16.86" />
                    <SPLIT distance="100" swimtime="00:01:45.95" />
                    <SPLIT distance="125" swimtime="00:02:15.90" />
                    <SPLIT distance="150" swimtime="00:02:45.99" />
                    <SPLIT distance="175" swimtime="00:03:16.05" />
                    <SPLIT distance="200" swimtime="00:03:46.20" />
                    <SPLIT distance="225" swimtime="00:04:16.35" />
                    <SPLIT distance="250" swimtime="00:04:45.59" />
                    <SPLIT distance="275" swimtime="00:05:14.92" />
                    <SPLIT distance="300" swimtime="00:05:44.37" />
                    <SPLIT distance="325" swimtime="00:06:13.42" />
                    <SPLIT distance="350" swimtime="00:06:43.13" />
                    <SPLIT distance="375" swimtime="00:07:12.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Ruslan" gender="M" lastname="Yakovenko" nation="RUS" athleteid="106888">
              <RESULTS>
                <RESULT eventid="98798" status="WDR" swimtime="00:00:00.00" resultid="106889" entrytime="00:00:30.00" />
                <RESULT eventid="106277" status="WDR" swimtime="00:00:00.00" resultid="106890" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Irina" gender="F" lastname="Titova" nation="RUS" athleteid="106752">
              <RESULTS>
                <RESULT eventid="98777" points="308" reactiontime="+101" swimtime="00:00:34.39" resultid="106753" heatid="110589" lane="7" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="310" swimtime="00:01:15.19" resultid="106754" heatid="110673" lane="4" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.67" />
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="106755" heatid="110767" lane="9" entrytime="00:02:47.00" />
                <RESULT eventid="99457" status="DNS" swimtime="00:00:00.00" resultid="106756" heatid="110840" lane="7" entrytime="00:05:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Aleksandr" gender="M" lastname="Tervinskii" nation="RUS" athleteid="106823">
              <RESULTS>
                <RESULT eventid="98798" points="219" reactiontime="+105" swimtime="00:00:33.58" resultid="106824" heatid="110600" lane="0" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="166" reactiontime="+84" swimtime="00:00:40.42" resultid="106825" heatid="110654" lane="8" entrytime="00:00:41.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="106826" heatid="110698" lane="8" entrytime="00:01:27.80" />
                <RESULT eventid="99091" points="200" reactiontime="+90" swimtime="00:01:35.07" resultid="106827" heatid="110729" lane="8" entrytime="00:01:36.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.41" />
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                    <SPLIT distance="75" swimtime="00:01:10.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="260" reactiontime="+85" swimtime="00:00:39.56" resultid="106828" heatid="110827" lane="8" entrytime="00:00:41.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Vitalii" gender="M" lastname="Galygin" nation="RUS" athleteid="106851">
              <RESULTS>
                <RESULT eventid="98924" points="172" reactiontime="+75" swimtime="00:00:39.91" resultid="106852" heatid="110655" lane="2" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="170" swimtime="00:00:39.35" resultid="106853" heatid="110744" lane="0" entrytime="00:00:35.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.79" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G3" eventid="99186" reactiontime="+85" status="DSQ" swimtime="00:00:00.00" resultid="106854" heatid="110759" lane="4" entrytime="00:01:25.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="175" reactiontime="+74" swimtime="00:02:41.53" resultid="106895" heatid="110716" lane="4" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.95" />
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                    <SPLIT distance="75" swimtime="00:01:01.20" />
                    <SPLIT distance="100" swimtime="00:01:22.85" />
                    <SPLIT distance="125" swimtime="00:01:40.02" />
                    <SPLIT distance="150" swimtime="00:02:01.67" />
                    <SPLIT distance="175" swimtime="00:02:20.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106843" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="106823" number="2" reactiontime="+6" />
                    <RELAYPOSITION athleteid="106805" number="3" />
                    <RELAYPOSITION athleteid="106818" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="220" swimtime="00:02:16.78" resultid="106899" heatid="110782" lane="0" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.51" />
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="75" swimtime="00:00:48.40" />
                    <SPLIT distance="100" swimtime="00:01:05.64" />
                    <SPLIT distance="125" swimtime="00:01:23.25" />
                    <SPLIT distance="150" swimtime="00:01:42.53" />
                    <SPLIT distance="175" swimtime="00:01:58.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106843" number="1" />
                    <RELAYPOSITION athleteid="106823" number="2" />
                    <RELAYPOSITION athleteid="106805" number="3" />
                    <RELAYPOSITION athleteid="106818" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="315" reactiontime="+75" swimtime="00:02:12.89" resultid="106896" heatid="110717" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.21" />
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="75" swimtime="00:00:48.89" />
                    <SPLIT distance="100" swimtime="00:01:08.65" />
                    <SPLIT distance="125" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:01:39.79" />
                    <SPLIT distance="175" swimtime="00:01:55.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106882" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="106855" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="106861" number="3" reactiontime="+13" />
                    <RELAYPOSITION athleteid="106851" number="4" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="382" reactiontime="+81" swimtime="00:01:53.75" resultid="106900" heatid="110782" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.47" />
                    <SPLIT distance="50" swimtime="00:00:27.29" />
                    <SPLIT distance="75" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:00:54.87" />
                    <SPLIT distance="125" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:25.41" />
                    <SPLIT distance="175" swimtime="00:01:38.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106882" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="106861" number="2" reactiontime="+4" />
                    <RELAYPOSITION athleteid="106870" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="106851" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="424" reactiontime="+71" swimtime="00:02:18.48" resultid="106891" heatid="110715" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.30" />
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="75" swimtime="00:00:55.42" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="125" swimtime="00:01:28.21" />
                    <SPLIT distance="150" swimtime="00:01:44.35" />
                    <SPLIT distance="175" swimtime="00:02:00.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106778" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="106784" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="106796" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="106752" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99234" points="173" reactiontime="+119" swimtime="00:02:49.10" resultid="106897" heatid="110780" lane="8" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.74" />
                    <SPLIT distance="50" swimtime="00:00:49.38" />
                    <SPLIT distance="75" swimtime="00:01:08.44" />
                    <SPLIT distance="100" swimtime="00:01:31.47" />
                    <SPLIT distance="125" swimtime="00:01:49.42" />
                    <SPLIT distance="150" swimtime="00:02:09.19" />
                    <SPLIT distance="175" swimtime="00:02:28.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106789" number="1" reactiontime="+119" />
                    <RELAYPOSITION athleteid="106745" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="106765" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="106772" number="4" reactiontime="+78" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="99234" points="435" reactiontime="+81" swimtime="00:02:04.37" resultid="106898" heatid="110780" lane="2" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.93" />
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="75" swimtime="00:00:47.65" />
                    <SPLIT distance="100" swimtime="00:01:03.05" />
                    <SPLIT distance="125" swimtime="00:01:16.42" />
                    <SPLIT distance="150" swimtime="00:01:30.76" />
                    <SPLIT distance="175" swimtime="00:01:46.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106778" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="106784" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="106796" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="106752" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="99036" points="209" reactiontime="+71" swimtime="00:02:55.15" resultid="106904" heatid="110715" lane="8" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.19" />
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                    <SPLIT distance="75" swimtime="00:01:07.51" />
                    <SPLIT distance="100" swimtime="00:01:32.16" />
                    <SPLIT distance="125" swimtime="00:01:53.40" />
                    <SPLIT distance="150" swimtime="00:02:20.21" />
                    <SPLIT distance="175" swimtime="00:02:37.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106765" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="106745" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="106772" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="106789" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="253" reactiontime="+79" swimtime="00:02:10.45" resultid="106892" heatid="110630" lane="3" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.97" />
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="75" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:01.45" />
                    <SPLIT distance="125" swimtime="00:01:16.55" />
                    <SPLIT distance="150" swimtime="00:01:32.86" />
                    <SPLIT distance="175" swimtime="00:01:50.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106778" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="106855" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="106843" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="106772" number="4" reactiontime="+80" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="373" reactiontime="+86" swimtime="00:01:54.70" resultid="106893" heatid="110631" lane="3" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.53" />
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                    <SPLIT distance="75" swimtime="00:00:40.64" />
                    <SPLIT distance="100" swimtime="00:00:54.93" />
                    <SPLIT distance="125" swimtime="00:01:08.10" />
                    <SPLIT distance="175" swimtime="00:01:37.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106882" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="106861" number="2" reactiontime="+11" />
                    <RELAYPOSITION athleteid="106796" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="106789" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="99441" points="169" reactiontime="+86" swimtime="00:02:43.60" resultid="106901" heatid="110836" lane="1" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.81" />
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                    <SPLIT distance="75" swimtime="00:01:01.21" />
                    <SPLIT distance="100" swimtime="00:01:25.71" />
                    <SPLIT distance="125" swimtime="00:01:42.69" />
                    <SPLIT distance="150" swimtime="00:02:04.86" />
                    <SPLIT distance="175" swimtime="00:02:23.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106823" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="106745" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="106805" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="106752" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="98846" points="189" reactiontime="+110" swimtime="00:02:23.77" resultid="110584" heatid="110630" lane="1" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.42" />
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="75" swimtime="00:00:49.89" />
                    <SPLIT distance="100" swimtime="00:01:06.77" />
                    <SPLIT distance="125" swimtime="00:01:25.64" />
                    <SPLIT distance="150" swimtime="00:01:35.57" />
                    <SPLIT distance="175" swimtime="00:02:04.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106752" number="1" reactiontime="+110" />
                    <RELAYPOSITION athleteid="106823" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="106745" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="106805" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="99441" points="221" reactiontime="+74" swimtime="00:02:29.63" resultid="106902" heatid="110836" lane="3" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.71" />
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="75" swimtime="00:00:58.25" />
                    <SPLIT distance="100" swimtime="00:01:18.94" />
                    <SPLIT distance="125" swimtime="00:01:35.01" />
                    <SPLIT distance="150" swimtime="00:01:53.97" />
                    <SPLIT distance="175" swimtime="00:02:10.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106778" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="106855" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="106851" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="106765" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="99441" reactiontime="+77" status="DSQ" swimtime="00:00:00.00" resultid="106903" heatid="110837" lane="4" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.14" />
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="75" swimtime="00:00:48.66" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="125" swimtime="00:01:21.58" />
                    <SPLIT distance="150" swimtime="00:01:37.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106882" number="1" reactiontime="+77" status="DSQ" />
                    <RELAYPOSITION athleteid="106784" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="106796" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="106861" number="4" reactiontime="-12" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="106905" name="Raduga">
          <CONTACT email="alkonter@gmail.com" name="Manevich" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Natalia" gender="F" lastname="Antsiferova" nation="RUS" athleteid="106941">
              <RESULTS>
                <RESULT eventid="98777" points="104" reactiontime="+111" swimtime="00:00:49.32" resultid="106942" heatid="110586" lane="4" entrytime="00:00:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="93" reactiontime="+95" swimtime="00:00:53.64" resultid="106943" heatid="110736" lane="2" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Mikhail" gender="M" lastname="Manevich" nation="RUS" athleteid="106936">
              <RESULTS>
                <RESULT eventid="98830" points="181" reactiontime="+82" swimtime="00:03:13.62" resultid="106937" heatid="110621" lane="2" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.07" />
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                    <SPLIT distance="75" swimtime="00:01:10.68" />
                    <SPLIT distance="100" swimtime="00:01:36.05" />
                    <SPLIT distance="125" swimtime="00:02:03.86" />
                    <SPLIT distance="150" swimtime="00:02:32.13" />
                    <SPLIT distance="175" swimtime="00:02:53.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="230" swimtime="00:01:13.27" resultid="106938" heatid="110681" lane="6" entrytime="00:01:14.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.81" />
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="75" swimtime="00:00:54.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="191" reactiontime="+95" swimtime="00:06:48.82" resultid="106939" heatid="110789" lane="8" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.05" />
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                    <SPLIT distance="75" swimtime="00:01:14.60" />
                    <SPLIT distance="100" swimtime="00:01:42.77" />
                    <SPLIT distance="125" swimtime="00:02:10.67" />
                    <SPLIT distance="150" swimtime="00:02:36.28" />
                    <SPLIT distance="175" swimtime="00:03:02.95" />
                    <SPLIT distance="200" swimtime="00:03:29.04" />
                    <SPLIT distance="225" swimtime="00:03:57.73" />
                    <SPLIT distance="250" swimtime="00:04:25.91" />
                    <SPLIT distance="275" swimtime="00:04:54.65" />
                    <SPLIT distance="300" swimtime="00:05:23.52" />
                    <SPLIT distance="325" swimtime="00:05:45.95" />
                    <SPLIT distance="350" swimtime="00:06:06.82" />
                    <SPLIT distance="375" swimtime="00:06:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="218" reactiontime="+113" swimtime="00:05:52.56" resultid="106940" heatid="110848" lane="1" entrytime="00:05:55.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.54" />
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="75" swimtime="00:00:59.33" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="125" swimtime="00:01:42.86" />
                    <SPLIT distance="150" swimtime="00:02:05.61" />
                    <SPLIT distance="175" swimtime="00:02:28.30" />
                    <SPLIT distance="200" swimtime="00:02:51.62" />
                    <SPLIT distance="225" swimtime="00:03:14.07" />
                    <SPLIT distance="250" swimtime="00:03:36.81" />
                    <SPLIT distance="275" swimtime="00:03:59.81" />
                    <SPLIT distance="300" swimtime="00:04:22.90" />
                    <SPLIT distance="325" swimtime="00:04:45.49" />
                    <SPLIT distance="350" swimtime="00:05:08.48" />
                    <SPLIT distance="375" swimtime="00:05:30.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Vladimir" gender="M" lastname="Efimets" nation="RUS" athleteid="106944">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="106945" heatid="110610" lane="3" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="107023" name="Redeco Wrocław">
          <CONTACT city="Wrocław" name="Wolny Dariusz" phone="603630870" state="DOL" street="Rogowska 52a" zip="55-440" />
          <ATHLETES>
            <ATHLETE birthdate="1969-12-31" firstname="Agata" gender="F" lastname="Szydło" nation="POL" athleteid="107038">
              <RESULTS>
                <RESULT eventid="98814" points="169" swimtime="00:03:40.33" resultid="107039" heatid="110615" lane="9" entrytime="00:03:49.37">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.52" />
                    <SPLIT distance="50" swimtime="00:00:49.84" />
                    <SPLIT distance="75" swimtime="00:01:19.27" />
                    <SPLIT distance="100" swimtime="00:01:49.51" />
                    <SPLIT distance="125" swimtime="00:02:18.41" />
                    <SPLIT distance="150" swimtime="00:02:48.50" />
                    <SPLIT distance="175" swimtime="00:03:14.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106254" points="178" reactiontime="+112" swimtime="00:27:14.12" resultid="107040" heatid="110640" lane="8" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.98" />
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="75" swimtime="00:01:15.45" />
                    <SPLIT distance="100" swimtime="00:01:41.57" />
                    <SPLIT distance="125" swimtime="00:02:08.11" />
                    <SPLIT distance="150" swimtime="00:02:34.24" />
                    <SPLIT distance="175" swimtime="00:03:01.15" />
                    <SPLIT distance="200" swimtime="00:03:28.33" />
                    <SPLIT distance="225" swimtime="00:03:55.46" />
                    <SPLIT distance="250" swimtime="00:04:22.58" />
                    <SPLIT distance="275" swimtime="00:04:49.82" />
                    <SPLIT distance="300" swimtime="00:05:17.53" />
                    <SPLIT distance="325" swimtime="00:05:44.64" />
                    <SPLIT distance="350" swimtime="00:06:12.29" />
                    <SPLIT distance="375" swimtime="00:06:40.00" />
                    <SPLIT distance="400" swimtime="00:07:07.89" />
                    <SPLIT distance="425" swimtime="00:07:34.95" />
                    <SPLIT distance="450" swimtime="00:08:02.40" />
                    <SPLIT distance="475" swimtime="00:08:30.05" />
                    <SPLIT distance="500" swimtime="00:08:57.50" />
                    <SPLIT distance="525" swimtime="00:09:24.99" />
                    <SPLIT distance="550" swimtime="00:09:52.48" />
                    <SPLIT distance="575" swimtime="00:10:20.01" />
                    <SPLIT distance="600" swimtime="00:10:47.40" />
                    <SPLIT distance="625" swimtime="00:11:15.02" />
                    <SPLIT distance="650" swimtime="00:11:42.63" />
                    <SPLIT distance="675" swimtime="00:12:10.22" />
                    <SPLIT distance="700" swimtime="00:12:37.83" />
                    <SPLIT distance="725" swimtime="00:13:05.76" />
                    <SPLIT distance="750" swimtime="00:13:33.47" />
                    <SPLIT distance="775" swimtime="00:14:01.10" />
                    <SPLIT distance="800" swimtime="00:14:28.27" />
                    <SPLIT distance="825" swimtime="00:14:56.41" />
                    <SPLIT distance="850" swimtime="00:15:23.47" />
                    <SPLIT distance="875" swimtime="00:15:51.10" />
                    <SPLIT distance="900" swimtime="00:16:19.09" />
                    <SPLIT distance="925" swimtime="00:16:46.68" />
                    <SPLIT distance="950" swimtime="00:17:14.15" />
                    <SPLIT distance="975" swimtime="00:17:42.01" />
                    <SPLIT distance="1000" swimtime="00:18:09.91" />
                    <SPLIT distance="1025" swimtime="00:18:37.70" />
                    <SPLIT distance="1050" swimtime="00:19:04.93" />
                    <SPLIT distance="1075" swimtime="00:19:32.69" />
                    <SPLIT distance="1100" swimtime="00:19:59.94" />
                    <SPLIT distance="1125" swimtime="00:20:27.83" />
                    <SPLIT distance="1150" swimtime="00:20:55.38" />
                    <SPLIT distance="1175" swimtime="00:21:22.87" />
                    <SPLIT distance="1200" swimtime="00:21:50.11" />
                    <SPLIT distance="1225" swimtime="00:22:17.28" />
                    <SPLIT distance="1250" swimtime="00:22:44.73" />
                    <SPLIT distance="1275" swimtime="00:23:12.19" />
                    <SPLIT distance="1300" swimtime="00:23:39.49" />
                    <SPLIT distance="1325" swimtime="00:24:06.87" />
                    <SPLIT distance="1350" swimtime="00:24:34.14" />
                    <SPLIT distance="1375" swimtime="00:25:01.68" />
                    <SPLIT distance="1400" swimtime="00:25:28.75" />
                    <SPLIT distance="1425" swimtime="00:25:56.06" />
                    <SPLIT distance="1450" swimtime="00:26:22.36" />
                    <SPLIT distance="1475" swimtime="00:26:48.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="207" reactiontime="+109" swimtime="00:03:47.15" resultid="107041" heatid="110662" lane="2" entrytime="00:03:44.83">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.39" />
                    <SPLIT distance="50" swimtime="00:00:53.17" />
                    <SPLIT distance="75" swimtime="00:01:22.14" />
                    <SPLIT distance="100" swimtime="00:01:50.72" />
                    <SPLIT distance="125" swimtime="00:02:20.05" />
                    <SPLIT distance="150" swimtime="00:02:49.26" />
                    <SPLIT distance="175" swimtime="00:03:18.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="172" reactiontime="+103" swimtime="00:01:41.81" resultid="107042" heatid="110691" lane="7" entrytime="00:01:42.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.20" />
                    <SPLIT distance="50" swimtime="00:00:50.78" />
                    <SPLIT distance="75" swimtime="00:01:18.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="195" reactiontime="+94" swimtime="00:01:47.36" resultid="107043" heatid="110722" lane="8" entrytime="00:01:46.64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.58" />
                    <SPLIT distance="50" swimtime="00:00:51.75" />
                    <SPLIT distance="75" swimtime="00:01:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="170" swimtime="00:07:47.88" resultid="107044" heatid="110785" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.33" />
                    <SPLIT distance="50" swimtime="00:00:54.86" />
                    <SPLIT distance="75" swimtime="00:01:25.07" />
                    <SPLIT distance="100" swimtime="00:01:56.65" />
                    <SPLIT distance="125" swimtime="00:02:27.10" />
                    <SPLIT distance="150" swimtime="00:02:58.46" />
                    <SPLIT distance="175" swimtime="00:03:28.78" />
                    <SPLIT distance="200" swimtime="00:04:01.80" />
                    <SPLIT distance="225" swimtime="00:04:31.02" />
                    <SPLIT distance="250" swimtime="00:05:01.59" />
                    <SPLIT distance="275" swimtime="00:05:31.69" />
                    <SPLIT distance="300" swimtime="00:06:02.05" />
                    <SPLIT distance="325" swimtime="00:06:28.42" />
                    <SPLIT distance="350" swimtime="00:06:55.65" />
                    <SPLIT distance="375" swimtime="00:07:22.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="194" reactiontime="+98" swimtime="00:00:49.71" resultid="107045" heatid="110819" lane="1" entrytime="00:00:49.96">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="175" reactiontime="+97" swimtime="00:06:59.03" resultid="107046" heatid="110842" lane="4" entrytime="00:06:49.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.16" />
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                    <SPLIT distance="75" swimtime="00:01:13.42" />
                    <SPLIT distance="100" swimtime="00:01:39.50" />
                    <SPLIT distance="125" swimtime="00:02:05.81" />
                    <SPLIT distance="150" swimtime="00:02:32.40" />
                    <SPLIT distance="175" swimtime="00:02:59.12" />
                    <SPLIT distance="200" swimtime="00:03:26.25" />
                    <SPLIT distance="225" swimtime="00:04:47.85" />
                    <SPLIT distance="250" swimtime="00:04:20.34" />
                    <SPLIT distance="275" swimtime="00:05:42.72" />
                    <SPLIT distance="300" swimtime="00:05:15.59" />
                    <SPLIT distance="350" swimtime="00:06:09.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-13" firstname="Małgorzata" gender="F" lastname="Bołtuć" nation="POL" athleteid="107030">
              <RESULTS>
                <RESULT eventid="98814" points="219" reactiontime="+112" swimtime="00:03:21.89" resultid="107031" heatid="110615" lane="3" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.66" />
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                    <SPLIT distance="75" swimtime="00:01:09.13" />
                    <SPLIT distance="100" swimtime="00:01:35.30" />
                    <SPLIT distance="125" swimtime="00:02:05.03" />
                    <SPLIT distance="150" swimtime="00:02:34.94" />
                    <SPLIT distance="175" swimtime="00:02:58.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106254" points="222" swimtime="00:25:17.64" resultid="107032" heatid="110640" lane="1" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.32" />
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                    <SPLIT distance="75" swimtime="00:01:08.11" />
                    <SPLIT distance="100" swimtime="00:01:31.39" />
                    <SPLIT distance="125" swimtime="00:01:56.60" />
                    <SPLIT distance="150" swimtime="00:02:21.05" />
                    <SPLIT distance="175" swimtime="00:02:45.73" />
                    <SPLIT distance="200" swimtime="00:03:11.42" />
                    <SPLIT distance="225" swimtime="00:03:36.04" />
                    <SPLIT distance="250" swimtime="00:04:01.44" />
                    <SPLIT distance="275" swimtime="00:04:26.56" />
                    <SPLIT distance="300" swimtime="00:04:52.76" />
                    <SPLIT distance="325" swimtime="00:05:19.26" />
                    <SPLIT distance="350" swimtime="00:05:44.70" />
                    <SPLIT distance="375" swimtime="00:06:10.05" />
                    <SPLIT distance="400" swimtime="00:06:35.84" />
                    <SPLIT distance="425" swimtime="00:07:01.32" />
                    <SPLIT distance="450" swimtime="00:07:27.11" />
                    <SPLIT distance="475" swimtime="00:07:52.83" />
                    <SPLIT distance="500" swimtime="00:08:18.44" />
                    <SPLIT distance="525" swimtime="00:08:43.16" />
                    <SPLIT distance="550" swimtime="00:09:08.42" />
                    <SPLIT distance="575" swimtime="00:09:33.76" />
                    <SPLIT distance="600" swimtime="00:09:59.41" />
                    <SPLIT distance="625" swimtime="00:10:25.32" />
                    <SPLIT distance="650" swimtime="00:10:51.09" />
                    <SPLIT distance="675" swimtime="00:11:16.62" />
                    <SPLIT distance="700" swimtime="00:11:42.03" />
                    <SPLIT distance="725" swimtime="00:12:07.52" />
                    <SPLIT distance="750" swimtime="00:12:33.23" />
                    <SPLIT distance="775" swimtime="00:12:58.84" />
                    <SPLIT distance="800" swimtime="00:13:24.44" />
                    <SPLIT distance="825" swimtime="00:13:50.59" />
                    <SPLIT distance="850" swimtime="00:14:15.63" />
                    <SPLIT distance="875" swimtime="00:14:42.27" />
                    <SPLIT distance="900" swimtime="00:15:07.18" />
                    <SPLIT distance="925" swimtime="00:15:33.79" />
                    <SPLIT distance="950" swimtime="00:15:59.57" />
                    <SPLIT distance="975" swimtime="00:16:25.37" />
                    <SPLIT distance="1000" swimtime="00:16:51.40" />
                    <SPLIT distance="1025" swimtime="00:17:16.78" />
                    <SPLIT distance="1050" swimtime="00:17:43.05" />
                    <SPLIT distance="1075" swimtime="00:18:09.29" />
                    <SPLIT distance="1100" swimtime="00:18:34.45" />
                    <SPLIT distance="1125" swimtime="00:19:00.36" />
                    <SPLIT distance="1150" swimtime="00:19:26.00" />
                    <SPLIT distance="1175" swimtime="00:19:52.53" />
                    <SPLIT distance="1200" swimtime="00:20:16.70" />
                    <SPLIT distance="1225" swimtime="00:20:42.20" />
                    <SPLIT distance="1250" swimtime="00:21:07.88" />
                    <SPLIT distance="1275" swimtime="00:21:33.86" />
                    <SPLIT distance="1300" swimtime="00:21:58.75" />
                    <SPLIT distance="1325" swimtime="00:22:24.81" />
                    <SPLIT distance="1350" swimtime="00:22:49.59" />
                    <SPLIT distance="1375" swimtime="00:23:14.53" />
                    <SPLIT distance="1400" swimtime="00:23:38.91" />
                    <SPLIT distance="1425" swimtime="00:24:04.00" />
                    <SPLIT distance="1450" swimtime="00:24:29.02" />
                    <SPLIT distance="1475" swimtime="00:24:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="205" reactiontime="+117" swimtime="00:01:35.99" resultid="107033" heatid="110691" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.55" />
                    <SPLIT distance="50" swimtime="00:00:45.72" />
                    <SPLIT distance="75" swimtime="00:01:14.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="192" swimtime="00:00:42.26" resultid="107034" heatid="110737" lane="6" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="216" swimtime="00:07:12.34" resultid="107035" heatid="110786" lane="8" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.73" />
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                    <SPLIT distance="75" swimtime="00:01:16.12" />
                    <SPLIT distance="100" swimtime="00:01:46.23" />
                    <SPLIT distance="125" swimtime="00:02:13.77" />
                    <SPLIT distance="150" swimtime="00:02:40.85" />
                    <SPLIT distance="175" swimtime="00:03:08.57" />
                    <SPLIT distance="200" swimtime="00:03:36.92" />
                    <SPLIT distance="225" swimtime="00:04:06.43" />
                    <SPLIT distance="250" swimtime="00:04:36.68" />
                    <SPLIT distance="275" swimtime="00:05:07.27" />
                    <SPLIT distance="300" swimtime="00:05:38.78" />
                    <SPLIT distance="325" swimtime="00:06:02.18" />
                    <SPLIT distance="350" swimtime="00:06:26.46" />
                    <SPLIT distance="375" swimtime="00:06:49.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="172" reactiontime="+115" swimtime="00:01:38.10" resultid="107036" heatid="110794" lane="1" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.19" />
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                    <SPLIT distance="75" swimtime="00:01:11.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="213" reactiontime="+102" swimtime="00:03:19.37" resultid="107037" heatid="110807" lane="7" entrytime="00:03:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.00" />
                    <SPLIT distance="50" swimtime="00:00:48.57" />
                    <SPLIT distance="75" swimtime="00:01:14.08" />
                    <SPLIT distance="100" swimtime="00:01:39.63" />
                    <SPLIT distance="125" swimtime="00:02:05.07" />
                    <SPLIT distance="150" swimtime="00:02:30.44" />
                    <SPLIT distance="175" swimtime="00:02:55.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-03-21" firstname="Dariusz" gender="M" lastname="Wolny" nation="POL" athleteid="107024">
              <RESULTS>
                <RESULT eventid="98830" points="391" reactiontime="+86" swimtime="00:02:29.84" resultid="107025" heatid="110626" lane="3" entrytime="00:02:31.31">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.65" />
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="75" swimtime="00:00:50.45" />
                    <SPLIT distance="100" swimtime="00:01:08.76" />
                    <SPLIT distance="125" swimtime="00:01:31.10" />
                    <SPLIT distance="150" swimtime="00:01:53.98" />
                    <SPLIT distance="175" swimtime="00:02:12.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="349" reactiontime="+71" swimtime="00:00:31.53" resultid="107026" heatid="110659" lane="8" entrytime="00:00:31.31">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="402" reactiontime="+87" swimtime="00:01:08.62" resultid="107027" heatid="110704" lane="1" entrytime="00:01:08.08">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.32" />
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="75" swimtime="00:00:52.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="365" reactiontime="+77" swimtime="00:01:08.41" resultid="107028" heatid="110762" lane="4" entrytime="00:01:07.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.44" />
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="75" swimtime="00:00:51.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="373" reactiontime="+73" swimtime="00:02:26.72" resultid="107029" heatid="110815" lane="5" entrytime="00:02:29.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.76" />
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="75" swimtime="00:00:52.68" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="125" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:01:49.01" />
                    <SPLIT distance="175" swimtime="00:02:08.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RMKS RYBNI" nation="POL" region="SLA" clubid="108264" name="RMKS Rybnik">
          <CONTACT city="Rybnik" email="aniaduda0511@tlen.pl" name="Duda Anna" phone="792666159" state="SLA" street="Powstańców sl 40/42" zip="44-200" />
          <ATHLETES>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="108265">
              <RESULTS>
                <RESULT eventid="98777" points="573" reactiontime="+79" swimtime="00:00:27.97" resultid="108266" heatid="110593" lane="8" entrytime="00:00:28.03">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="441" reactiontime="+87" swimtime="00:02:40.06" resultid="108267" heatid="110618" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.03" />
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="75" swimtime="00:00:54.70" />
                    <SPLIT distance="100" swimtime="00:01:15.54" />
                    <SPLIT distance="125" swimtime="00:01:39.33" />
                    <SPLIT distance="150" swimtime="00:02:03.86" />
                    <SPLIT distance="175" swimtime="00:02:22.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="526" reactiontime="+89" swimtime="00:01:03.04" resultid="108268" heatid="110676" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.21" />
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                    <SPLIT distance="75" swimtime="00:00:46.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="294" reactiontime="+91" swimtime="00:02:59.84" resultid="108269" heatid="110708" lane="5" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.68" />
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="75" swimtime="00:00:59.54" />
                    <SPLIT distance="100" swimtime="00:01:24.47" />
                    <SPLIT distance="125" swimtime="00:01:49.44" />
                    <SPLIT distance="150" swimtime="00:02:14.09" />
                    <SPLIT distance="175" swimtime="00:02:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="549" reactiontime="+77" swimtime="00:00:29.76" resultid="108270" heatid="110740" lane="5" entrytime="00:00:29.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="399" reactiontime="+93" swimtime="00:05:52.24" resultid="108271" heatid="110787" lane="5" entrytime="00:05:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.20" />
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="75" swimtime="00:00:57.04" />
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="125" swimtime="00:01:43.31" />
                    <SPLIT distance="150" swimtime="00:02:06.82" />
                    <SPLIT distance="175" swimtime="00:02:30.60" />
                    <SPLIT distance="200" swimtime="00:02:54.36" />
                    <SPLIT distance="225" swimtime="00:03:19.23" />
                    <SPLIT distance="250" swimtime="00:03:44.74" />
                    <SPLIT distance="275" swimtime="00:04:09.92" />
                    <SPLIT distance="300" swimtime="00:04:36.38" />
                    <SPLIT distance="325" swimtime="00:04:57.10" />
                    <SPLIT distance="350" swimtime="00:05:16.38" />
                    <SPLIT distance="375" swimtime="00:05:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="487" reactiontime="+69" swimtime="00:01:09.39" resultid="108272" heatid="110796" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.41" />
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="75" swimtime="00:00:50.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="428" swimtime="00:00:38.20" resultid="108273" heatid="110822" lane="0" entrytime="00:00:39.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="108152" name="Rydułtowska Akademia Aktywnego Seniora 60+" shortname="Rydułtowska Akademia Aktywnego">
          <CONTACT email="otelom.080966@interia.pl" name="OTLIK MARIAN" />
          <ATHLETES>
            <ATHLETE birthdate="1966-09-08" firstname="Marian" gender="M" lastname="Otlik" nation="POL" athleteid="108179">
              <RESULTS>
                <RESULT comment="O4" eventid="98798" status="DSQ" swimtime="00:00:00.00" resultid="108180" heatid="110604" lane="9" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="204" reactiontime="+66" swimtime="00:03:05.97" resultid="108181" heatid="110621" lane="6" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.65" />
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="75" swimtime="00:01:02.09" />
                    <SPLIT distance="100" swimtime="00:01:25.67" />
                    <SPLIT distance="125" swimtime="00:01:53.66" />
                    <SPLIT distance="150" swimtime="00:02:21.45" />
                    <SPLIT distance="175" swimtime="00:02:44.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="269" reactiontime="+57" swimtime="00:01:09.58" resultid="108182" heatid="110682" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.66" />
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="75" swimtime="00:00:51.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="241" swimtime="00:01:21.30" resultid="108183" heatid="110698" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.74" />
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="75" swimtime="00:01:02.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="259" reactiontime="+78" swimtime="00:00:34.16" resultid="108184" heatid="110744" lane="2" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="108185" heatid="110789" lane="9" entrytime="00:07:10.00" />
                <RESULT eventid="99361" points="202" reactiontime="+72" swimtime="00:01:22.55" resultid="108186" heatid="110800" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.14" />
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="75" swimtime="00:00:59.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="108187" heatid="110848" lane="9" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="108171">
              <RESULTS>
                <RESULT eventid="98830" points="67" reactiontime="+96" swimtime="00:04:29.37" resultid="108172" heatid="110619" lane="4" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.63" />
                    <SPLIT distance="50" swimtime="00:01:02.53" />
                    <SPLIT distance="75" swimtime="00:01:35.07" />
                    <SPLIT distance="100" swimtime="00:02:11.07" />
                    <SPLIT distance="125" swimtime="00:02:48.89" />
                    <SPLIT distance="150" swimtime="00:03:25.57" />
                    <SPLIT distance="175" swimtime="00:03:57.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="52" reactiontime="+85" swimtime="00:00:59.36" resultid="108173" heatid="110652" lane="2" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="43" reactiontime="+110" swimtime="00:05:09.64" resultid="108174" heatid="110710" lane="1" entrytime="00:04:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.65" />
                    <SPLIT distance="50" swimtime="00:01:07.56" />
                    <SPLIT distance="75" swimtime="00:01:46.09" />
                    <SPLIT distance="100" swimtime="00:02:24.86" />
                    <SPLIT distance="125" swimtime="00:03:03.67" />
                    <SPLIT distance="150" swimtime="00:03:44.58" />
                    <SPLIT distance="175" swimtime="00:04:26.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="49" swimtime="00:00:59.43" resultid="108175" heatid="110742" lane="0" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="55" reactiontime="+115" swimtime="00:10:18.09" resultid="108176" heatid="110788" lane="1" entrytime="00:09:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.05" />
                    <SPLIT distance="50" swimtime="00:01:10.82" />
                    <SPLIT distance="75" swimtime="00:01:51.44" />
                    <SPLIT distance="100" swimtime="00:02:35.57" />
                    <SPLIT distance="125" swimtime="00:03:14.80" />
                    <SPLIT distance="150" swimtime="00:03:54.07" />
                    <SPLIT distance="175" swimtime="00:04:33.59" />
                    <SPLIT distance="200" swimtime="00:05:13.49" />
                    <SPLIT distance="225" swimtime="00:05:55.19" />
                    <SPLIT distance="250" swimtime="00:06:34.87" />
                    <SPLIT distance="275" swimtime="00:07:14.63" />
                    <SPLIT distance="300" swimtime="00:07:55.85" />
                    <SPLIT distance="325" swimtime="00:08:30.47" />
                    <SPLIT distance="350" swimtime="00:09:06.84" />
                    <SPLIT distance="375" swimtime="00:09:43.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="39" reactiontime="+115" swimtime="00:02:22.16" resultid="108177" heatid="110798" lane="1" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.25" />
                    <SPLIT distance="50" swimtime="00:01:04.11" />
                    <SPLIT distance="75" swimtime="00:01:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="48" reactiontime="+97" swimtime="00:04:48.84" resultid="108178" heatid="110811" lane="0" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.61" />
                    <SPLIT distance="50" swimtime="00:01:09.41" />
                    <SPLIT distance="75" swimtime="00:01:47.97" />
                    <SPLIT distance="100" swimtime="00:02:24.89" />
                    <SPLIT distance="125" swimtime="00:03:02.37" />
                    <SPLIT distance="150" swimtime="00:03:39.05" />
                    <SPLIT distance="175" swimtime="00:04:15.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-07" firstname="Leon" gender="M" lastname="Irczyk" nation="POL" athleteid="108162">
              <RESULTS>
                <RESULT eventid="98830" points="95" reactiontime="+126" swimtime="00:04:00.12" resultid="108163" heatid="110620" lane="7" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.27" />
                    <SPLIT distance="50" swimtime="00:00:55.05" />
                    <SPLIT distance="75" swimtime="00:01:33.90" />
                    <SPLIT distance="100" swimtime="00:02:09.58" />
                    <SPLIT distance="125" swimtime="00:02:37.84" />
                    <SPLIT distance="150" swimtime="00:03:07.19" />
                    <SPLIT distance="175" swimtime="00:03:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="119" reactiontime="+135" swimtime="00:28:40.68" resultid="108164" heatid="110643" lane="0" entrytime="00:32:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.37" />
                    <SPLIT distance="50" swimtime="00:00:50.49" />
                    <SPLIT distance="75" swimtime="00:01:18.92" />
                    <SPLIT distance="100" swimtime="00:01:47.66" />
                    <SPLIT distance="125" swimtime="00:02:16.43" />
                    <SPLIT distance="150" swimtime="00:02:45.76" />
                    <SPLIT distance="175" swimtime="00:03:14.25" />
                    <SPLIT distance="200" swimtime="00:03:42.60" />
                    <SPLIT distance="225" swimtime="00:04:10.67" />
                    <SPLIT distance="250" swimtime="00:04:39.22" />
                    <SPLIT distance="275" swimtime="00:05:07.66" />
                    <SPLIT distance="300" swimtime="00:05:36.26" />
                    <SPLIT distance="325" swimtime="00:06:04.71" />
                    <SPLIT distance="350" swimtime="00:06:33.64" />
                    <SPLIT distance="375" swimtime="00:07:02.15" />
                    <SPLIT distance="400" swimtime="00:07:31.20" />
                    <SPLIT distance="425" swimtime="00:08:00.00" />
                    <SPLIT distance="450" swimtime="00:08:29.33" />
                    <SPLIT distance="475" swimtime="00:08:58.30" />
                    <SPLIT distance="500" swimtime="00:09:27.12" />
                    <SPLIT distance="525" swimtime="00:09:55.90" />
                    <SPLIT distance="550" swimtime="00:10:24.72" />
                    <SPLIT distance="575" swimtime="00:10:53.73" />
                    <SPLIT distance="600" swimtime="00:11:22.65" />
                    <SPLIT distance="625" swimtime="00:11:50.82" />
                    <SPLIT distance="650" swimtime="00:12:19.98" />
                    <SPLIT distance="675" swimtime="00:12:48.37" />
                    <SPLIT distance="700" swimtime="00:13:17.75" />
                    <SPLIT distance="725" swimtime="00:13:45.51" />
                    <SPLIT distance="750" swimtime="00:14:15.32" />
                    <SPLIT distance="775" swimtime="00:14:44.19" />
                    <SPLIT distance="800" swimtime="00:15:13.81" />
                    <SPLIT distance="825" swimtime="00:15:42.09" />
                    <SPLIT distance="850" swimtime="00:16:11.63" />
                    <SPLIT distance="875" swimtime="00:16:39.93" />
                    <SPLIT distance="900" swimtime="00:17:09.75" />
                    <SPLIT distance="925" swimtime="00:17:38.10" />
                    <SPLIT distance="950" swimtime="00:18:07.71" />
                    <SPLIT distance="975" swimtime="00:18:36.11" />
                    <SPLIT distance="1000" swimtime="00:19:05.47" />
                    <SPLIT distance="1025" swimtime="00:19:33.41" />
                    <SPLIT distance="1050" swimtime="00:20:02.73" />
                    <SPLIT distance="1075" swimtime="00:20:31.44" />
                    <SPLIT distance="1100" swimtime="00:21:00.90" />
                    <SPLIT distance="1125" swimtime="00:21:29.29" />
                    <SPLIT distance="1150" swimtime="00:21:58.98" />
                    <SPLIT distance="1175" swimtime="00:22:27.55" />
                    <SPLIT distance="1200" swimtime="00:22:57.60" />
                    <SPLIT distance="1225" swimtime="00:23:25.68" />
                    <SPLIT distance="1250" swimtime="00:23:54.93" />
                    <SPLIT distance="1275" swimtime="00:24:23.83" />
                    <SPLIT distance="1300" swimtime="00:24:52.98" />
                    <SPLIT distance="1325" swimtime="00:25:22.63" />
                    <SPLIT distance="1350" swimtime="00:25:51.32" />
                    <SPLIT distance="1375" swimtime="00:26:20.99" />
                    <SPLIT distance="1400" swimtime="00:26:50.34" />
                    <SPLIT distance="1425" swimtime="00:27:19.39" />
                    <SPLIT distance="1450" swimtime="00:27:47.55" />
                    <SPLIT distance="1475" swimtime="00:28:16.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="142" reactiontime="+113" swimtime="00:03:50.87" resultid="108165" heatid="110666" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.66" />
                    <SPLIT distance="50" swimtime="00:00:52.45" />
                    <SPLIT distance="75" swimtime="00:01:20.95" />
                    <SPLIT distance="100" swimtime="00:01:50.39" />
                    <SPLIT distance="125" swimtime="00:02:20.55" />
                    <SPLIT distance="150" swimtime="00:02:50.57" />
                    <SPLIT distance="175" swimtime="00:03:21.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="79" reactiontime="+129" swimtime="00:01:57.60" resultid="108166" heatid="110697" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.79" />
                    <SPLIT distance="50" swimtime="00:01:03.70" />
                    <SPLIT distance="75" swimtime="00:01:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="132" reactiontime="+115" swimtime="00:01:49.14" resultid="108167" heatid="110728" lane="3" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.02" />
                    <SPLIT distance="50" swimtime="00:00:51.23" />
                    <SPLIT distance="75" swimtime="00:01:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="98" swimtime="00:08:30.52" resultid="108168" heatid="110788" lane="6" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.96" />
                    <SPLIT distance="50" swimtime="00:00:56.27" />
                    <SPLIT distance="75" swimtime="00:01:28.77" />
                    <SPLIT distance="100" swimtime="00:02:02.55" />
                    <SPLIT distance="125" swimtime="00:02:43.88" />
                    <SPLIT distance="150" swimtime="00:03:21.32" />
                    <SPLIT distance="175" swimtime="00:03:58.01" />
                    <SPLIT distance="200" swimtime="00:04:36.25" />
                    <SPLIT distance="225" swimtime="00:05:06.23" />
                    <SPLIT distance="250" swimtime="00:05:37.40" />
                    <SPLIT distance="275" swimtime="00:06:08.48" />
                    <SPLIT distance="300" swimtime="00:06:38.88" />
                    <SPLIT distance="325" swimtime="00:07:08.44" />
                    <SPLIT distance="350" swimtime="00:07:37.62" />
                    <SPLIT distance="375" swimtime="00:08:05.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="65" reactiontime="+130" swimtime="00:02:00.12" resultid="108169" heatid="110798" lane="4" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.43" />
                    <SPLIT distance="50" swimtime="00:00:56.37" />
                    <SPLIT distance="75" swimtime="00:01:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="108170" heatid="110851" lane="6" entrytime="00:07:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="108153">
              <RESULTS>
                <RESULT eventid="98830" points="173" reactiontime="+92" swimtime="00:03:16.44" resultid="108154" heatid="110621" lane="7" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.55" />
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="75" swimtime="00:01:06.49" />
                    <SPLIT distance="100" swimtime="00:01:31.64" />
                    <SPLIT distance="125" swimtime="00:02:02.70" />
                    <SPLIT distance="150" swimtime="00:02:32.97" />
                    <SPLIT distance="175" swimtime="00:02:55.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="186" reactiontime="+96" swimtime="00:24:43.08" resultid="108155" heatid="110643" lane="3" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.81" />
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="75" swimtime="00:01:06.38" />
                    <SPLIT distance="100" swimtime="00:01:29.94" />
                    <SPLIT distance="125" swimtime="00:01:53.94" />
                    <SPLIT distance="150" swimtime="00:02:18.13" />
                    <SPLIT distance="175" swimtime="00:02:42.65" />
                    <SPLIT distance="200" swimtime="00:03:06.99" />
                    <SPLIT distance="225" swimtime="00:03:31.67" />
                    <SPLIT distance="250" swimtime="00:03:56.38" />
                    <SPLIT distance="275" swimtime="00:04:21.46" />
                    <SPLIT distance="300" swimtime="00:04:46.34" />
                    <SPLIT distance="325" swimtime="00:05:10.83" />
                    <SPLIT distance="350" swimtime="00:05:35.73" />
                    <SPLIT distance="375" swimtime="00:06:00.81" />
                    <SPLIT distance="400" swimtime="00:06:25.77" />
                    <SPLIT distance="425" swimtime="00:06:50.76" />
                    <SPLIT distance="450" swimtime="00:07:15.71" />
                    <SPLIT distance="475" swimtime="00:07:40.44" />
                    <SPLIT distance="500" swimtime="00:08:05.59" />
                    <SPLIT distance="525" swimtime="00:08:30.47" />
                    <SPLIT distance="550" swimtime="00:08:55.28" />
                    <SPLIT distance="575" swimtime="00:09:20.13" />
                    <SPLIT distance="600" swimtime="00:09:45.11" />
                    <SPLIT distance="625" swimtime="00:10:09.96" />
                    <SPLIT distance="650" swimtime="00:10:35.12" />
                    <SPLIT distance="675" swimtime="00:11:00.09" />
                    <SPLIT distance="700" swimtime="00:11:25.48" />
                    <SPLIT distance="725" swimtime="00:11:50.21" />
                    <SPLIT distance="750" swimtime="00:12:15.21" />
                    <SPLIT distance="775" swimtime="00:12:39.99" />
                    <SPLIT distance="800" swimtime="00:13:05.24" />
                    <SPLIT distance="825" swimtime="00:13:30.35" />
                    <SPLIT distance="850" swimtime="00:13:55.47" />
                    <SPLIT distance="875" swimtime="00:14:20.45" />
                    <SPLIT distance="900" swimtime="00:14:45.59" />
                    <SPLIT distance="925" swimtime="00:15:10.79" />
                    <SPLIT distance="950" swimtime="00:15:35.88" />
                    <SPLIT distance="975" swimtime="00:16:00.80" />
                    <SPLIT distance="1000" swimtime="00:16:25.70" />
                    <SPLIT distance="1025" swimtime="00:16:50.41" />
                    <SPLIT distance="1050" swimtime="00:17:15.35" />
                    <SPLIT distance="1075" swimtime="00:17:40.29" />
                    <SPLIT distance="1100" swimtime="00:18:05.46" />
                    <SPLIT distance="1125" swimtime="00:18:30.27" />
                    <SPLIT distance="1150" swimtime="00:18:55.42" />
                    <SPLIT distance="1175" swimtime="00:19:20.34" />
                    <SPLIT distance="1200" swimtime="00:19:45.41" />
                    <SPLIT distance="1225" swimtime="00:20:10.44" />
                    <SPLIT distance="1250" swimtime="00:20:35.37" />
                    <SPLIT distance="1275" swimtime="00:21:00.18" />
                    <SPLIT distance="1300" swimtime="00:21:25.06" />
                    <SPLIT distance="1325" swimtime="00:21:49.96" />
                    <SPLIT distance="1350" swimtime="00:22:15.05" />
                    <SPLIT distance="1375" swimtime="00:22:40.20" />
                    <SPLIT distance="1400" swimtime="00:23:05.01" />
                    <SPLIT distance="1425" swimtime="00:23:30.03" />
                    <SPLIT distance="1450" swimtime="00:23:54.74" />
                    <SPLIT distance="1475" swimtime="00:24:19.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="156" reactiontime="+86" swimtime="00:00:41.26" resultid="108156" heatid="110653" lane="5" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="106" swimtime="00:03:49.07" resultid="108157" heatid="110711" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.57" />
                    <SPLIT distance="50" swimtime="00:00:47.56" />
                    <SPLIT distance="75" swimtime="00:01:16.29" />
                    <SPLIT distance="100" swimtime="00:01:46.53" />
                    <SPLIT distance="125" swimtime="00:02:16.58" />
                    <SPLIT distance="150" swimtime="00:02:48.14" />
                    <SPLIT distance="175" swimtime="00:03:19.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="145" reactiontime="+71" swimtime="00:01:33.05" resultid="108158" heatid="110759" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.13" />
                    <SPLIT distance="50" swimtime="00:00:45.63" />
                    <SPLIT distance="75" swimtime="00:01:09.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="153" reactiontime="+94" swimtime="00:07:19.95" resultid="108159" heatid="110788" lane="5" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.60" />
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                    <SPLIT distance="75" swimtime="00:01:15.18" />
                    <SPLIT distance="100" swimtime="00:01:45.55" />
                    <SPLIT distance="125" swimtime="00:02:13.89" />
                    <SPLIT distance="150" swimtime="00:03:39.30" />
                    <SPLIT distance="175" swimtime="00:03:11.08" />
                    <SPLIT distance="200" swimtime="00:04:43.09" />
                    <SPLIT distance="225" swimtime="00:04:11.39" />
                    <SPLIT distance="250" swimtime="00:05:43.56" />
                    <SPLIT distance="275" swimtime="00:05:12.88" />
                    <SPLIT distance="325" swimtime="00:06:07.64" />
                    <SPLIT distance="350" swimtime="00:06:31.88" />
                    <SPLIT distance="375" swimtime="00:06:56.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="156" swimtime="00:01:29.81" resultid="108160" heatid="110800" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.77" />
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="75" swimtime="00:01:05.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="142" reactiontime="+89" swimtime="00:03:22.06" resultid="108161" heatid="110812" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.24" />
                    <SPLIT distance="50" swimtime="00:00:46.32" />
                    <SPLIT distance="75" swimtime="00:01:12.10" />
                    <SPLIT distance="100" swimtime="00:01:38.33" />
                    <SPLIT distance="125" swimtime="00:02:04.69" />
                    <SPLIT distance="150" swimtime="00:02:31.23" />
                    <SPLIT distance="175" swimtime="00:02:57.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="110218" name="Sikret Gliwice">
          <CONTACT city="Gliwice" email="joannaeco@wp.pl" internet="www.sikret-plywanie.pl" name="Joanna Zagała" street="Jagielońska 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="110228">
              <RESULTS>
                <RESULT eventid="98777" points="190" reactiontime="+87" swimtime="00:00:40.39" resultid="110229" heatid="110587" lane="6" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="160" reactiontime="+81" swimtime="00:04:07.55" resultid="110230" heatid="110661" lane="5" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.78" />
                    <SPLIT distance="50" swimtime="00:00:53.59" />
                    <SPLIT distance="75" swimtime="00:01:23.82" />
                    <SPLIT distance="100" swimtime="00:01:55.59" />
                    <SPLIT distance="125" swimtime="00:02:28.58" />
                    <SPLIT distance="150" swimtime="00:03:01.81" />
                    <SPLIT distance="175" swimtime="00:03:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="69" reactiontime="+98" swimtime="00:04:50.38" resultid="110231" heatid="110707" lane="3" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.25" />
                    <SPLIT distance="50" swimtime="00:01:05.55" />
                    <SPLIT distance="75" swimtime="00:01:40.70" />
                    <SPLIT distance="100" swimtime="00:02:20.21" />
                    <SPLIT distance="125" swimtime="00:02:57.69" />
                    <SPLIT distance="150" swimtime="00:03:37.76" />
                    <SPLIT distance="175" swimtime="00:04:16.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="179" reactiontime="+97" swimtime="00:01:50.55" resultid="110232" heatid="110721" lane="4" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.54" />
                    <SPLIT distance="50" swimtime="00:00:52.49" />
                    <SPLIT distance="75" swimtime="00:01:21.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="107" reactiontime="+101" swimtime="00:09:06.17" resultid="110233" heatid="110785" lane="5" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.00" />
                    <SPLIT distance="50" swimtime="00:01:00.12" />
                    <SPLIT distance="75" swimtime="00:01:34.15" />
                    <SPLIT distance="175" swimtime="00:04:09.06" />
                    <SPLIT distance="200" swimtime="00:04:47.31" />
                    <SPLIT distance="225" swimtime="00:05:21.80" />
                    <SPLIT distance="250" swimtime="00:05:56.81" />
                    <SPLIT distance="275" swimtime="00:06:29.94" />
                    <SPLIT distance="300" swimtime="00:07:05.17" />
                    <SPLIT distance="350" swimtime="00:08:07.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="90" reactiontime="+93" swimtime="00:02:01.62" resultid="110234" heatid="110793" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.97" />
                    <SPLIT distance="50" swimtime="00:00:56.41" />
                    <SPLIT distance="75" swimtime="00:01:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="190" reactiontime="+72" swimtime="00:00:50.09" resultid="110235" heatid="110819" lane="7" entrytime="00:00:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="110219">
              <RESULTS>
                <RESULT eventid="98777" points="246" reactiontime="+80" swimtime="00:00:37.06" resultid="110220" heatid="110588" lane="3" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="193" reactiontime="+88" swimtime="00:13:49.44" resultid="110221" heatid="110634" lane="7" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.56" />
                    <SPLIT distance="50" swimtime="00:00:45.49" />
                    <SPLIT distance="75" swimtime="00:01:10.52" />
                    <SPLIT distance="100" swimtime="00:01:36.70" />
                    <SPLIT distance="125" swimtime="00:02:03.43" />
                    <SPLIT distance="150" swimtime="00:02:30.45" />
                    <SPLIT distance="175" swimtime="00:02:56.75" />
                    <SPLIT distance="200" swimtime="00:03:23.28" />
                    <SPLIT distance="225" swimtime="00:03:49.86" />
                    <SPLIT distance="250" swimtime="00:04:16.50" />
                    <SPLIT distance="275" swimtime="00:04:43.67" />
                    <SPLIT distance="300" swimtime="00:05:10.55" />
                    <SPLIT distance="325" swimtime="00:05:36.91" />
                    <SPLIT distance="350" swimtime="00:06:03.30" />
                    <SPLIT distance="375" swimtime="00:06:30.14" />
                    <SPLIT distance="400" swimtime="00:06:57.31" />
                    <SPLIT distance="425" swimtime="00:07:23.28" />
                    <SPLIT distance="450" swimtime="00:07:49.53" />
                    <SPLIT distance="475" swimtime="00:08:16.09" />
                    <SPLIT distance="500" swimtime="00:08:42.56" />
                    <SPLIT distance="525" swimtime="00:09:08.75" />
                    <SPLIT distance="550" swimtime="00:09:34.82" />
                    <SPLIT distance="575" swimtime="00:10:01.04" />
                    <SPLIT distance="600" swimtime="00:10:27.73" />
                    <SPLIT distance="625" swimtime="00:10:53.14" />
                    <SPLIT distance="650" swimtime="00:11:19.91" />
                    <SPLIT distance="675" swimtime="00:11:45.31" />
                    <SPLIT distance="700" swimtime="00:12:11.44" />
                    <SPLIT distance="725" swimtime="00:12:36.97" />
                    <SPLIT distance="750" swimtime="00:13:03.16" />
                    <SPLIT distance="775" swimtime="00:13:27.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="183" reactiontime="+78" swimtime="00:00:45.21" resultid="110222" heatid="110647" lane="1" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="164" reactiontime="+91" swimtime="00:01:40.48" resultid="110224" heatid="110754" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.82" />
                    <SPLIT distance="75" swimtime="00:01:15.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="197" reactiontime="+61" swimtime="00:03:10.19" resultid="110225" heatid="110765" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.26" />
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="75" swimtime="00:01:09.83" />
                    <SPLIT distance="100" swimtime="00:01:34.47" />
                    <SPLIT distance="125" swimtime="00:01:59.50" />
                    <SPLIT distance="150" swimtime="00:02:24.63" />
                    <SPLIT distance="175" swimtime="00:02:48.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="158" reactiontime="+41" swimtime="00:03:40.17" resultid="110226" heatid="110807" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.69" />
                    <SPLIT distance="50" swimtime="00:00:53.16" />
                    <SPLIT distance="75" swimtime="00:01:20.68" />
                    <SPLIT distance="100" swimtime="00:01:48.69" />
                    <SPLIT distance="125" swimtime="00:02:16.43" />
                    <SPLIT distance="150" swimtime="00:03:40.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="218" reactiontime="+84" swimtime="00:00:47.83" resultid="110227" heatid="110818" lane="5" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="202" reactiontime="+74" swimtime="00:01:36.55" resultid="110353" heatid="110691" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.99" />
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                    <SPLIT distance="75" swimtime="00:01:14.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-11" firstname="Agnieszka" gender="F" lastname="Drejka" nation="POL" athleteid="110236">
              <RESULTS>
                <RESULT eventid="98777" points="218" reactiontime="+84" swimtime="00:00:38.58" resultid="110237" heatid="110587" lane="5" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="196" reactiontime="+85" swimtime="00:03:51.49" resultid="110238" heatid="110662" lane="8" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.51" />
                    <SPLIT distance="50" swimtime="00:00:50.86" />
                    <SPLIT distance="75" swimtime="00:01:19.48" />
                    <SPLIT distance="100" swimtime="00:01:49.01" />
                    <SPLIT distance="125" swimtime="00:02:19.12" />
                    <SPLIT distance="150" swimtime="00:02:50.01" />
                    <SPLIT distance="175" swimtime="00:03:20.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="173" swimtime="00:01:31.34" resultid="110239" heatid="110672" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.12" />
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                    <SPLIT distance="75" swimtime="00:01:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="181" swimtime="00:01:50.10" resultid="110240" heatid="110722" lane="9" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.54" />
                    <SPLIT distance="50" swimtime="00:00:51.36" />
                    <SPLIT distance="75" swimtime="00:01:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="169" reactiontime="+85" swimtime="00:03:19.99" resultid="110241" heatid="110764" lane="4" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.28" />
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                    <SPLIT distance="75" swimtime="00:01:06.75" />
                    <SPLIT distance="100" swimtime="00:01:32.61" />
                    <SPLIT distance="125" swimtime="00:01:59.51" />
                    <SPLIT distance="150" swimtime="00:02:26.79" />
                    <SPLIT distance="175" swimtime="00:02:54.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="180" swimtime="00:00:50.96" resultid="110242" heatid="110819" lane="0" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-14" firstname="Dawid" gender="M" lastname="Zimkowski" nation="POL" athleteid="110243">
              <RESULTS>
                <RESULT eventid="98798" points="354" reactiontime="+72" swimtime="00:00:28.63" resultid="110244" heatid="110604" lane="5" entrytime="00:00:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="271" reactiontime="+94" swimtime="00:02:49.21" resultid="110245" heatid="110623" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.88" />
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="75" swimtime="00:00:55.76" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="125" swimtime="00:01:43.06" />
                    <SPLIT distance="150" swimtime="00:02:09.42" />
                    <SPLIT distance="175" swimtime="00:02:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="110246" heatid="110656" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="110247" heatid="110700" lane="5" entrytime="00:01:15.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="110248" heatid="110747" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="110249" heatid="110760" lane="5" entrytime="00:01:18.00" />
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="110250" heatid="110849" lane="4" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-15" firstname="Mieczysław" gender="M" lastname="Mydłowski" nation="POL" athleteid="110251">
              <RESULTS>
                <RESULT eventid="98798" status="WDR" swimtime="00:00:00.00" resultid="110252" entrytime="00:00:31.00" />
                <RESULT eventid="106277" status="WDR" swimtime="00:00:00.00" resultid="110253" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" status="DNS" swimtime="00:00:00.00" resultid="110254" heatid="110630" lane="8" entrytime="00:02:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110251" number="1" />
                    <RELAYPOSITION athleteid="110236" number="2" />
                    <RELAYPOSITION athleteid="110228" number="3" />
                    <RELAYPOSITION athleteid="110243" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="109310" name="SKP Legia Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1993-01-01" firstname="Krzysztof " gender="M" lastname="Micorek" nation="POL" swrid="4086676" athleteid="109301">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="109311" heatid="110613" lane="9" entrytime="00:00:24.36" entrycourse="SCM" />
                <RESULT eventid="98924" points="355" reactiontime="+59" swimtime="00:00:31.37" resultid="109312" heatid="110659" lane="0" entrytime="00:00:31.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="109313" heatid="110834" lane="1" entrytime="00:00:31.16" entrycourse="SCM" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="109314" heatid="110750" lane="6" entrytime="00:00:27.11" entrycourse="SCM" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="110857" heatid="110797" lane="2" late="yes" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SOPMAST" nation="POL" region="POM" clubid="107683" name="Sopot Masters">
          <CONTACT city="SOPOT" email="sopotmasters@o2.pl" internet="strona www chwilowo nieczynna" name="Gorbaczow Mirosław" phone="696 258 185" state="POMOR" street="ul. Haffnera 57" zip="81-715" />
          <ATHLETES>
            <ATHLETE birthdate="1971-06-03" firstname="Leszek" gender="M" lastname="Wilkowski" nation="POL" athleteid="107684">
              <RESULTS>
                <RESULT eventid="98830" points="242" reactiontime="+99" swimtime="00:02:55.77" resultid="107685" heatid="110622" lane="2" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.79" />
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="75" swimtime="00:00:59.68" />
                    <SPLIT distance="100" swimtime="00:01:21.38" />
                    <SPLIT distance="125" swimtime="00:01:47.78" />
                    <SPLIT distance="150" swimtime="00:02:15.00" />
                    <SPLIT distance="175" swimtime="00:02:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="233" reactiontime="+118" swimtime="00:22:57.69" resultid="107686" heatid="110642" lane="0" entrytime="00:23:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.67" />
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="75" swimtime="00:00:59.54" />
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                    <SPLIT distance="125" swimtime="00:01:43.82" />
                    <SPLIT distance="150" swimtime="00:02:06.42" />
                    <SPLIT distance="175" swimtime="00:02:28.77" />
                    <SPLIT distance="200" swimtime="00:02:52.30" />
                    <SPLIT distance="225" swimtime="00:03:15.21" />
                    <SPLIT distance="250" swimtime="00:03:38.27" />
                    <SPLIT distance="275" swimtime="00:04:01.11" />
                    <SPLIT distance="300" swimtime="00:04:24.47" />
                    <SPLIT distance="325" swimtime="00:04:47.86" />
                    <SPLIT distance="350" swimtime="00:05:11.20" />
                    <SPLIT distance="375" swimtime="00:05:34.99" />
                    <SPLIT distance="400" swimtime="00:05:58.63" />
                    <SPLIT distance="425" swimtime="00:06:21.89" />
                    <SPLIT distance="450" swimtime="00:06:45.34" />
                    <SPLIT distance="475" swimtime="00:07:09.08" />
                    <SPLIT distance="500" swimtime="00:07:32.84" />
                    <SPLIT distance="525" swimtime="00:07:56.48" />
                    <SPLIT distance="550" swimtime="00:08:20.36" />
                    <SPLIT distance="575" swimtime="00:08:43.88" />
                    <SPLIT distance="600" swimtime="00:09:07.73" />
                    <SPLIT distance="625" swimtime="00:09:31.21" />
                    <SPLIT distance="650" swimtime="00:09:54.85" />
                    <SPLIT distance="675" swimtime="00:10:17.86" />
                    <SPLIT distance="700" swimtime="00:10:41.63" />
                    <SPLIT distance="725" swimtime="00:11:05.04" />
                    <SPLIT distance="750" swimtime="00:11:28.52" />
                    <SPLIT distance="775" swimtime="00:11:51.71" />
                    <SPLIT distance="800" swimtime="00:12:14.71" />
                    <SPLIT distance="825" swimtime="00:12:37.22" />
                    <SPLIT distance="850" swimtime="00:13:00.04" />
                    <SPLIT distance="875" swimtime="00:13:23.00" />
                    <SPLIT distance="900" swimtime="00:13:46.14" />
                    <SPLIT distance="925" swimtime="00:14:08.96" />
                    <SPLIT distance="950" swimtime="00:14:32.27" />
                    <SPLIT distance="975" swimtime="00:14:55.18" />
                    <SPLIT distance="1000" swimtime="00:15:18.22" />
                    <SPLIT distance="1025" swimtime="00:15:41.02" />
                    <SPLIT distance="1050" swimtime="00:16:04.42" />
                    <SPLIT distance="1075" swimtime="00:16:27.68" />
                    <SPLIT distance="1100" swimtime="00:16:51.20" />
                    <SPLIT distance="1125" swimtime="00:17:14.39" />
                    <SPLIT distance="1150" swimtime="00:17:37.68" />
                    <SPLIT distance="1175" swimtime="00:18:00.99" />
                    <SPLIT distance="1200" swimtime="00:18:23.99" />
                    <SPLIT distance="1225" swimtime="00:18:46.88" />
                    <SPLIT distance="1250" swimtime="00:19:10.35" />
                    <SPLIT distance="1275" swimtime="00:19:33.59" />
                    <SPLIT distance="1300" swimtime="00:19:57.16" />
                    <SPLIT distance="1325" swimtime="00:20:20.61" />
                    <SPLIT distance="1350" swimtime="00:20:44.91" />
                    <SPLIT distance="1375" swimtime="00:21:07.38" />
                    <SPLIT distance="1400" swimtime="00:21:30.71" />
                    <SPLIT distance="1425" swimtime="00:21:53.54" />
                    <SPLIT distance="1450" swimtime="00:22:16.93" />
                    <SPLIT distance="1475" swimtime="00:22:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="203" reactiontime="+80" swimtime="00:00:37.78" resultid="107687" heatid="110655" lane="8" entrytime="00:00:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="324" reactiontime="+107" swimtime="00:01:05.38" resultid="107688" heatid="110683" lane="4" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.73" />
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="75" swimtime="00:00:47.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="214" reactiontime="+82" swimtime="00:01:21.73" resultid="107689" heatid="110760" lane="6" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.27" />
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="75" swimtime="00:01:01.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="198" swimtime="00:06:43.46" resultid="107690" heatid="110790" lane="0" entrytime="00:06:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.42" />
                    <SPLIT distance="50" swimtime="00:00:45.33" />
                    <SPLIT distance="75" swimtime="00:01:11.21" />
                    <SPLIT distance="100" swimtime="00:01:38.17" />
                    <SPLIT distance="125" swimtime="00:02:05.50" />
                    <SPLIT distance="150" swimtime="00:02:29.87" />
                    <SPLIT distance="175" swimtime="00:02:55.26" />
                    <SPLIT distance="200" swimtime="00:03:21.36" />
                    <SPLIT distance="225" swimtime="00:03:50.54" />
                    <SPLIT distance="250" swimtime="00:04:18.73" />
                    <SPLIT distance="275" swimtime="00:04:47.03" />
                    <SPLIT distance="300" swimtime="00:05:15.96" />
                    <SPLIT distance="325" swimtime="00:05:39.21" />
                    <SPLIT distance="350" swimtime="00:06:01.17" />
                    <SPLIT distance="375" swimtime="00:06:23.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="174" reactiontime="+83" swimtime="00:03:09.06" resultid="107691" heatid="110813" lane="8" entrytime="00:03:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.39" />
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="75" swimtime="00:01:05.13" />
                    <SPLIT distance="125" swimtime="00:01:54.71" />
                    <SPLIT distance="150" swimtime="00:02:20.24" />
                    <SPLIT distance="175" swimtime="00:02:46.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="238" reactiontime="+111" swimtime="00:05:42.40" resultid="107692" heatid="110847" lane="3" entrytime="00:05:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                    <SPLIT distance="75" swimtime="00:00:56.57" />
                    <SPLIT distance="100" swimtime="00:01:17.38" />
                    <SPLIT distance="125" swimtime="00:01:38.33" />
                    <SPLIT distance="150" swimtime="00:02:00.33" />
                    <SPLIT distance="175" swimtime="00:02:22.29" />
                    <SPLIT distance="200" swimtime="00:02:44.34" />
                    <SPLIT distance="225" swimtime="00:03:06.51" />
                    <SPLIT distance="250" swimtime="00:03:29.17" />
                    <SPLIT distance="275" swimtime="00:03:51.39" />
                    <SPLIT distance="300" swimtime="00:04:14.13" />
                    <SPLIT distance="325" swimtime="00:04:36.24" />
                    <SPLIT distance="350" swimtime="00:04:59.33" />
                    <SPLIT distance="375" swimtime="00:05:22.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-20" firstname="Piotr" gender="M" lastname="Suwara" nation="POL" athleteid="107693">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="107694" heatid="110607" lane="5" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="98891" points="316" reactiontime="+97" swimtime="00:10:50.97" resultid="107695" heatid="110636" lane="3" entrytime="00:10:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.35" />
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="75" swimtime="00:00:55.77" />
                    <SPLIT distance="100" swimtime="00:01:15.88" />
                    <SPLIT distance="125" swimtime="00:01:36.50" />
                    <SPLIT distance="150" swimtime="00:01:57.15" />
                    <SPLIT distance="175" swimtime="00:02:17.95" />
                    <SPLIT distance="200" swimtime="00:02:38.66" />
                    <SPLIT distance="225" swimtime="00:02:59.54" />
                    <SPLIT distance="250" swimtime="00:03:20.41" />
                    <SPLIT distance="275" swimtime="00:03:41.50" />
                    <SPLIT distance="300" swimtime="00:04:02.30" />
                    <SPLIT distance="325" swimtime="00:04:23.27" />
                    <SPLIT distance="350" swimtime="00:04:44.17" />
                    <SPLIT distance="375" swimtime="00:05:05.16" />
                    <SPLIT distance="400" swimtime="00:05:25.80" />
                    <SPLIT distance="425" swimtime="00:05:46.50" />
                    <SPLIT distance="450" swimtime="00:06:07.07" />
                    <SPLIT distance="475" swimtime="00:06:28.01" />
                    <SPLIT distance="500" swimtime="00:06:49.27" />
                    <SPLIT distance="525" swimtime="00:07:10.11" />
                    <SPLIT distance="550" swimtime="00:07:30.81" />
                    <SPLIT distance="575" swimtime="00:07:51.83" />
                    <SPLIT distance="600" swimtime="00:08:12.10" />
                    <SPLIT distance="625" swimtime="00:08:32.28" />
                    <SPLIT distance="650" swimtime="00:08:52.55" />
                    <SPLIT distance="675" swimtime="00:09:12.58" />
                    <SPLIT distance="700" swimtime="00:09:32.74" />
                    <SPLIT distance="725" swimtime="00:09:52.44" />
                    <SPLIT distance="750" swimtime="00:10:12.35" />
                    <SPLIT distance="775" swimtime="00:10:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="273" reactiontime="+87" swimtime="00:00:34.23" resultid="107696" heatid="110655" lane="6" entrytime="00:00:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="365" swimtime="00:01:02.87" resultid="107697" heatid="110686" lane="0" entrytime="00:01:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.26" />
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="75" swimtime="00:00:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="317" reactiontime="+88" swimtime="00:01:11.69" resultid="107698" heatid="110761" lane="9" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.22" />
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="75" swimtime="00:00:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="356" reactiontime="+91" swimtime="00:02:20.11" resultid="107699" heatid="110775" lane="8" entrytime="00:02:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.93" />
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="75" swimtime="00:00:49.59" />
                    <SPLIT distance="100" swimtime="00:01:07.50" />
                    <SPLIT distance="125" swimtime="00:01:25.82" />
                    <SPLIT distance="150" swimtime="00:01:44.53" />
                    <SPLIT distance="175" swimtime="00:02:02.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="305" reactiontime="+92" swimtime="00:02:36.85" resultid="107700" heatid="110814" lane="5" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.67" />
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="75" swimtime="00:00:56.08" />
                    <SPLIT distance="100" swimtime="00:01:16.17" />
                    <SPLIT distance="125" swimtime="00:01:36.27" />
                    <SPLIT distance="150" swimtime="00:01:56.83" />
                    <SPLIT distance="175" swimtime="00:02:17.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="327" reactiontime="+93" swimtime="00:05:08.07" resultid="107701" heatid="110846" lane="4" entrytime="00:05:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.77" />
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="75" swimtime="00:00:52.82" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="125" swimtime="00:01:31.71" />
                    <SPLIT distance="150" swimtime="00:01:51.62" />
                    <SPLIT distance="175" swimtime="00:02:11.51" />
                    <SPLIT distance="200" swimtime="00:02:31.49" />
                    <SPLIT distance="225" swimtime="00:02:51.40" />
                    <SPLIT distance="250" swimtime="00:03:11.46" />
                    <SPLIT distance="275" swimtime="00:03:31.50" />
                    <SPLIT distance="300" swimtime="00:03:51.62" />
                    <SPLIT distance="325" swimtime="00:04:11.32" />
                    <SPLIT distance="350" swimtime="00:04:31.06" />
                    <SPLIT distance="375" swimtime="00:04:50.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="109146" name="SPK Kúpele Piešťany– KUPI ">
          <ATHLETES>
            <ATHLETE birthdate="1969-10-28" firstname=" Pavel" gender="M" lastname="Škodný" nation="SVK" athleteid="109169">
              <RESULTS>
                <RESULT eventid="98924" points="290" reactiontime="+81" swimtime="00:00:33.56" resultid="109170" heatid="110657" lane="1" entrytime="00:00:33.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="290" reactiontime="+95" swimtime="00:02:43.92" resultid="109171" heatid="110712" lane="3" entrytime="00:02:49.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.35" />
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="75" swimtime="00:00:55.89" />
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                    <SPLIT distance="125" swimtime="00:01:38.35" />
                    <SPLIT distance="150" swimtime="00:02:00.06" />
                    <SPLIT distance="175" swimtime="00:02:22.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="318" reactiontime="+76" swimtime="00:01:11.60" resultid="109172" heatid="110762" lane="8" entrytime="00:01:11.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.15" />
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="75" swimtime="00:00:53.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="340" reactiontime="+98" swimtime="00:05:37.16" resultid="109173" heatid="110791" lane="5" entrytime="00:05:39.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.96" />
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="75" swimtime="00:00:55.50" />
                    <SPLIT distance="100" swimtime="00:01:16.77" />
                    <SPLIT distance="125" swimtime="00:01:38.72" />
                    <SPLIT distance="150" swimtime="00:02:00.41" />
                    <SPLIT distance="175" swimtime="00:02:21.99" />
                    <SPLIT distance="200" swimtime="00:02:43.12" />
                    <SPLIT distance="225" swimtime="00:03:07.72" />
                    <SPLIT distance="250" swimtime="00:03:33.33" />
                    <SPLIT distance="275" swimtime="00:03:57.49" />
                    <SPLIT distance="300" swimtime="00:04:22.87" />
                    <SPLIT distance="325" swimtime="00:04:42.24" />
                    <SPLIT distance="350" swimtime="00:05:01.35" />
                    <SPLIT distance="375" swimtime="00:05:20.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="318" reactiontime="+84" swimtime="00:02:34.62" resultid="109174" heatid="110815" lane="1" entrytime="00:02:35.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.03" />
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="75" swimtime="00:00:55.39" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="125" swimtime="00:01:35.14" />
                    <SPLIT distance="150" swimtime="00:01:55.52" />
                    <SPLIT distance="175" swimtime="00:02:15.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-04-21" firstname=" Anna" gender="F" lastname="Kičinova " nation="SVK" athleteid="109175">
              <RESULTS>
                <RESULT eventid="98940" points="276" reactiontime="+118" swimtime="00:03:26.55" resultid="109176" heatid="110663" lane="2" entrytime="00:03:24.94">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.75" />
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="75" swimtime="00:01:11.63" />
                    <SPLIT distance="100" swimtime="00:01:37.76" />
                    <SPLIT distance="125" swimtime="00:02:04.17" />
                    <SPLIT distance="150" swimtime="00:02:31.42" />
                    <SPLIT distance="175" swimtime="00:02:59.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="207" reactiontime="+90" swimtime="00:03:22.12" resultid="109177" heatid="110708" lane="6" entrytime="00:03:14.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.49" />
                    <SPLIT distance="50" swimtime="00:00:43.57" />
                    <SPLIT distance="75" swimtime="00:01:07.88" />
                    <SPLIT distance="100" swimtime="00:01:32.99" />
                    <SPLIT distance="125" swimtime="00:01:58.61" />
                    <SPLIT distance="150" swimtime="00:02:25.99" />
                    <SPLIT distance="175" swimtime="00:02:52.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="280" swimtime="00:01:35.26" resultid="109178" heatid="110723" lane="4" entrytime="00:01:34.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.19" />
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                    <SPLIT distance="75" swimtime="00:01:10.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="238" reactiontime="+88" swimtime="00:00:39.32" resultid="109179" heatid="110738" lane="8" entrytime="00:00:38.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="247" reactiontime="+89" swimtime="00:01:26.98" resultid="109180" heatid="110795" lane="8" entrytime="00:01:27.03">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.65" />
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="75" swimtime="00:01:02.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="270" swimtime="00:00:44.51" resultid="109181" heatid="110820" lane="4" entrytime="00:00:43.74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="106496" name="Start Poznań">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" phone="512111513" street="os. Batorego 8/67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1964-06-06" firstname="Krzysztof" gender="M" lastname="Kapałczyński" nation="POL" athleteid="106511">
              <RESULTS>
                <RESULT eventid="98830" points="302" reactiontime="+104" swimtime="00:02:43.23" resultid="110263" heatid="110624" lane="0" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.07" />
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="75" swimtime="00:00:57.43" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="125" swimtime="00:01:41.61" />
                    <SPLIT distance="150" swimtime="00:02:05.84" />
                    <SPLIT distance="175" swimtime="00:02:25.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="223" reactiontime="+82" swimtime="00:02:58.92" resultid="110264" heatid="110712" lane="7" entrytime="00:02:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.69" />
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="75" swimtime="00:01:00.37" />
                    <SPLIT distance="100" swimtime="00:01:24.12" />
                    <SPLIT distance="125" swimtime="00:01:47.68" />
                    <SPLIT distance="150" swimtime="00:02:12.01" />
                    <SPLIT distance="175" swimtime="00:02:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="110265" heatid="110732" lane="4" entrytime="00:01:20.00" entrycourse="SCM" />
                <RESULT eventid="99282" points="291" swimtime="00:05:55.05" resultid="110266" heatid="110791" lane="0" entrytime="00:05:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.00" />
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="75" swimtime="00:00:57.17" />
                    <SPLIT distance="100" swimtime="00:01:20.09" />
                    <SPLIT distance="125" swimtime="00:01:44.41" />
                    <SPLIT distance="150" swimtime="00:02:07.53" />
                    <SPLIT distance="175" swimtime="00:02:30.14" />
                    <SPLIT distance="200" swimtime="00:02:52.73" />
                    <SPLIT distance="225" swimtime="00:03:18.07" />
                    <SPLIT distance="250" swimtime="00:03:43.97" />
                    <SPLIT distance="275" swimtime="00:04:08.64" />
                    <SPLIT distance="300" swimtime="00:04:34.31" />
                    <SPLIT distance="325" swimtime="00:04:55.28" />
                    <SPLIT distance="350" swimtime="00:05:16.68" />
                    <SPLIT distance="375" swimtime="00:05:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="261" swimtime="00:01:15.73" resultid="110267" heatid="110801" lane="6" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.50" />
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="75" swimtime="00:00:55.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="267" swimtime="00:00:39.19" resultid="110268" heatid="110830" lane="0" entrytime="00:00:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-06-06" firstname="Anna" gender="F" lastname="Rostkowska-Kaczmarek" nation="POL" athleteid="106557">
              <RESULTS>
                <RESULT eventid="98777" points="307" reactiontime="+96" swimtime="00:00:34.44" resultid="110303" heatid="110589" lane="3" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="265" reactiontime="+102" swimtime="00:01:19.25" resultid="110304" heatid="110673" lane="7" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.98" />
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="75" swimtime="00:00:57.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="110305" heatid="110692" lane="7" entrytime="00:01:32.00" />
                <RESULT eventid="99154" points="217" reactiontime="+96" swimtime="00:00:40.54" resultid="110306" heatid="110737" lane="7" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="215" swimtime="00:03:04.80" resultid="110307" heatid="110765" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.50" />
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                    <SPLIT distance="75" swimtime="00:01:05.08" />
                    <SPLIT distance="100" swimtime="00:01:28.98" />
                    <SPLIT distance="150" swimtime="00:02:17.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="258" swimtime="00:00:45.19" resultid="110308" heatid="110820" lane="9" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="206" reactiontime="+98" swimtime="00:06:36.50" resultid="110309" heatid="110842" lane="5" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.20" />
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                    <SPLIT distance="75" swimtime="00:01:07.97" />
                    <SPLIT distance="100" swimtime="00:01:32.99" />
                    <SPLIT distance="125" swimtime="00:01:57.83" />
                    <SPLIT distance="150" swimtime="00:02:22.83" />
                    <SPLIT distance="175" swimtime="00:03:40.28" />
                    <SPLIT distance="200" swimtime="00:03:14.01" />
                    <SPLIT distance="225" swimtime="00:05:22.88" />
                    <SPLIT distance="250" swimtime="00:04:57.99" />
                    <SPLIT distance="275" swimtime="00:06:13.14" />
                    <SPLIT distance="300" swimtime="00:05:48.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-06-06" firstname="Maja" gender="F" lastname="Spychalska" nation="POL" athleteid="106535">
              <RESULTS>
                <RESULT eventid="98777" points="458" reactiontime="+85" swimtime="00:00:30.14" resultid="110284" heatid="110590" lane="6" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" status="DNS" swimtime="00:00:00.00" resultid="110285" heatid="110649" lane="0" entrytime="00:00:39.00" />
                <RESULT eventid="99409" points="444" swimtime="00:00:37.74" resultid="110286" heatid="110822" lane="2" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-06" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="106502">
              <RESULTS>
                <RESULT eventid="98798" points="495" reactiontime="+79" swimtime="00:00:25.61" resultid="110255" heatid="110609" lane="4" entrytime="00:00:26.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="110256" heatid="110626" lane="1" entrytime="00:02:35.00" entrycourse="SCM" />
                <RESULT eventid="106277" points="489" reactiontime="+90" swimtime="00:00:57.02" resultid="110257" heatid="110678" lane="1" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                    <SPLIT distance="75" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="500" reactiontime="+85" swimtime="00:01:03.80" resultid="110258" heatid="110705" lane="3" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.24" />
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                    <SPLIT distance="75" swimtime="00:00:48.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="460" reactiontime="+81" swimtime="00:00:28.22" resultid="110259" heatid="110749" lane="8" entrytime="00:00:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="413" reactiontime="+66" swimtime="00:01:05.65" resultid="110260" heatid="110763" lane="0" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.24" />
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="75" swimtime="00:00:48.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="462" swimtime="00:01:02.64" resultid="110261" heatid="110803" lane="3" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.43" />
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                    <SPLIT distance="75" swimtime="00:00:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="110262" heatid="110816" lane="0" entrytime="00:02:25.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-06" firstname="Aneta" gender="F" lastname="Maduzia" nation="POL" athleteid="106548">
              <RESULTS>
                <RESULT eventid="98777" points="346" reactiontime="+97" swimtime="00:00:33.09" resultid="110295" heatid="110590" lane="1" entrytime="00:00:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="290" reactiontime="+99" swimtime="00:12:03.60" resultid="110296" heatid="110633" lane="0" entrytime="00:11:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.49" />
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="75" swimtime="00:01:03.52" />
                    <SPLIT distance="100" swimtime="00:01:25.92" />
                    <SPLIT distance="125" swimtime="00:01:48.65" />
                    <SPLIT distance="150" swimtime="00:02:11.55" />
                    <SPLIT distance="175" swimtime="00:02:34.18" />
                    <SPLIT distance="200" swimtime="00:02:57.00" />
                    <SPLIT distance="225" swimtime="00:03:19.48" />
                    <SPLIT distance="250" swimtime="00:03:42.43" />
                    <SPLIT distance="275" swimtime="00:04:05.00" />
                    <SPLIT distance="300" swimtime="00:04:28.04" />
                    <SPLIT distance="325" swimtime="00:04:51.10" />
                    <SPLIT distance="350" swimtime="00:05:14.26" />
                    <SPLIT distance="375" swimtime="00:05:37.02" />
                    <SPLIT distance="400" swimtime="00:06:00.09" />
                    <SPLIT distance="425" swimtime="00:06:22.90" />
                    <SPLIT distance="450" swimtime="00:06:45.68" />
                    <SPLIT distance="475" swimtime="00:07:08.19" />
                    <SPLIT distance="500" swimtime="00:07:30.69" />
                    <SPLIT distance="525" swimtime="00:07:53.70" />
                    <SPLIT distance="550" swimtime="00:08:16.60" />
                    <SPLIT distance="575" swimtime="00:08:39.47" />
                    <SPLIT distance="600" swimtime="00:09:02.35" />
                    <SPLIT distance="625" swimtime="00:09:25.05" />
                    <SPLIT distance="650" swimtime="00:09:48.38" />
                    <SPLIT distance="675" swimtime="00:10:11.23" />
                    <SPLIT distance="700" swimtime="00:10:33.95" />
                    <SPLIT distance="725" swimtime="00:10:56.55" />
                    <SPLIT distance="750" swimtime="00:11:19.85" />
                    <SPLIT distance="775" swimtime="00:11:42.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="345" reactiontime="+88" swimtime="00:01:12.55" resultid="110297" heatid="110674" lane="5" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.42" />
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="75" swimtime="00:00:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="238" reactiontime="+93" swimtime="00:03:12.78" resultid="110298" heatid="110708" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.54" />
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                    <SPLIT distance="75" swimtime="00:01:08.34" />
                    <SPLIT distance="100" swimtime="00:01:33.19" />
                    <SPLIT distance="125" swimtime="00:01:57.93" />
                    <SPLIT distance="150" swimtime="00:02:23.36" />
                    <SPLIT distance="175" swimtime="00:02:48.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="318" reactiontime="+90" swimtime="00:00:35.69" resultid="110299" heatid="110738" lane="4" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="309" reactiontime="+90" swimtime="00:02:43.74" resultid="110300" heatid="110766" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.87" />
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="75" swimtime="00:00:58.75" />
                    <SPLIT distance="100" swimtime="00:01:19.72" />
                    <SPLIT distance="125" swimtime="00:01:41.04" />
                    <SPLIT distance="150" swimtime="00:02:02.79" />
                    <SPLIT distance="175" swimtime="00:02:23.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="278" reactiontime="+95" swimtime="00:01:23.61" resultid="110301" heatid="110795" lane="1" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.08" />
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="75" swimtime="00:01:01.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="294" reactiontime="+91" swimtime="00:05:52.45" resultid="110302" heatid="110840" lane="1" entrytime="00:05:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.01" />
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="75" swimtime="00:01:01.77" />
                    <SPLIT distance="100" swimtime="00:01:23.97" />
                    <SPLIT distance="125" swimtime="00:01:46.42" />
                    <SPLIT distance="150" swimtime="00:02:09.05" />
                    <SPLIT distance="175" swimtime="00:02:31.44" />
                    <SPLIT distance="200" swimtime="00:02:53.65" />
                    <SPLIT distance="225" swimtime="00:03:16.03" />
                    <SPLIT distance="250" swimtime="00:03:38.85" />
                    <SPLIT distance="275" swimtime="00:04:01.07" />
                    <SPLIT distance="300" swimtime="00:04:23.39" />
                    <SPLIT distance="325" swimtime="00:04:45.76" />
                    <SPLIT distance="350" swimtime="00:05:08.21" />
                    <SPLIT distance="375" swimtime="00:05:30.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-06" firstname="Joanna" gender="F" lastname="Kostencka" nation="POL" athleteid="106526">
              <RESULTS>
                <RESULT eventid="98814" points="414" reactiontime="+107" swimtime="00:02:43.43" resultid="110276" heatid="110615" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.92" />
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="75" swimtime="00:00:56.45" />
                    <SPLIT distance="100" swimtime="00:01:15.93" />
                    <SPLIT distance="125" swimtime="00:01:40.39" />
                    <SPLIT distance="150" swimtime="00:02:05.60" />
                    <SPLIT distance="175" swimtime="00:02:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="395" reactiontime="+95" swimtime="00:10:52.89" resultid="110277" heatid="110633" lane="7" entrytime="00:11:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.54" />
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="75" swimtime="00:00:56.37" />
                    <SPLIT distance="100" swimtime="00:01:16.11" />
                    <SPLIT distance="125" swimtime="00:01:36.17" />
                    <SPLIT distance="150" swimtime="00:01:56.43" />
                    <SPLIT distance="175" swimtime="00:02:16.77" />
                    <SPLIT distance="200" swimtime="00:02:37.37" />
                    <SPLIT distance="225" swimtime="00:02:57.98" />
                    <SPLIT distance="250" swimtime="00:03:18.52" />
                    <SPLIT distance="275" swimtime="00:03:39.16" />
                    <SPLIT distance="300" swimtime="00:04:00.09" />
                    <SPLIT distance="325" swimtime="00:04:20.94" />
                    <SPLIT distance="350" swimtime="00:04:41.81" />
                    <SPLIT distance="375" swimtime="00:05:02.56" />
                    <SPLIT distance="400" swimtime="00:05:23.49" />
                    <SPLIT distance="425" swimtime="00:05:44.39" />
                    <SPLIT distance="450" swimtime="00:06:05.40" />
                    <SPLIT distance="475" swimtime="00:06:26.13" />
                    <SPLIT distance="500" swimtime="00:06:47.14" />
                    <SPLIT distance="525" swimtime="00:07:08.10" />
                    <SPLIT distance="550" swimtime="00:07:28.91" />
                    <SPLIT distance="575" swimtime="00:07:49.37" />
                    <SPLIT distance="600" swimtime="00:08:10.09" />
                    <SPLIT distance="625" swimtime="00:08:30.58" />
                    <SPLIT distance="650" swimtime="00:08:50.97" />
                    <SPLIT distance="675" swimtime="00:09:11.36" />
                    <SPLIT distance="700" swimtime="00:09:31.94" />
                    <SPLIT distance="725" swimtime="00:09:52.70" />
                    <SPLIT distance="750" swimtime="00:10:13.09" />
                    <SPLIT distance="775" swimtime="00:10:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="403" reactiontime="+79" swimtime="00:00:34.73" resultid="110278" heatid="110649" lane="4" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="454" swimtime="00:01:06.23" resultid="110279" heatid="110675" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.62" />
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="75" swimtime="00:00:49.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="426" reactiontime="+89" swimtime="00:01:13.12" resultid="110280" heatid="110755" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.72" />
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="75" swimtime="00:00:54.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="448" reactiontime="+93" swimtime="00:02:24.75" resultid="110281" heatid="110767" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.11" />
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="75" swimtime="00:00:51.91" />
                    <SPLIT distance="100" swimtime="00:01:10.40" />
                    <SPLIT distance="125" swimtime="00:01:28.96" />
                    <SPLIT distance="150" swimtime="00:01:47.71" />
                    <SPLIT distance="175" swimtime="00:02:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="439" reactiontime="+85" swimtime="00:02:36.87" resultid="110282" heatid="110809" lane="5" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.46" />
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="75" swimtime="00:00:57.12" />
                    <SPLIT distance="100" swimtime="00:01:17.00" />
                    <SPLIT distance="125" swimtime="00:01:37.08" />
                    <SPLIT distance="150" swimtime="00:01:57.39" />
                    <SPLIT distance="175" swimtime="00:02:17.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="402" reactiontime="+98" swimtime="00:05:17.76" resultid="110283" heatid="110841" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.30" />
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                    <SPLIT distance="75" swimtime="00:00:56.41" />
                    <SPLIT distance="100" swimtime="00:01:16.27" />
                    <SPLIT distance="125" swimtime="00:01:36.44" />
                    <SPLIT distance="150" swimtime="00:01:56.69" />
                    <SPLIT distance="175" swimtime="00:02:17.23" />
                    <SPLIT distance="200" swimtime="00:02:37.09" />
                    <SPLIT distance="225" swimtime="00:02:57.69" />
                    <SPLIT distance="250" swimtime="00:03:17.92" />
                    <SPLIT distance="275" swimtime="00:03:38.45" />
                    <SPLIT distance="300" swimtime="00:03:58.72" />
                    <SPLIT distance="325" swimtime="00:04:19.04" />
                    <SPLIT distance="350" swimtime="00:04:39.30" />
                    <SPLIT distance="375" swimtime="00:04:59.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-06" firstname="Joanna" gender="F" lastname="Krzyśków" nation="POL" athleteid="106565">
              <RESULTS>
                <RESULT comment="Z-2G3" eventid="98972" status="DSQ" swimtime="00:00:00.00" resultid="110310" heatid="110693" lane="6" entrytime="00:01:25.00" />
                <RESULT eventid="99089" points="349" reactiontime="+92" swimtime="00:01:28.55" resultid="110311" heatid="110724" lane="5" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.23" />
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="75" swimtime="00:01:04.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="290" reactiontime="+98" swimtime="00:00:36.80" resultid="110312" heatid="110738" lane="2" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="350" reactiontime="+107" swimtime="00:00:40.86" resultid="110865" heatid="110822" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-06-06" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="106518">
              <RESULTS>
                <RESULT eventid="98798" points="446" reactiontime="+77" swimtime="00:00:26.50" resultid="110269" heatid="110608" lane="4" entrytime="00:00:27.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="397" reactiontime="+59" swimtime="00:02:29.16" resultid="110270" heatid="110627" lane="7" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.54" />
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="75" swimtime="00:00:51.90" />
                    <SPLIT distance="100" swimtime="00:01:11.04" />
                    <SPLIT distance="125" swimtime="00:01:32.92" />
                    <SPLIT distance="150" swimtime="00:01:55.50" />
                    <SPLIT distance="175" swimtime="00:02:13.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="490" reactiontime="+61" swimtime="00:00:56.98" resultid="110271" heatid="110688" lane="7" entrytime="00:00:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.43" />
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="75" swimtime="00:00:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="422" reactiontime="+76" swimtime="00:01:07.52" resultid="110272" heatid="110704" lane="2" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="75" swimtime="00:00:51.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="478" swimtime="00:02:07.04" resultid="110273" heatid="110777" lane="6" entrytime="00:02:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.09" />
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="75" swimtime="00:00:46.61" />
                    <SPLIT distance="100" swimtime="00:01:02.68" />
                    <SPLIT distance="125" swimtime="00:01:18.87" />
                    <SPLIT distance="150" swimtime="00:01:35.09" />
                    <SPLIT distance="175" swimtime="00:01:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="376" reactiontime="+87" swimtime="00:05:26.00" resultid="110274" heatid="110791" lane="4" entrytime="00:05:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.52" />
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="75" swimtime="00:00:53.63" />
                    <SPLIT distance="100" swimtime="00:01:13.76" />
                    <SPLIT distance="125" swimtime="00:01:35.88" />
                    <SPLIT distance="150" swimtime="00:01:56.62" />
                    <SPLIT distance="175" swimtime="00:02:17.81" />
                    <SPLIT distance="200" swimtime="00:02:38.88" />
                    <SPLIT distance="225" swimtime="00:03:02.93" />
                    <SPLIT distance="250" swimtime="00:03:26.81" />
                    <SPLIT distance="275" swimtime="00:03:51.23" />
                    <SPLIT distance="300" swimtime="00:04:16.81" />
                    <SPLIT distance="325" swimtime="00:04:34.26" />
                    <SPLIT distance="350" swimtime="00:04:51.80" />
                    <SPLIT distance="375" swimtime="00:05:09.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="433" swimtime="00:04:40.40" resultid="110275" heatid="110844" lane="6" entrytime="00:04:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="75" swimtime="00:00:50.07" />
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                    <SPLIT distance="125" swimtime="00:01:26.32" />
                    <SPLIT distance="150" swimtime="00:01:43.98" />
                    <SPLIT distance="175" swimtime="00:02:01.93" />
                    <SPLIT distance="200" swimtime="00:02:20.10" />
                    <SPLIT distance="225" swimtime="00:02:38.16" />
                    <SPLIT distance="250" swimtime="00:02:56.24" />
                    <SPLIT distance="275" swimtime="00:03:14.34" />
                    <SPLIT distance="300" swimtime="00:03:32.75" />
                    <SPLIT distance="325" swimtime="00:03:50.01" />
                    <SPLIT distance="350" swimtime="00:04:07.62" />
                    <SPLIT distance="375" swimtime="00:04:24.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-06-06" firstname="Mateusz" gender="M" lastname="Pałczyński" nation="POL" athleteid="106539">
              <RESULTS>
                <RESULT eventid="98830" points="359" reactiontime="+70" swimtime="00:02:34.18" resultid="110287" heatid="110626" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.80" />
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="75" swimtime="00:00:50.44" />
                    <SPLIT distance="100" swimtime="00:01:10.10" />
                    <SPLIT distance="125" swimtime="00:01:31.04" />
                    <SPLIT distance="150" swimtime="00:01:53.63" />
                    <SPLIT distance="175" swimtime="00:02:14.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="225" reactiontime="+100" swimtime="00:12:08.23" resultid="110288" heatid="110635" lane="3" entrytime="00:09:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.00" />
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="75" swimtime="00:00:54.46" />
                    <SPLIT distance="100" swimtime="00:01:14.28" />
                    <SPLIT distance="125" swimtime="00:01:34.13" />
                    <SPLIT distance="150" swimtime="00:01:54.44" />
                    <SPLIT distance="175" swimtime="00:02:14.99" />
                    <SPLIT distance="200" swimtime="00:02:36.31" />
                    <SPLIT distance="225" swimtime="00:02:57.25" />
                    <SPLIT distance="250" swimtime="00:03:19.04" />
                    <SPLIT distance="275" swimtime="00:03:41.46" />
                    <SPLIT distance="300" swimtime="00:04:05.24" />
                    <SPLIT distance="325" swimtime="00:04:27.89" />
                    <SPLIT distance="350" swimtime="00:04:50.82" />
                    <SPLIT distance="375" swimtime="00:05:14.32" />
                    <SPLIT distance="400" swimtime="00:05:38.14" />
                    <SPLIT distance="425" swimtime="00:06:02.86" />
                    <SPLIT distance="450" swimtime="00:06:26.95" />
                    <SPLIT distance="475" swimtime="00:06:50.90" />
                    <SPLIT distance="500" swimtime="00:07:14.20" />
                    <SPLIT distance="525" swimtime="00:07:38.65" />
                    <SPLIT distance="550" swimtime="00:08:03.19" />
                    <SPLIT distance="575" swimtime="00:08:28.87" />
                    <SPLIT distance="600" swimtime="00:08:53.02" />
                    <SPLIT distance="625" swimtime="00:09:17.93" />
                    <SPLIT distance="650" swimtime="00:09:43.19" />
                    <SPLIT distance="675" swimtime="00:10:08.34" />
                    <SPLIT distance="700" swimtime="00:10:32.65" />
                    <SPLIT distance="725" swimtime="00:10:57.18" />
                    <SPLIT distance="750" swimtime="00:11:21.03" />
                    <SPLIT distance="775" swimtime="00:11:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="349" reactiontime="+43" swimtime="00:02:51.04" resultid="110289" heatid="110670" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.89" />
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="75" swimtime="00:00:56.63" />
                    <SPLIT distance="100" swimtime="00:01:17.72" />
                    <SPLIT distance="125" swimtime="00:01:39.80" />
                    <SPLIT distance="150" swimtime="00:02:02.69" />
                    <SPLIT distance="175" swimtime="00:02:26.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="252" swimtime="00:02:51.72" resultid="110290" heatid="110713" lane="9" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.72" />
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="75" swimtime="00:00:57.80" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="125" swimtime="00:01:40.40" />
                    <SPLIT distance="150" swimtime="00:02:03.25" />
                    <SPLIT distance="175" swimtime="00:02:27.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="458" reactiontime="+78" swimtime="00:01:12.13" resultid="110291" heatid="110733" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.35" />
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="75" swimtime="00:00:52.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="299" reactiontime="+92" swimtime="00:05:52.02" resultid="110292" heatid="110792" lane="7" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.95" />
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="75" swimtime="00:00:53.74" />
                    <SPLIT distance="100" swimtime="00:01:15.14" />
                    <SPLIT distance="125" swimtime="00:01:37.65" />
                    <SPLIT distance="150" swimtime="00:01:59.74" />
                    <SPLIT distance="175" swimtime="00:02:21.96" />
                    <SPLIT distance="200" swimtime="00:02:45.21" />
                    <SPLIT distance="225" swimtime="00:03:09.14" />
                    <SPLIT distance="250" swimtime="00:03:33.26" />
                    <SPLIT distance="275" swimtime="00:03:57.53" />
                    <SPLIT distance="300" swimtime="00:04:22.81" />
                    <SPLIT distance="325" swimtime="00:04:46.03" />
                    <SPLIT distance="350" swimtime="00:05:08.35" />
                    <SPLIT distance="375" swimtime="00:05:30.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="246" reactiontime="+105" swimtime="00:02:48.39" resultid="110293" heatid="110814" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.68" />
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="75" swimtime="00:00:58.75" />
                    <SPLIT distance="100" swimtime="00:01:19.52" />
                    <SPLIT distance="125" swimtime="00:01:40.91" />
                    <SPLIT distance="150" swimtime="00:02:02.84" />
                    <SPLIT distance="175" swimtime="00:02:25.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="466" swimtime="00:00:32.55" resultid="110294" heatid="110834" lane="9" entrytime="00:00:32.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="394" reactiontime="+74" swimtime="00:02:03.41" resultid="110315" heatid="110718" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.23" />
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="75" swimtime="00:00:45.46" />
                    <SPLIT distance="100" swimtime="00:01:03.21" />
                    <SPLIT distance="125" swimtime="00:01:18.32" />
                    <SPLIT distance="150" swimtime="00:01:36.87" />
                    <SPLIT distance="175" swimtime="00:01:49.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106502" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="106539" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="106511" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="106518" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="99250" points="422" swimtime="00:01:50.09" resultid="110318" heatid="110783" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.96" />
                    <SPLIT distance="50" swimtime="00:00:26.12" />
                    <SPLIT distance="75" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:00:56.16" />
                    <SPLIT distance="125" swimtime="00:01:08.98" />
                    <SPLIT distance="150" swimtime="00:01:23.12" />
                    <SPLIT distance="175" swimtime="00:01:36.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106502" number="1" />
                    <RELAYPOSITION athleteid="106511" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="106539" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="106518" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="99036" points="404" reactiontime="+93" swimtime="00:02:20.70" resultid="110314" heatid="110715" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.30" />
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="75" swimtime="00:00:53.22" />
                    <SPLIT distance="100" swimtime="00:01:14.98" />
                    <SPLIT distance="125" swimtime="00:01:31.29" />
                    <SPLIT distance="150" swimtime="00:01:50.70" />
                    <SPLIT distance="175" swimtime="00:02:05.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106526" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="106565" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="106548" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="106535" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="99234" points="384" reactiontime="+88" swimtime="00:02:09.59" resultid="110317" heatid="110780" lane="7" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.18" />
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="75" swimtime="00:00:47.82" />
                    <SPLIT distance="100" swimtime="00:01:06.20" />
                    <SPLIT distance="125" swimtime="00:01:22.08" />
                    <SPLIT distance="150" swimtime="00:01:39.60" />
                    <SPLIT distance="175" swimtime="00:01:54.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106526" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="106565" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="106548" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="106535" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="99441" points="381" reactiontime="+87" swimtime="00:02:04.75" resultid="110316" heatid="110838" lane="2" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.35" />
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="75" swimtime="00:00:49.75" />
                    <SPLIT distance="100" swimtime="00:01:07.16" />
                    <SPLIT distance="125" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:01:35.01" />
                    <SPLIT distance="175" swimtime="00:01:49.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106526" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="106539" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="106502" number="3" />
                    <RELAYPOSITION athleteid="106535" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="107087" name="Steef Wroclaw">
          <CONTACT city="rocław" email="ste1@wp.pl" name="Skrzypek Stefan" phone="500388374" street="Edyty Stein 6/1" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="107095">
              <RESULTS>
                <RESULT eventid="98830" points="182" reactiontime="+106" swimtime="00:03:13.13" resultid="107096" heatid="110622" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.09" />
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="75" swimtime="00:01:08.79" />
                    <SPLIT distance="100" swimtime="00:01:34.66" />
                    <SPLIT distance="125" swimtime="00:02:02.28" />
                    <SPLIT distance="150" swimtime="00:02:30.30" />
                    <SPLIT distance="175" swimtime="00:02:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="198" reactiontime="+105" swimtime="00:24:13.44" resultid="107097" heatid="110643" lane="2" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.27" />
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="75" swimtime="00:01:05.62" />
                    <SPLIT distance="100" swimtime="00:01:28.52" />
                    <SPLIT distance="125" swimtime="00:01:51.65" />
                    <SPLIT distance="150" swimtime="00:02:14.90" />
                    <SPLIT distance="175" swimtime="00:02:38.53" />
                    <SPLIT distance="200" swimtime="00:03:02.80" />
                    <SPLIT distance="225" swimtime="00:03:26.67" />
                    <SPLIT distance="250" swimtime="00:03:51.37" />
                    <SPLIT distance="275" swimtime="00:04:15.22" />
                    <SPLIT distance="300" swimtime="00:04:39.11" />
                    <SPLIT distance="325" swimtime="00:05:03.19" />
                    <SPLIT distance="350" swimtime="00:05:27.44" />
                    <SPLIT distance="375" swimtime="00:05:51.98" />
                    <SPLIT distance="400" swimtime="00:06:16.61" />
                    <SPLIT distance="425" swimtime="00:06:40.37" />
                    <SPLIT distance="450" swimtime="00:07:04.76" />
                    <SPLIT distance="475" swimtime="00:07:28.83" />
                    <SPLIT distance="500" swimtime="00:07:52.88" />
                    <SPLIT distance="525" swimtime="00:08:16.66" />
                    <SPLIT distance="550" swimtime="00:08:41.09" />
                    <SPLIT distance="575" swimtime="00:09:05.04" />
                    <SPLIT distance="600" swimtime="00:09:29.64" />
                    <SPLIT distance="625" swimtime="00:09:53.45" />
                    <SPLIT distance="650" swimtime="00:10:17.91" />
                    <SPLIT distance="675" swimtime="00:10:41.77" />
                    <SPLIT distance="700" swimtime="00:11:05.79" />
                    <SPLIT distance="725" swimtime="00:11:29.61" />
                    <SPLIT distance="750" swimtime="00:11:54.60" />
                    <SPLIT distance="775" swimtime="00:12:18.71" />
                    <SPLIT distance="800" swimtime="00:12:43.00" />
                    <SPLIT distance="825" swimtime="00:13:06.66" />
                    <SPLIT distance="850" swimtime="00:13:31.00" />
                    <SPLIT distance="875" swimtime="00:13:55.13" />
                    <SPLIT distance="900" swimtime="00:14:19.35" />
                    <SPLIT distance="925" swimtime="00:14:44.21" />
                    <SPLIT distance="950" swimtime="00:15:09.44" />
                    <SPLIT distance="975" swimtime="00:15:33.62" />
                    <SPLIT distance="1000" swimtime="00:15:58.65" />
                    <SPLIT distance="1025" swimtime="00:16:23.18" />
                    <SPLIT distance="1050" swimtime="00:16:48.10" />
                    <SPLIT distance="1075" swimtime="00:17:12.95" />
                    <SPLIT distance="1100" swimtime="00:17:38.11" />
                    <SPLIT distance="1125" swimtime="00:18:03.18" />
                    <SPLIT distance="1150" swimtime="00:18:28.04" />
                    <SPLIT distance="1175" swimtime="00:18:53.92" />
                    <SPLIT distance="1200" swimtime="00:19:19.69" />
                    <SPLIT distance="1225" swimtime="00:19:45.29" />
                    <SPLIT distance="1250" swimtime="00:20:10.25" />
                    <SPLIT distance="1275" swimtime="00:20:34.91" />
                    <SPLIT distance="1300" swimtime="00:20:59.74" />
                    <SPLIT distance="1325" swimtime="00:21:24.85" />
                    <SPLIT distance="1350" swimtime="00:21:49.30" />
                    <SPLIT distance="1375" swimtime="00:22:14.19" />
                    <SPLIT distance="1400" swimtime="00:22:38.15" />
                    <SPLIT distance="1425" swimtime="00:23:02.77" />
                    <SPLIT distance="1450" swimtime="00:23:26.24" />
                    <SPLIT distance="1475" swimtime="00:23:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="107098" heatid="110711" lane="7" entrytime="00:03:30.00" />
                <RESULT eventid="99218" points="223" swimtime="00:02:43.71" resultid="107099" heatid="110772" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.81" />
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="75" swimtime="00:00:58.16" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                    <SPLIT distance="125" swimtime="00:01:39.98" />
                    <SPLIT distance="150" swimtime="00:02:01.05" />
                    <SPLIT distance="175" swimtime="00:02:22.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="144" reactiontime="+102" swimtime="00:01:32.23" resultid="107100" heatid="110799" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.84" />
                    <SPLIT distance="50" swimtime="00:00:44.07" />
                    <SPLIT distance="75" swimtime="00:01:07.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="215" reactiontime="+102" swimtime="00:05:54.07" resultid="107101" heatid="110849" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.07" />
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="75" swimtime="00:01:01.75" />
                    <SPLIT distance="100" swimtime="00:01:23.81" />
                    <SPLIT distance="125" swimtime="00:01:46.02" />
                    <SPLIT distance="150" swimtime="00:02:08.41" />
                    <SPLIT distance="175" swimtime="00:02:31.38" />
                    <SPLIT distance="200" swimtime="00:02:53.89" />
                    <SPLIT distance="225" swimtime="00:03:16.13" />
                    <SPLIT distance="250" swimtime="00:03:38.30" />
                    <SPLIT distance="275" swimtime="00:04:01.05" />
                    <SPLIT distance="300" swimtime="00:04:23.70" />
                    <SPLIT distance="325" swimtime="00:04:46.61" />
                    <SPLIT distance="350" swimtime="00:05:09.91" />
                    <SPLIT distance="375" swimtime="00:05:32.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="107088">
              <RESULTS>
                <RESULT eventid="98814" points="294" reactiontime="+88" swimtime="00:03:03.11" resultid="107089" heatid="110617" lane="1" entrytime="00:02:58.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.08" />
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="75" swimtime="00:01:03.24" />
                    <SPLIT distance="100" swimtime="00:01:25.59" />
                    <SPLIT distance="125" swimtime="00:01:52.05" />
                    <SPLIT distance="150" swimtime="00:02:18.49" />
                    <SPLIT distance="175" swimtime="00:02:41.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106254" points="296" reactiontime="+104" swimtime="00:22:58.53" resultid="107090" heatid="110640" lane="2" entrytime="00:23:43.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.17" />
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="75" swimtime="00:01:03.34" />
                    <SPLIT distance="100" swimtime="00:01:25.48" />
                    <SPLIT distance="125" swimtime="00:01:47.99" />
                    <SPLIT distance="150" swimtime="00:02:10.66" />
                    <SPLIT distance="175" swimtime="00:02:33.53" />
                    <SPLIT distance="200" swimtime="00:02:56.54" />
                    <SPLIT distance="225" swimtime="00:03:19.57" />
                    <SPLIT distance="250" swimtime="00:03:42.74" />
                    <SPLIT distance="275" swimtime="00:04:05.54" />
                    <SPLIT distance="300" swimtime="00:04:28.42" />
                    <SPLIT distance="325" swimtime="00:04:51.57" />
                    <SPLIT distance="350" swimtime="00:05:14.79" />
                    <SPLIT distance="375" swimtime="00:05:37.91" />
                    <SPLIT distance="400" swimtime="00:06:00.83" />
                    <SPLIT distance="425" swimtime="00:06:23.61" />
                    <SPLIT distance="450" swimtime="00:06:46.31" />
                    <SPLIT distance="475" swimtime="00:07:09.62" />
                    <SPLIT distance="500" swimtime="00:07:32.79" />
                    <SPLIT distance="525" swimtime="00:07:56.02" />
                    <SPLIT distance="550" swimtime="00:08:19.24" />
                    <SPLIT distance="575" swimtime="00:08:42.46" />
                    <SPLIT distance="600" swimtime="00:09:05.54" />
                    <SPLIT distance="625" swimtime="00:09:28.88" />
                    <SPLIT distance="650" swimtime="00:09:51.88" />
                    <SPLIT distance="675" swimtime="00:10:14.98" />
                    <SPLIT distance="700" swimtime="00:10:38.32" />
                    <SPLIT distance="725" swimtime="00:11:01.51" />
                    <SPLIT distance="750" swimtime="00:11:24.83" />
                    <SPLIT distance="775" swimtime="00:11:48.23" />
                    <SPLIT distance="800" swimtime="00:12:11.30" />
                    <SPLIT distance="825" swimtime="00:12:34.47" />
                    <SPLIT distance="850" swimtime="00:12:57.80" />
                    <SPLIT distance="875" swimtime="00:13:20.95" />
                    <SPLIT distance="900" swimtime="00:13:44.51" />
                    <SPLIT distance="925" swimtime="00:14:07.31" />
                    <SPLIT distance="950" swimtime="00:14:30.80" />
                    <SPLIT distance="975" swimtime="00:14:53.83" />
                    <SPLIT distance="1000" swimtime="00:15:17.31" />
                    <SPLIT distance="1025" swimtime="00:15:40.02" />
                    <SPLIT distance="1050" swimtime="00:16:03.34" />
                    <SPLIT distance="1075" swimtime="00:16:26.70" />
                    <SPLIT distance="1100" swimtime="00:16:49.77" />
                    <SPLIT distance="1125" swimtime="00:17:13.03" />
                    <SPLIT distance="1150" swimtime="00:17:36.11" />
                    <SPLIT distance="1175" swimtime="00:17:59.20" />
                    <SPLIT distance="1200" swimtime="00:18:22.97" />
                    <SPLIT distance="1225" swimtime="00:18:46.37" />
                    <SPLIT distance="1250" swimtime="00:19:09.20" />
                    <SPLIT distance="1275" swimtime="00:19:32.31" />
                    <SPLIT distance="1300" swimtime="00:19:56.09" />
                    <SPLIT distance="1325" swimtime="00:20:19.00" />
                    <SPLIT distance="1350" swimtime="00:20:42.05" />
                    <SPLIT distance="1375" swimtime="00:21:05.24" />
                    <SPLIT distance="1400" swimtime="00:21:28.81" />
                    <SPLIT distance="1425" swimtime="00:21:51.78" />
                    <SPLIT distance="1450" swimtime="00:22:14.69" />
                    <SPLIT distance="1475" swimtime="00:22:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="248" reactiontime="+90" swimtime="00:01:27.50" resultid="107091" heatid="110756" lane="9" entrytime="00:01:23.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.31" />
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="75" swimtime="00:01:04.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="295" reactiontime="+97" swimtime="00:06:29.52" resultid="107092" heatid="110787" lane="8" entrytime="00:06:25.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.84" />
                    <SPLIT distance="50" swimtime="00:00:42.51" />
                    <SPLIT distance="75" swimtime="00:01:08.60" />
                    <SPLIT distance="100" swimtime="00:01:34.32" />
                    <SPLIT distance="125" swimtime="00:01:59.22" />
                    <SPLIT distance="150" swimtime="00:02:23.15" />
                    <SPLIT distance="175" swimtime="00:02:47.19" />
                    <SPLIT distance="200" swimtime="00:03:11.04" />
                    <SPLIT distance="225" swimtime="00:03:38.18" />
                    <SPLIT distance="250" swimtime="00:04:05.30" />
                    <SPLIT distance="275" swimtime="00:04:32.36" />
                    <SPLIT distance="300" swimtime="00:05:00.19" />
                    <SPLIT distance="325" swimtime="00:05:23.13" />
                    <SPLIT distance="350" swimtime="00:05:45.54" />
                    <SPLIT distance="375" swimtime="00:06:08.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="262" reactiontime="+102" swimtime="00:03:06.21" resultid="107093" heatid="110809" lane="1" entrytime="00:02:58.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.27" />
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="75" swimtime="00:01:06.86" />
                    <SPLIT distance="100" swimtime="00:01:30.81" />
                    <SPLIT distance="125" swimtime="00:01:54.50" />
                    <SPLIT distance="150" swimtime="00:02:18.93" />
                    <SPLIT distance="175" swimtime="00:02:43.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="269" swimtime="00:06:03.00" resultid="107094" heatid="110840" lane="0" entrytime="00:05:50.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.54" />
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="75" swimtime="00:01:01.96" />
                    <SPLIT distance="100" swimtime="00:01:24.38" />
                    <SPLIT distance="125" swimtime="00:01:46.63" />
                    <SPLIT distance="150" swimtime="00:02:09.43" />
                    <SPLIT distance="175" swimtime="00:02:31.80" />
                    <SPLIT distance="200" swimtime="00:02:55.34" />
                    <SPLIT distance="225" swimtime="00:03:18.94" />
                    <SPLIT distance="250" swimtime="00:03:42.26" />
                    <SPLIT distance="275" swimtime="00:04:06.00" />
                    <SPLIT distance="300" swimtime="00:04:29.58" />
                    <SPLIT distance="325" swimtime="00:04:53.18" />
                    <SPLIT distance="350" swimtime="00:05:17.06" />
                    <SPLIT distance="375" swimtime="00:05:40.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WA" clubid="106570" name="Swimmers St. Pływackie">
          <CONTACT city="WARSZAWA" email="remog@swimmersteam.pl" name="GOŁĘBIOWSKI REMO" phone="601333 782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1978-08-12" firstname="Jan" gender="M" lastname="Rekowski" nation="POL" athleteid="106578">
              <RESULTS>
                <RESULT eventid="98798" points="481" reactiontime="+77" swimtime="00:00:25.84" resultid="106579" heatid="110611" lane="8" entrytime="00:00:25.85">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="469" reactiontime="+84" swimtime="00:00:57.81" resultid="106580" heatid="110686" lane="3" entrytime="00:01:01.09">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.38" />
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="75" swimtime="00:00:42.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="355" reactiontime="+99" swimtime="00:01:11.50" resultid="106581" heatid="110702" lane="1" entrytime="00:01:12.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.10" />
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="75" swimtime="00:00:54.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="401" swimtime="00:00:29.56" resultid="106582" heatid="110749" lane="0" entrytime="00:00:29.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="106583" heatid="110774" lane="2" entrytime="00:02:26.25" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="106584" heatid="110831" lane="7" entrytime="00:00:35.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-11-27" firstname="Sopolińska" gender="F" lastname="Emilia" nation="POL" athleteid="106591">
              <RESULTS>
                <RESULT eventid="98777" points="230" swimtime="00:00:37.92" resultid="106592" heatid="110589" lane="9" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="157" reactiontime="+99" swimtime="00:03:45.45" resultid="106593" heatid="110615" lane="8" entrytime="00:03:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.37" />
                    <SPLIT distance="50" swimtime="00:00:53.24" />
                    <SPLIT distance="75" swimtime="00:01:25.45" />
                    <SPLIT distance="100" swimtime="00:01:54.36" />
                    <SPLIT distance="125" swimtime="00:02:24.99" />
                    <SPLIT distance="150" swimtime="00:02:56.51" />
                    <SPLIT distance="175" swimtime="00:03:21.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="210" reactiontime="+115" swimtime="00:01:25.64" resultid="106594" heatid="110673" lane="1" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.88" />
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="75" swimtime="00:01:03.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="171" reactiontime="+95" swimtime="00:01:42.09" resultid="106595" heatid="110691" lane="5" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.41" />
                    <SPLIT distance="50" swimtime="00:00:51.40" />
                    <SPLIT distance="75" swimtime="00:01:20.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="106596" heatid="110765" lane="3" entrytime="00:03:11.00" />
                <RESULT eventid="99266" points="151" swimtime="00:08:06.31" resultid="106597" heatid="110786" lane="0" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.29" />
                    <SPLIT distance="50" swimtime="00:00:58.28" />
                    <SPLIT distance="75" swimtime="00:01:30.46" />
                    <SPLIT distance="100" swimtime="00:02:04.70" />
                    <SPLIT distance="125" swimtime="00:02:38.67" />
                    <SPLIT distance="150" swimtime="00:03:11.89" />
                    <SPLIT distance="175" swimtime="00:03:44.79" />
                    <SPLIT distance="200" swimtime="00:04:18.29" />
                    <SPLIT distance="225" swimtime="00:04:48.60" />
                    <SPLIT distance="250" swimtime="00:05:21.67" />
                    <SPLIT distance="275" swimtime="00:05:51.42" />
                    <SPLIT distance="300" swimtime="00:06:23.32" />
                    <SPLIT distance="325" swimtime="00:06:48.91" />
                    <SPLIT distance="350" swimtime="00:07:15.57" />
                    <SPLIT distance="375" swimtime="00:07:41.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="205" swimtime="00:06:37.29" resultid="106598" heatid="110841" lane="9" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.09" />
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                    <SPLIT distance="75" swimtime="00:01:07.16" />
                    <SPLIT distance="100" swimtime="00:01:31.67" />
                    <SPLIT distance="125" swimtime="00:01:56.59" />
                    <SPLIT distance="150" swimtime="00:02:21.37" />
                    <SPLIT distance="175" swimtime="00:02:46.89" />
                    <SPLIT distance="200" swimtime="00:03:12.53" />
                    <SPLIT distance="225" swimtime="00:03:38.82" />
                    <SPLIT distance="250" swimtime="00:04:04.62" />
                    <SPLIT distance="275" swimtime="00:04:30.65" />
                    <SPLIT distance="300" swimtime="00:04:56.12" />
                    <SPLIT distance="325" swimtime="00:05:21.73" />
                    <SPLIT distance="350" swimtime="00:05:47.36" />
                    <SPLIT distance="375" swimtime="00:06:13.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brożyna" nation="POL" athleteid="106599">
              <RESULTS>
                <RESULT eventid="98924" points="283" reactiontime="+81" swimtime="00:00:33.83" resultid="106600" heatid="110657" lane="2" entrytime="00:00:33.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="325" reactiontime="+78" swimtime="00:01:13.67" resultid="106601" heatid="110702" lane="8" entrytime="00:01:13.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.79" />
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="75" swimtime="00:00:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="307" reactiontime="+74" swimtime="00:01:12.48" resultid="106602" heatid="110761" lane="4" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.63" />
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="75" swimtime="00:00:54.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="298" reactiontime="+95" swimtime="00:02:38.09" resultid="106603" heatid="110815" lane="9" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.45" />
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="75" swimtime="00:00:57.02" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="125" swimtime="00:01:37.44" />
                    <SPLIT distance="150" swimtime="00:01:57.64" />
                    <SPLIT distance="175" swimtime="00:02:18.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-04" firstname="Norbert" gender="M" lastname="Tchorzewski" nation="POL" athleteid="106609">
              <RESULTS>
                <RESULT eventid="98830" points="229" reactiontime="+89" swimtime="00:02:58.98" resultid="106610" heatid="110622" lane="5" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.17" />
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="75" swimtime="00:01:00.07" />
                    <SPLIT distance="100" swimtime="00:01:23.51" />
                    <SPLIT distance="125" swimtime="00:01:51.35" />
                    <SPLIT distance="150" swimtime="00:02:18.62" />
                    <SPLIT distance="175" swimtime="00:02:39.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="222" reactiontime="+107" swimtime="00:23:19.79" resultid="106611" heatid="110642" lane="7" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.74" />
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                    <SPLIT distance="75" swimtime="00:00:59.27" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="125" swimtime="00:01:42.51" />
                    <SPLIT distance="150" swimtime="00:02:03.82" />
                    <SPLIT distance="175" swimtime="00:02:25.32" />
                    <SPLIT distance="200" swimtime="00:02:47.17" />
                    <SPLIT distance="225" swimtime="00:03:09.06" />
                    <SPLIT distance="250" swimtime="00:03:31.37" />
                    <SPLIT distance="275" swimtime="00:03:53.89" />
                    <SPLIT distance="300" swimtime="00:04:16.83" />
                    <SPLIT distance="325" swimtime="00:04:39.70" />
                    <SPLIT distance="350" swimtime="00:05:03.07" />
                    <SPLIT distance="375" swimtime="00:05:26.16" />
                    <SPLIT distance="400" swimtime="00:05:49.17" />
                    <SPLIT distance="425" swimtime="00:06:11.96" />
                    <SPLIT distance="450" swimtime="00:06:34.84" />
                    <SPLIT distance="475" swimtime="00:06:58.21" />
                    <SPLIT distance="500" swimtime="00:07:21.66" />
                    <SPLIT distance="525" swimtime="00:07:45.15" />
                    <SPLIT distance="550" swimtime="00:08:08.48" />
                    <SPLIT distance="575" swimtime="00:08:32.81" />
                    <SPLIT distance="600" swimtime="00:08:56.65" />
                    <SPLIT distance="625" swimtime="00:09:20.53" />
                    <SPLIT distance="650" swimtime="00:09:44.54" />
                    <SPLIT distance="675" swimtime="00:10:08.56" />
                    <SPLIT distance="700" swimtime="00:10:31.85" />
                    <SPLIT distance="725" swimtime="00:10:54.78" />
                    <SPLIT distance="750" swimtime="00:11:17.67" />
                    <SPLIT distance="775" swimtime="00:11:42.19" />
                    <SPLIT distance="800" swimtime="00:12:05.02" />
                    <SPLIT distance="825" swimtime="00:12:27.85" />
                    <SPLIT distance="850" swimtime="00:12:51.27" />
                    <SPLIT distance="875" swimtime="00:13:14.49" />
                    <SPLIT distance="900" swimtime="00:13:38.69" />
                    <SPLIT distance="925" swimtime="00:14:03.04" />
                    <SPLIT distance="950" swimtime="00:14:27.16" />
                    <SPLIT distance="975" swimtime="00:14:51.41" />
                    <SPLIT distance="1000" swimtime="00:15:15.35" />
                    <SPLIT distance="1025" swimtime="00:15:38.91" />
                    <SPLIT distance="1050" swimtime="00:16:02.75" />
                    <SPLIT distance="1075" swimtime="00:16:27.47" />
                    <SPLIT distance="1100" swimtime="00:16:51.47" />
                    <SPLIT distance="1125" swimtime="00:17:15.76" />
                    <SPLIT distance="1150" swimtime="00:17:39.86" />
                    <SPLIT distance="1175" swimtime="00:18:03.49" />
                    <SPLIT distance="1200" swimtime="00:18:27.25" />
                    <SPLIT distance="1225" swimtime="00:18:51.14" />
                    <SPLIT distance="1250" swimtime="00:19:15.22" />
                    <SPLIT distance="1275" swimtime="00:19:39.57" />
                    <SPLIT distance="1300" swimtime="00:20:03.43" />
                    <SPLIT distance="1325" swimtime="00:20:27.45" />
                    <SPLIT distance="1350" swimtime="00:20:51.77" />
                    <SPLIT distance="1375" swimtime="00:21:16.34" />
                    <SPLIT distance="1400" swimtime="00:21:40.43" />
                    <SPLIT distance="1425" swimtime="00:22:05.55" />
                    <SPLIT distance="1450" swimtime="00:22:30.27" />
                    <SPLIT distance="1475" swimtime="00:22:54.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="308" reactiontime="+87" swimtime="00:01:06.52" resultid="106612" heatid="110683" lane="7" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.25" />
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="75" swimtime="00:00:49.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="161" reactiontime="+96" swimtime="00:03:19.45" resultid="106613" heatid="110711" lane="6" entrytime="00:03:19.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.20" />
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="75" swimtime="00:01:04.78" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="125" swimtime="00:01:56.48" />
                    <SPLIT distance="150" swimtime="00:02:23.51" />
                    <SPLIT distance="175" swimtime="00:02:50.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="275" reactiontime="+87" swimtime="00:02:32.74" resultid="106614" heatid="110773" lane="6" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.08" />
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="75" swimtime="00:00:52.27" />
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                    <SPLIT distance="125" swimtime="00:01:31.97" />
                    <SPLIT distance="150" swimtime="00:01:52.91" />
                    <SPLIT distance="175" swimtime="00:02:13.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="106615" heatid="110789" lane="7" entrytime="00:06:59.00" />
                <RESULT eventid="99361" points="197" swimtime="00:01:23.14" resultid="106616" heatid="110801" lane="9" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.26" />
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="75" swimtime="00:01:01.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="246" swimtime="00:05:38.49" resultid="106617" heatid="110847" lane="0" entrytime="00:05:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.88" />
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                    <SPLIT distance="75" swimtime="00:00:58.47" />
                    <SPLIT distance="100" swimtime="00:01:19.69" />
                    <SPLIT distance="125" swimtime="00:01:41.54" />
                    <SPLIT distance="150" swimtime="00:02:03.55" />
                    <SPLIT distance="175" swimtime="00:02:26.34" />
                    <SPLIT distance="200" swimtime="00:02:48.97" />
                    <SPLIT distance="225" swimtime="00:03:10.83" />
                    <SPLIT distance="250" swimtime="00:03:33.03" />
                    <SPLIT distance="275" swimtime="00:03:54.98" />
                    <SPLIT distance="300" swimtime="00:04:17.04" />
                    <SPLIT distance="325" swimtime="00:04:38.84" />
                    <SPLIT distance="350" swimtime="00:05:00.39" />
                    <SPLIT distance="375" swimtime="00:05:21.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-07-31" firstname="Katarzyna" gender="F" lastname="Herczyńska" nation="POL" athleteid="106618">
              <RESULTS>
                <RESULT eventid="99154" points="280" reactiontime="+94" swimtime="00:00:37.23" resultid="106619" heatid="110737" lane="1" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-27" firstname="Remigiusz" gender="M" lastname="Miklewski" nation="POL" athleteid="106604">
              <RESULTS>
                <RESULT eventid="98798" points="336" reactiontime="+74" swimtime="00:00:29.14" resultid="106605" heatid="110604" lane="0" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="268" swimtime="00:01:09.62" resultid="106606" heatid="110682" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.97" />
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="75" swimtime="00:00:50.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="186" reactiontime="+49" swimtime="00:02:53.96" resultid="106607" heatid="110771" lane="2" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.23" />
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="75" swimtime="00:01:00.34" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="125" swimtime="00:01:45.75" />
                    <SPLIT distance="150" swimtime="00:02:09.06" />
                    <SPLIT distance="175" swimtime="00:02:32.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="106608" heatid="110828" lane="7" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Bolesław" gender="M" lastname="Porolniczak" nation="POL" athleteid="109147">
              <RESULTS>
                <RESULT eventid="98798" points="439" reactiontime="+95" swimtime="00:00:26.65" resultid="109148" heatid="110608" lane="1" entrytime="00:00:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="435" reactiontime="+93" swimtime="00:00:59.30" resultid="109149" heatid="110685" lane="2" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                    <SPLIT distance="75" swimtime="00:00:43.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="379" reactiontime="+58" swimtime="00:01:09.99" resultid="109150" heatid="110701" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.33" />
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="75" swimtime="00:00:54.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="109151" heatid="110746" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="99218" points="400" reactiontime="+90" swimtime="00:02:14.77" resultid="110210" heatid="110776" lane="8" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.66" />
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="75" swimtime="00:00:46.94" />
                    <SPLIT distance="100" swimtime="00:01:04.10" />
                    <SPLIT distance="125" swimtime="00:01:21.71" />
                    <SPLIT distance="150" swimtime="00:01:39.57" />
                    <SPLIT distance="175" swimtime="00:01:57.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-01" firstname="Katarzyna" gender="F" lastname="Koba-Gołaszewska" nation="POL" athleteid="106585">
              <RESULTS>
                <RESULT eventid="98777" points="404" reactiontime="+79" swimtime="00:00:31.43" resultid="106586" heatid="110591" lane="4" entrytime="00:00:30.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="391" reactiontime="+83" swimtime="00:01:09.60" resultid="106587" heatid="110675" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.59" />
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="75" swimtime="00:00:51.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="369" reactiontime="+86" swimtime="00:00:33.96" resultid="106588" heatid="110739" lane="1" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="321" reactiontime="+74" swimtime="00:02:41.71" resultid="106589" heatid="110767" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.49" />
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="75" swimtime="00:00:54.74" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="125" swimtime="00:01:36.58" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                    <SPLIT distance="175" swimtime="00:02:20.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="263" swimtime="00:01:25.17" resultid="106590" heatid="110795" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.48" />
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="75" swimtime="00:01:02.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-07-07" firstname="Remigiusz" gender="M" lastname="Gołębiowski" nation="POL" athleteid="106571">
              <RESULTS>
                <RESULT eventid="98798" points="443" reactiontime="+77" swimtime="00:00:26.56" resultid="106572" heatid="110609" lane="1" entrytime="00:00:26.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="421" reactiontime="+63" swimtime="00:09:51.27" resultid="106573" heatid="110635" lane="5" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.97" />
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="75" swimtime="00:00:49.76" />
                    <SPLIT distance="100" swimtime="00:01:07.65" />
                    <SPLIT distance="125" swimtime="00:01:25.96" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                    <SPLIT distance="175" swimtime="00:02:02.79" />
                    <SPLIT distance="200" swimtime="00:02:21.40" />
                    <SPLIT distance="225" swimtime="00:02:39.79" />
                    <SPLIT distance="250" swimtime="00:02:58.33" />
                    <SPLIT distance="275" swimtime="00:03:16.64" />
                    <SPLIT distance="300" swimtime="00:03:35.31" />
                    <SPLIT distance="325" swimtime="00:03:53.85" />
                    <SPLIT distance="350" swimtime="00:04:12.22" />
                    <SPLIT distance="375" swimtime="00:04:30.55" />
                    <SPLIT distance="400" swimtime="00:04:49.35" />
                    <SPLIT distance="425" swimtime="00:05:07.43" />
                    <SPLIT distance="450" swimtime="00:05:26.32" />
                    <SPLIT distance="475" swimtime="00:05:45.00" />
                    <SPLIT distance="500" swimtime="00:06:03.96" />
                    <SPLIT distance="525" swimtime="00:06:22.61" />
                    <SPLIT distance="550" swimtime="00:06:41.72" />
                    <SPLIT distance="575" swimtime="00:07:00.29" />
                    <SPLIT distance="600" swimtime="00:07:19.19" />
                    <SPLIT distance="625" swimtime="00:07:38.13" />
                    <SPLIT distance="650" swimtime="00:07:57.16" />
                    <SPLIT distance="675" swimtime="00:08:16.37" />
                    <SPLIT distance="700" swimtime="00:08:35.31" />
                    <SPLIT distance="725" swimtime="00:08:54.15" />
                    <SPLIT distance="750" swimtime="00:09:13.41" />
                    <SPLIT distance="775" swimtime="00:09:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="484" reactiontime="+74" swimtime="00:00:27.75" resultid="106574" heatid="110750" lane="4" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="425" reactiontime="+72" swimtime="00:02:12.13" resultid="106575" heatid="110777" lane="4" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.18" />
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="75" swimtime="00:00:46.53" />
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                    <SPLIT distance="125" swimtime="00:01:20.18" />
                    <SPLIT distance="150" swimtime="00:01:37.40" />
                    <SPLIT distance="175" swimtime="00:01:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="106576" heatid="110804" lane="6" entrytime="00:01:05.00" />
                <RESULT eventid="99473" points="378" reactiontime="+83" swimtime="00:04:53.40" resultid="106577" heatid="110844" lane="4" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.60" />
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="75" swimtime="00:00:50.97" />
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                    <SPLIT distance="125" swimtime="00:01:28.04" />
                    <SPLIT distance="150" swimtime="00:01:46.84" />
                    <SPLIT distance="175" swimtime="00:02:05.79" />
                    <SPLIT distance="200" swimtime="00:02:24.61" />
                    <SPLIT distance="225" swimtime="00:02:43.24" />
                    <SPLIT distance="250" swimtime="00:03:02.45" />
                    <SPLIT distance="275" swimtime="00:03:21.14" />
                    <SPLIT distance="300" swimtime="00:03:40.02" />
                    <SPLIT distance="325" swimtime="00:03:58.63" />
                    <SPLIT distance="350" swimtime="00:04:17.10" />
                    <SPLIT distance="375" swimtime="00:04:36.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="395" reactiontime="+73" swimtime="00:02:03.34" resultid="106622" heatid="110718" lane="1" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.07" />
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="75" swimtime="00:00:50.21" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="125" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:01:36.62" />
                    <SPLIT distance="175" swimtime="00:01:49.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106599" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="106578" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="106571" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="109147" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="451" reactiontime="+73" swimtime="00:01:47.64" resultid="106623" heatid="110783" lane="7" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                    <SPLIT distance="75" swimtime="00:00:40.81" />
                    <SPLIT distance="100" swimtime="00:00:55.96" />
                    <SPLIT distance="125" swimtime="00:01:08.39" />
                    <SPLIT distance="150" swimtime="00:01:21.88" />
                    <SPLIT distance="175" swimtime="00:01:34.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106571" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="106609" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="106604" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="106578" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="328" reactiontime="+82" swimtime="00:01:59.66" resultid="106620" heatid="110631" lane="8" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.85" />
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="75" swimtime="00:00:42.53" />
                    <SPLIT distance="100" swimtime="00:00:56.00" />
                    <SPLIT distance="125" swimtime="00:01:14.11" />
                    <SPLIT distance="150" swimtime="00:01:22.93" />
                    <SPLIT distance="175" swimtime="00:01:46.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106585" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="106578" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="106571" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="106591" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="260" reactiontime="+81" swimtime="00:02:21.78" resultid="106621" heatid="110837" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="75" swimtime="00:00:48.96" />
                    <SPLIT distance="100" swimtime="00:01:07.10" />
                    <SPLIT distance="125" swimtime="00:01:24.24" />
                    <SPLIT distance="150" swimtime="00:01:44.62" />
                    <SPLIT distance="175" swimtime="00:02:02.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106591" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="106599" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="106618" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="106578" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="108604" name="Swimming Masters Team Szczecin">
          <CONTACT city="Szczecin" email="aga.krzyzostaniak@gmail.com" name="Krzyżostaniak Agnieszka" phone="603772862" street="Żupańskiego 12/8" zip="71-440" />
          <ATHLETES>
            <ATHLETE birthdate="1996-02-15" firstname="Filip" gender="M" lastname="Przybyłowki" nation="POL" athleteid="108701">
              <RESULTS>
                <RESULT eventid="98798" points="427" reactiontime="+70" swimtime="00:00:26.89" resultid="108702" heatid="110605" lane="5" entrytime="00:00:28.74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="426" reactiontime="+66" swimtime="00:00:59.71" resultid="108703" heatid="110684" lane="5" entrytime="00:01:03.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.17" />
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                    <SPLIT distance="75" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="396" swimtime="00:00:29.68" resultid="108704" heatid="110746" lane="6" entrytime="00:00:31.64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="374" reactiontime="+80" swimtime="00:02:17.87" resultid="108705" heatid="110773" lane="1" entrytime="00:02:34.53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.30" />
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="75" swimtime="00:00:48.06" />
                    <SPLIT distance="100" swimtime="00:01:06.03" />
                    <SPLIT distance="125" swimtime="00:01:24.08" />
                    <SPLIT distance="150" swimtime="00:01:42.29" />
                    <SPLIT distance="175" swimtime="00:02:00.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="378" reactiontime="+68" swimtime="00:01:06.95" resultid="108706" heatid="110802" lane="5" entrytime="00:01:10.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.10" />
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="75" swimtime="00:00:48.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-14" firstname="Kinga" gender="F" lastname="Maciupa" nation="POL" athleteid="108671">
              <RESULTS>
                <RESULT eventid="98777" points="482" reactiontime="+74" swimtime="00:00:29.64" resultid="108672" heatid="110592" lane="8" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="469" reactiontime="+78" swimtime="00:02:36.75" resultid="108673" heatid="110618" lane="8" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.87" />
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="75" swimtime="00:00:53.64" />
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="125" swimtime="00:01:35.88" />
                    <SPLIT distance="150" swimtime="00:01:58.66" />
                    <SPLIT distance="175" swimtime="00:02:18.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="511" reactiontime="+74" swimtime="00:00:32.10" resultid="108674" heatid="110650" lane="1" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="506" reactiontime="+90" swimtime="00:01:11.09" resultid="108675" heatid="110695" lane="1" entrytime="00:01:13.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.62" />
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="75" swimtime="00:00:53.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="516" reactiontime="+65" swimtime="00:01:08.57" resultid="108676" heatid="110756" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.26" />
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="75" swimtime="00:00:51.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="485" reactiontime="+43" swimtime="00:05:30.06" resultid="108677" heatid="110787" lane="4" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.83" />
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="75" swimtime="00:00:51.48" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="125" swimtime="00:01:33.85" />
                    <SPLIT distance="150" swimtime="00:01:54.95" />
                    <SPLIT distance="175" swimtime="00:02:16.14" />
                    <SPLIT distance="200" swimtime="00:02:37.20" />
                    <SPLIT distance="225" swimtime="00:03:00.90" />
                    <SPLIT distance="250" swimtime="00:03:24.88" />
                    <SPLIT distance="275" swimtime="00:03:48.56" />
                    <SPLIT distance="300" swimtime="00:04:12.36" />
                    <SPLIT distance="325" swimtime="00:04:32.61" />
                    <SPLIT distance="350" swimtime="00:04:52.24" />
                    <SPLIT distance="375" swimtime="00:05:11.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="466" swimtime="00:01:10.41" resultid="108678" heatid="110796" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.63" />
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="75" swimtime="00:00:50.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-07" firstname="Marta" gender="F" lastname="Pachuc" nation="POL" athleteid="108666">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="108667" heatid="110590" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="108668" heatid="110675" lane="1" entrytime="00:01:12.00" />
                <RESULT eventid="99089" status="DNS" swimtime="00:00:00.00" resultid="108669" heatid="110723" lane="8" entrytime="00:01:40.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="108670" heatid="110820" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="Roenig" nation="POL" athleteid="108628">
              <RESULTS>
                <RESULT eventid="98798" points="429" reactiontime="+79" swimtime="00:00:26.86" resultid="108629" heatid="110607" lane="6" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="403" reactiontime="+86" swimtime="00:01:00.81" resultid="108630" heatid="110685" lane="6" entrytime="00:01:02.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                    <SPLIT distance="75" swimtime="00:00:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="345" swimtime="00:01:19.26" resultid="108631" heatid="110729" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.01" />
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="75" swimtime="00:00:59.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="355" swimtime="00:00:30.76" resultid="108632" heatid="110747" lane="0" entrytime="00:00:31.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="108633" heatid="110800" lane="1" entrytime="00:01:30.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="108634" heatid="110831" lane="2" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-02-07" firstname="Szymon" gender="M" lastname="Klimkowski" nation="POL" athleteid="108688">
              <RESULTS>
                <RESULT eventid="98798" points="386" reactiontime="+77" swimtime="00:00:27.82" resultid="108689" heatid="110607" lane="8" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="341" reactiontime="+85" swimtime="00:02:36.86" resultid="108690" heatid="110624" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.70" />
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="75" swimtime="00:00:53.36" />
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                    <SPLIT distance="125" swimtime="00:01:37.05" />
                    <SPLIT distance="150" swimtime="00:02:01.44" />
                    <SPLIT distance="175" swimtime="00:02:20.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="280" reactiontime="+78" swimtime="00:00:33.95" resultid="108691" heatid="110657" lane="9" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="348" reactiontime="+81" swimtime="00:01:11.97" resultid="108692" heatid="110700" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="75" swimtime="00:00:55.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="382" swimtime="00:00:30.04" resultid="108693" heatid="110748" lane="3" entrytime="00:00:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="260" reactiontime="+78" swimtime="00:00:39.52" resultid="108694" heatid="110829" lane="1" entrytime="00:00:38.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-12" firstname="Marek" gender="M" lastname="Zienkiewicz" nation="POL" athleteid="108657">
              <RESULTS>
                <RESULT eventid="98798" points="320" reactiontime="+68" swimtime="00:00:29.59" resultid="108658" heatid="110603" lane="7" entrytime="00:00:30.35">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="217" swimtime="00:03:02.18" resultid="108659" heatid="110624" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="75" swimtime="00:01:03.46" />
                    <SPLIT distance="100" swimtime="00:01:28.78" />
                    <SPLIT distance="125" swimtime="00:01:53.34" />
                    <SPLIT distance="150" swimtime="00:02:18.48" />
                    <SPLIT distance="175" swimtime="00:02:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="282" reactiontime="+48" swimtime="00:01:08.52" resultid="108660" heatid="110682" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.35" />
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="75" swimtime="00:00:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="256" reactiontime="+85" swimtime="00:01:19.71" resultid="108661" heatid="110698" lane="3" entrytime="00:01:22.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.86" />
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                    <SPLIT distance="75" swimtime="00:01:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="289" swimtime="00:00:32.97" resultid="108662" heatid="110745" lane="9" entrytime="00:00:33.75">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="202" swimtime="00:02:49.11" resultid="108663" heatid="110774" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.08" />
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="75" swimtime="00:00:58.58" />
                    <SPLIT distance="100" swimtime="00:01:20.63" />
                    <SPLIT distance="125" swimtime="00:01:42.11" />
                    <SPLIT distance="150" swimtime="00:02:04.24" />
                    <SPLIT distance="175" swimtime="00:02:26.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="315" reactiontime="+71" swimtime="00:00:37.09" resultid="108664" heatid="110829" lane="5" entrytime="00:00:37.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="191" swimtime="00:06:07.99" resultid="108665" heatid="110849" lane="6" entrytime="00:06:09.46">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.96" />
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                    <SPLIT distance="75" swimtime="00:01:01.08" />
                    <SPLIT distance="100" swimtime="00:01:23.59" />
                    <SPLIT distance="125" swimtime="00:01:46.46" />
                    <SPLIT distance="150" swimtime="00:02:09.81" />
                    <SPLIT distance="175" swimtime="00:02:33.14" />
                    <SPLIT distance="200" swimtime="00:02:56.45" />
                    <SPLIT distance="225" swimtime="00:03:20.74" />
                    <SPLIT distance="250" swimtime="00:03:44.70" />
                    <SPLIT distance="275" swimtime="00:04:09.13" />
                    <SPLIT distance="300" swimtime="00:04:33.58" />
                    <SPLIT distance="325" swimtime="00:04:57.02" />
                    <SPLIT distance="350" swimtime="00:05:21.31" />
                    <SPLIT distance="375" swimtime="00:05:45.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-11-04" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="108707">
              <RESULTS>
                <RESULT eventid="98798" points="219" reactiontime="+105" swimtime="00:00:33.59" resultid="108708" heatid="110600" lane="7" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-10" firstname="Krzysztof" gender="M" lastname="Kwieciński" nation="POL" athleteid="108709">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="108710" heatid="110598" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="108711" heatid="110679" lane="2" entrytime="00:01:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-12" firstname="Dominika" gender="F" lastname="Zielińska" nation="POL" athleteid="108679">
              <RESULTS>
                <RESULT eventid="98814" points="354" reactiontime="+93" swimtime="00:02:52.23" resultid="108680" heatid="110617" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.29" />
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="75" swimtime="00:00:57.78" />
                    <SPLIT distance="100" swimtime="00:01:18.93" />
                    <SPLIT distance="125" swimtime="00:01:44.02" />
                    <SPLIT distance="150" swimtime="00:02:10.52" />
                    <SPLIT distance="175" swimtime="00:02:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="333" reactiontime="+105" swimtime="00:11:31.11" resultid="108681" heatid="110633" lane="3" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.74" />
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="75" swimtime="00:00:57.43" />
                    <SPLIT distance="100" swimtime="00:01:18.06" />
                    <SPLIT distance="125" swimtime="00:01:38.69" />
                    <SPLIT distance="150" swimtime="00:01:59.53" />
                    <SPLIT distance="175" swimtime="00:02:20.80" />
                    <SPLIT distance="200" swimtime="00:02:42.33" />
                    <SPLIT distance="225" swimtime="00:03:03.89" />
                    <SPLIT distance="250" swimtime="00:03:25.90" />
                    <SPLIT distance="275" swimtime="00:03:47.88" />
                    <SPLIT distance="300" swimtime="00:04:09.97" />
                    <SPLIT distance="325" swimtime="00:04:32.03" />
                    <SPLIT distance="350" swimtime="00:04:54.05" />
                    <SPLIT distance="375" swimtime="00:05:16.33" />
                    <SPLIT distance="400" swimtime="00:05:38.70" />
                    <SPLIT distance="425" swimtime="00:06:01.06" />
                    <SPLIT distance="450" swimtime="00:06:23.34" />
                    <SPLIT distance="475" swimtime="00:06:45.62" />
                    <SPLIT distance="500" swimtime="00:07:08.04" />
                    <SPLIT distance="525" swimtime="00:07:30.47" />
                    <SPLIT distance="550" swimtime="00:07:53.47" />
                    <SPLIT distance="575" swimtime="00:08:15.94" />
                    <SPLIT distance="600" swimtime="00:08:38.48" />
                    <SPLIT distance="625" swimtime="00:09:01.28" />
                    <SPLIT distance="650" swimtime="00:09:23.77" />
                    <SPLIT distance="675" swimtime="00:09:46.20" />
                    <SPLIT distance="700" swimtime="00:10:08.36" />
                    <SPLIT distance="725" swimtime="00:10:30.17" />
                    <SPLIT distance="750" swimtime="00:10:51.93" />
                    <SPLIT distance="775" swimtime="00:11:12.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="384" reactiontime="+114" swimtime="00:01:10.04" resultid="108682" heatid="110673" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.42" />
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="75" swimtime="00:00:51.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="363" reactiontime="+82" swimtime="00:01:19.43" resultid="108683" heatid="110693" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.74" />
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="75" swimtime="00:01:01.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="345" reactiontime="+87" swimtime="00:01:18.44" resultid="108684" heatid="110756" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                    <SPLIT distance="75" swimtime="00:00:57.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="352" reactiontime="+92" swimtime="00:02:36.89" resultid="108685" heatid="110766" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.32" />
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="75" swimtime="00:00:56.14" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="125" swimtime="00:01:37.08" />
                    <SPLIT distance="150" swimtime="00:01:57.68" />
                    <SPLIT distance="175" swimtime="00:02:18.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="313" reactiontime="+85" swimtime="00:01:20.38" resultid="108686" heatid="110795" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.08" />
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="75" swimtime="00:00:58.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="337" reactiontime="+78" swimtime="00:02:51.26" resultid="108687" heatid="110809" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.01" />
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="75" swimtime="00:01:02.68" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                    <SPLIT distance="125" swimtime="00:01:47.05" />
                    <SPLIT distance="150" swimtime="00:02:09.26" />
                    <SPLIT distance="175" swimtime="00:02:30.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="Brodacki" nation="POL" athleteid="108648">
              <RESULTS>
                <RESULT eventid="98798" points="520" reactiontime="+75" swimtime="00:00:25.19" resultid="108649" heatid="110610" lane="8" entrytime="00:00:26.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="471" reactiontime="+80" swimtime="00:02:20.88" resultid="108650" heatid="110627" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.41" />
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="75" swimtime="00:00:47.38" />
                    <SPLIT distance="100" swimtime="00:01:05.03" />
                    <SPLIT distance="125" swimtime="00:01:26.26" />
                    <SPLIT distance="150" swimtime="00:01:48.17" />
                    <SPLIT distance="175" swimtime="00:02:05.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="542" reactiontime="+86" swimtime="00:00:55.09" resultid="108651" heatid="110688" lane="1" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.44" />
                    <SPLIT distance="50" swimtime="00:00:26.22" />
                    <SPLIT distance="75" swimtime="00:00:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="509" reactiontime="+73" swimtime="00:01:03.41" resultid="108652" heatid="110705" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.93" />
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="75" swimtime="00:00:48.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="466" reactiontime="+83" swimtime="00:00:28.10" resultid="108653" heatid="110749" lane="1" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="390" swimtime="00:05:22.17" resultid="108654" heatid="110792" lane="9" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="75" swimtime="00:00:50.97" />
                    <SPLIT distance="100" swimtime="00:01:10.38" />
                    <SPLIT distance="125" swimtime="00:01:31.20" />
                    <SPLIT distance="150" swimtime="00:01:51.73" />
                    <SPLIT distance="175" swimtime="00:02:12.77" />
                    <SPLIT distance="200" swimtime="00:02:33.97" />
                    <SPLIT distance="225" swimtime="00:02:57.43" />
                    <SPLIT distance="250" swimtime="00:03:21.15" />
                    <SPLIT distance="275" swimtime="00:03:44.73" />
                    <SPLIT distance="300" swimtime="00:04:08.61" />
                    <SPLIT distance="325" swimtime="00:04:27.29" />
                    <SPLIT distance="350" swimtime="00:04:45.74" />
                    <SPLIT distance="375" swimtime="00:05:04.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="388" reactiontime="+89" swimtime="00:00:34.61" resultid="108655" heatid="110833" lane="1" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="388" swimtime="00:04:50.94" resultid="108656" heatid="110845" lane="6" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.87" />
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="75" swimtime="00:00:48.67" />
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                    <SPLIT distance="125" swimtime="00:01:24.17" />
                    <SPLIT distance="150" swimtime="00:01:42.31" />
                    <SPLIT distance="175" swimtime="00:02:00.59" />
                    <SPLIT distance="200" swimtime="00:02:19.09" />
                    <SPLIT distance="225" swimtime="00:02:38.23" />
                    <SPLIT distance="250" swimtime="00:02:57.76" />
                    <SPLIT distance="275" swimtime="00:03:16.81" />
                    <SPLIT distance="300" swimtime="00:03:36.03" />
                    <SPLIT distance="325" swimtime="00:03:55.69" />
                    <SPLIT distance="350" swimtime="00:04:14.99" />
                    <SPLIT distance="375" swimtime="00:04:33.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-29" firstname="Robert" gender="M" lastname="Szota" nation="POL" athleteid="108695">
              <RESULTS>
                <RESULT eventid="98798" points="304" reactiontime="+93" swimtime="00:00:30.12" resultid="108696" heatid="110602" lane="1" entrytime="00:00:31.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="307" reactiontime="+78" swimtime="00:01:06.59" resultid="108697" heatid="110681" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.37" />
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="75" swimtime="00:00:50.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="280" reactiontime="+77" swimtime="00:01:17.35" resultid="108698" heatid="110699" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.85" />
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="75" swimtime="00:00:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="248" reactiontime="+84" swimtime="00:00:34.68" resultid="108699" heatid="110744" lane="8" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="287" swimtime="00:00:38.25" resultid="108700" heatid="110828" lane="9" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-12" firstname="Kamila" gender="F" lastname="Gębka" nation="POL" athleteid="108643">
              <RESULTS>
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="108644" heatid="110617" lane="8" entrytime="00:03:00.00" />
                <RESULT eventid="98940" points="339" swimtime="00:03:12.84" resultid="108645" heatid="110664" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.96" />
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                    <SPLIT distance="75" swimtime="00:01:07.67" />
                    <SPLIT distance="100" swimtime="00:01:32.61" />
                    <SPLIT distance="125" swimtime="00:01:57.15" />
                    <SPLIT distance="150" swimtime="00:02:22.95" />
                    <SPLIT distance="175" swimtime="00:02:47.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="321" reactiontime="+107" swimtime="00:01:31.01" resultid="108646" heatid="110723" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.11" />
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                    <SPLIT distance="75" swimtime="00:01:07.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="333" reactiontime="+102" swimtime="00:00:41.53" resultid="108647" heatid="110821" lane="8" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-09" firstname="Helena" gender="F" lastname="Szulc" nation="POL" athleteid="108620">
              <RESULTS>
                <RESULT eventid="98777" points="360" reactiontime="+81" swimtime="00:00:32.64" resultid="108621" heatid="110590" lane="4" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="331" reactiontime="+92" swimtime="00:02:56.05" resultid="108622" heatid="110617" lane="6" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.38" />
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="75" swimtime="00:01:01.73" />
                    <SPLIT distance="100" swimtime="00:01:23.63" />
                    <SPLIT distance="125" swimtime="00:01:49.41" />
                    <SPLIT distance="150" swimtime="00:02:15.03" />
                    <SPLIT distance="175" swimtime="00:02:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="344" reactiontime="+79" swimtime="00:01:20.85" resultid="108623" heatid="110694" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.78" />
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="75" swimtime="00:01:01.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="221" reactiontime="+100" swimtime="00:03:17.82" resultid="108624" heatid="110708" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.06" />
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                    <SPLIT distance="75" swimtime="00:01:10.11" />
                    <SPLIT distance="100" swimtime="00:01:35.76" />
                    <SPLIT distance="125" swimtime="00:02:01.29" />
                    <SPLIT distance="150" swimtime="00:02:27.01" />
                    <SPLIT distance="175" swimtime="00:02:52.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="295" swimtime="00:00:36.60" resultid="108625" heatid="110739" lane="9" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="321" reactiontime="+79" swimtime="00:06:18.90" resultid="108626" heatid="110787" lane="2" entrytime="00:06:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.29" />
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                    <SPLIT distance="75" swimtime="00:01:05.61" />
                    <SPLIT distance="100" swimtime="00:01:31.10" />
                    <SPLIT distance="125" swimtime="00:01:56.23" />
                    <SPLIT distance="150" swimtime="00:02:19.50" />
                    <SPLIT distance="175" swimtime="00:02:43.02" />
                    <SPLIT distance="200" swimtime="00:03:05.84" />
                    <SPLIT distance="225" swimtime="00:03:32.37" />
                    <SPLIT distance="250" swimtime="00:03:59.39" />
                    <SPLIT distance="275" swimtime="00:04:25.98" />
                    <SPLIT distance="300" swimtime="00:04:53.00" />
                    <SPLIT distance="325" swimtime="00:05:15.40" />
                    <SPLIT distance="350" swimtime="00:05:37.50" />
                    <SPLIT distance="375" swimtime="00:05:59.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="277" swimtime="00:01:23.72" resultid="108627" heatid="110795" lane="0" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.20" />
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="75" swimtime="00:01:00.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-20" firstname="Agnieszka" gender="F" lastname="Krzyżostaniak" nation="POL" athleteid="108635">
              <RESULTS>
                <RESULT eventid="98777" points="559" swimtime="00:00:28.20" resultid="108636" heatid="110593" lane="9" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="498" reactiontime="+79" swimtime="00:02:33.68" resultid="108637" heatid="110618" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.78" />
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="75" swimtime="00:00:52.81" />
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                    <SPLIT distance="125" swimtime="00:01:35.37" />
                    <SPLIT distance="150" swimtime="00:01:58.38" />
                    <SPLIT distance="175" swimtime="00:02:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="594" reactiontime="+77" swimtime="00:00:30.53" resultid="108638" heatid="110650" lane="5" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="525" reactiontime="+81" swimtime="00:01:10.21" resultid="108639" heatid="110695" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.44" />
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="75" swimtime="00:00:53.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="544" reactiontime="+73" swimtime="00:01:07.41" resultid="108640" heatid="110756" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.93" />
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="75" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="510" reactiontime="+82" swimtime="00:02:18.59" resultid="108641" heatid="110768" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.69" />
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="75" swimtime="00:00:48.36" />
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="125" swimtime="00:01:23.60" />
                    <SPLIT distance="150" swimtime="00:01:42.24" />
                    <SPLIT distance="175" swimtime="00:02:00.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="500" reactiontime="+94" swimtime="00:04:55.36" resultid="108642" heatid="110839" lane="3" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.65" />
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="75" swimtime="00:00:51.27" />
                    <SPLIT distance="100" swimtime="00:01:09.26" />
                    <SPLIT distance="125" swimtime="00:01:27.88" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                    <SPLIT distance="175" swimtime="00:02:05.86" />
                    <SPLIT distance="200" swimtime="00:02:24.71" />
                    <SPLIT distance="225" swimtime="00:02:43.97" />
                    <SPLIT distance="250" swimtime="00:03:02.81" />
                    <SPLIT distance="275" swimtime="00:03:22.20" />
                    <SPLIT distance="300" swimtime="00:03:41.19" />
                    <SPLIT distance="325" swimtime="00:04:00.06" />
                    <SPLIT distance="350" swimtime="00:04:18.97" />
                    <SPLIT distance="375" swimtime="00:04:37.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="SMT Szczecin 1" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="354" reactiontime="+48" swimtime="00:02:07.90" resultid="108720" heatid="110718" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.19" />
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="75" swimtime="00:00:46.44" />
                    <SPLIT distance="100" swimtime="00:01:05.18" />
                    <SPLIT distance="125" swimtime="00:01:20.19" />
                    <SPLIT distance="150" swimtime="00:01:38.35" />
                    <SPLIT distance="175" swimtime="00:01:52.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108648" number="1" reactiontime="+48" />
                    <RELAYPOSITION athleteid="108628" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="108695" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="108657" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="397" swimtime="00:01:52.38" resultid="108721" heatid="110784" lane="9" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.01" />
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="75" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:00:56.75" />
                    <SPLIT distance="125" swimtime="00:01:11.32" />
                    <SPLIT distance="150" swimtime="00:01:27.39" />
                    <SPLIT distance="175" swimtime="00:01:39.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108628" number="1" />
                    <RELAYPOSITION athleteid="108657" number="2" />
                    <RELAYPOSITION athleteid="108695" number="3" />
                    <RELAYPOSITION athleteid="108648" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="96" agetotalmin="80" gender="M" name="SMT Szczecin 2" number="2">
              <RESULTS>
                <RESULT eventid="99059" status="DNS" swimtime="00:00:00.00" resultid="108722" heatid="110717" lane="2" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108688" number="1" />
                    <RELAYPOSITION athleteid="108707" number="2" />
                    <RELAYPOSITION athleteid="108701" number="3" />
                    <RELAYPOSITION athleteid="108709" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" status="DNS" swimtime="00:00:00.00" resultid="108723" heatid="110782" lane="3" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108701" number="1" />
                    <RELAYPOSITION athleteid="108709" number="2" />
                    <RELAYPOSITION athleteid="108707" number="3" />
                    <RELAYPOSITION athleteid="108688" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="SMT Szczecin 1" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="392" reactiontime="+77" status="EXH" swimtime="00:02:22.04" resultid="108718" heatid="110715" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="75" swimtime="00:00:51.06" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="125" swimtime="00:01:29.44" />
                    <SPLIT distance="150" swimtime="00:01:50.51" />
                    <SPLIT distance="175" swimtime="00:02:05.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108679" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="108643" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="108620" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="108666" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99234" status="DNS" swimtime="00:00:00.00" resultid="108719" heatid="110780" lane="3" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108666" number="1" />
                    <RELAYPOSITION athleteid="108643" number="2" />
                    <RELAYPOSITION athleteid="108620" number="3" />
                    <RELAYPOSITION athleteid="108679" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="SMT Szczecin 1" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="283" reactiontime="+94" swimtime="00:02:05.80" resultid="108712" heatid="110632" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.50" />
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="75" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:00.82" />
                    <SPLIT distance="125" swimtime="00:01:16.72" />
                    <SPLIT distance="150" swimtime="00:01:34.00" />
                    <SPLIT distance="175" swimtime="00:01:49.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108620" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="108709" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="108707" number="3" reactiontime="+84" />
                    <RELAYPOSITION athleteid="108643" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="320" reactiontime="+86" swimtime="00:02:12.29" resultid="108713" heatid="110837" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.59" />
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="75" swimtime="00:00:52.30" />
                    <SPLIT distance="100" swimtime="00:01:11.04" />
                    <SPLIT distance="125" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:01:46.99" />
                    <SPLIT distance="175" swimtime="00:01:58.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108679" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="108628" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="108643" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="108648" number="4" reactiontime="+3" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="SMT Szczecin 2" number="2">
              <RESULTS>
                <RESULT eventid="98846" status="DNS" swimtime="00:00:00.00" resultid="108714" heatid="110632" lane="7" entrytime="00:01:50.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108679" number="1" />
                    <RELAYPOSITION athleteid="108695" number="2" />
                    <RELAYPOSITION athleteid="108666" number="3" />
                    <RELAYPOSITION athleteid="108628" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="108715" heatid="110836" lane="6" entrytime="00:02:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108643" number="1" />
                    <RELAYPOSITION athleteid="108657" number="2" />
                    <RELAYPOSITION athleteid="108695" number="3" />
                    <RELAYPOSITION athleteid="108666" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="96" agetotalmin="80" gender="X" name="SMT Szczecin 3" number="3">
              <RESULTS>
                <RESULT comment="O4/ III ZMIANA" eventid="98846" reactiontime="+92" status="DSQ" swimtime="00:00:00.00" resultid="108716" heatid="110632" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="75" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:00:58.14" />
                    <SPLIT distance="125" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:25.70" />
                    <SPLIT distance="175" swimtime="00:01:39.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108671" number="1" reactiontime="+92" status="DSQ" />
                    <RELAYPOSITION athleteid="108701" number="2" reactiontime="+29" status="DSQ" />
                    <RELAYPOSITION athleteid="108635" number="3" reactiontime="-11" status="DSQ" />
                    <RELAYPOSITION athleteid="108688" number="4" reactiontime="+78" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="350" reactiontime="+78" swimtime="00:02:08.43" resultid="108717" heatid="110837" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.62" />
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="75" swimtime="00:00:49.92" />
                    <SPLIT distance="100" swimtime="00:01:11.64" />
                    <SPLIT distance="125" swimtime="00:01:25.67" />
                    <SPLIT distance="150" swimtime="00:01:41.90" />
                    <SPLIT distance="175" swimtime="00:01:54.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108635" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="108671" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="108701" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="108688" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="109046" name="Szczecin">
          <CONTACT name="Hanczewska" phone="664935249" />
          <ATHLETES>
            <ATHLETE birthdate="1984-10-05" firstname="Marta" gender="F" lastname="Hanczewska" nation="POL" athleteid="109047">
              <RESULTS>
                <RESULT eventid="98777" points="344" reactiontime="+86" swimtime="00:00:33.16" resultid="109048" heatid="110590" lane="7" entrytime="00:00:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="294" swimtime="00:01:16.49" resultid="109049" heatid="110674" lane="6" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.67" />
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                    <SPLIT distance="75" swimtime="00:00:55.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="295" reactiontime="+99" swimtime="00:01:33.64" resultid="109050" heatid="110724" lane="1" entrytime="00:01:30.28">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.92" />
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                    <SPLIT distance="75" swimtime="00:01:07.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="268" swimtime="00:02:51.65" resultid="109051" heatid="110766" lane="6" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.15" />
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="75" swimtime="00:00:57.74" />
                    <SPLIT distance="100" swimtime="00:01:19.79" />
                    <SPLIT distance="125" swimtime="00:01:41.78" />
                    <SPLIT distance="150" swimtime="00:02:04.97" />
                    <SPLIT distance="175" swimtime="00:02:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="318" reactiontime="+95" swimtime="00:00:42.15" resultid="109052" heatid="110821" lane="4" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STP" nation="POL" region="ZAC" clubid="107796" name="Szczecineckie Towarzystwo Pływackie Masters" shortname="Szczecineckie TP Masters">
          <CONTACT city="Szczecinek" email="szczecinekmasters@wp.pl" internet="www.masters.szczecinek.pl" name="Wojnicz Andrzej" phone="887550761" street="Szczecinecka" zip="78-400" />
          <ATHLETES>
            <ATHLETE birthdate="1933-02-19" firstname="Zbigniew" gender="M" lastname="Ludwiczak" nation="POL" athleteid="107819">
              <RESULTS>
                <RESULT eventid="98798" points="55" swimtime="00:00:53.20" resultid="107820" heatid="110595" lane="6" entrytime="00:00:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="59" swimtime="00:18:52.99" resultid="107821" heatid="110638" lane="0" entrytime="00:20:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.17" />
                    <SPLIT distance="50" swimtime="00:01:00.00" />
                    <SPLIT distance="75" swimtime="00:01:31.24" />
                    <SPLIT distance="100" swimtime="00:02:04.08" />
                    <SPLIT distance="125" swimtime="00:02:37.41" />
                    <SPLIT distance="150" swimtime="00:03:11.66" />
                    <SPLIT distance="175" swimtime="00:03:45.92" />
                    <SPLIT distance="200" swimtime="00:04:20.45" />
                    <SPLIT distance="225" swimtime="00:04:54.93" />
                    <SPLIT distance="250" swimtime="00:05:29.17" />
                    <SPLIT distance="275" swimtime="00:06:03.47" />
                    <SPLIT distance="300" swimtime="00:06:37.95" />
                    <SPLIT distance="325" swimtime="00:07:12.45" />
                    <SPLIT distance="350" swimtime="00:07:47.14" />
                    <SPLIT distance="375" swimtime="00:08:21.70" />
                    <SPLIT distance="400" swimtime="00:08:56.13" />
                    <SPLIT distance="425" swimtime="00:09:30.94" />
                    <SPLIT distance="450" swimtime="00:10:06.42" />
                    <SPLIT distance="475" swimtime="00:10:41.15" />
                    <SPLIT distance="500" swimtime="00:11:16.52" />
                    <SPLIT distance="525" swimtime="00:11:51.60" />
                    <SPLIT distance="550" swimtime="00:12:26.49" />
                    <SPLIT distance="575" swimtime="00:13:02.23" />
                    <SPLIT distance="600" swimtime="00:13:37.98" />
                    <SPLIT distance="625" swimtime="00:14:13.67" />
                    <SPLIT distance="650" swimtime="00:16:05.07" />
                    <SPLIT distance="675" swimtime="00:15:29.87" />
                    <SPLIT distance="700" swimtime="00:17:17.30" />
                    <SPLIT distance="725" swimtime="00:16:41.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="42" reactiontime="+124" swimtime="00:01:03.49" resultid="107822" heatid="110651" lane="3" entrytime="00:00:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="54" swimtime="00:01:58.73" resultid="107823" heatid="110678" lane="3" entrytime="00:01:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.16" />
                    <SPLIT distance="50" swimtime="00:00:57.96" />
                    <SPLIT distance="75" swimtime="00:01:28.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="44" reactiontime="+111" swimtime="00:02:17.80" resultid="107824" heatid="110757" lane="6" entrytime="00:02:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.54" />
                    <SPLIT distance="50" swimtime="00:01:07.78" />
                    <SPLIT distance="75" swimtime="00:01:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="62" swimtime="00:04:10.50" resultid="107825" heatid="110769" lane="2" entrytime="00:04:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.40" />
                    <SPLIT distance="50" swimtime="00:00:59.50" />
                    <SPLIT distance="75" swimtime="00:01:30.59" />
                    <SPLIT distance="100" swimtime="00:02:02.55" />
                    <SPLIT distance="125" swimtime="00:02:35.43" />
                    <SPLIT distance="150" swimtime="00:03:07.86" />
                    <SPLIT distance="175" swimtime="00:03:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="42" swimtime="00:05:02.83" resultid="107826" heatid="110810" lane="3" entrytime="00:05:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.77" />
                    <SPLIT distance="50" swimtime="00:01:09.84" />
                    <SPLIT distance="75" swimtime="00:01:48.79" />
                    <SPLIT distance="100" swimtime="00:02:26.53" />
                    <SPLIT distance="125" swimtime="00:03:06.48" />
                    <SPLIT distance="150" swimtime="00:03:46.67" />
                    <SPLIT distance="175" swimtime="00:04:25.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="63" swimtime="00:08:53.29" resultid="107827" heatid="110852" lane="5" entrytime="00:10:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.33" />
                    <SPLIT distance="50" swimtime="00:01:00.35" />
                    <SPLIT distance="75" swimtime="00:01:31.92" />
                    <SPLIT distance="100" swimtime="00:02:05.18" />
                    <SPLIT distance="125" swimtime="00:02:38.33" />
                    <SPLIT distance="150" swimtime="00:03:12.45" />
                    <SPLIT distance="175" swimtime="00:03:45.68" />
                    <SPLIT distance="200" swimtime="00:04:19.44" />
                    <SPLIT distance="225" swimtime="00:04:53.30" />
                    <SPLIT distance="250" swimtime="00:05:28.12" />
                    <SPLIT distance="275" swimtime="00:06:02.11" />
                    <SPLIT distance="300" swimtime="00:06:36.29" />
                    <SPLIT distance="325" swimtime="00:07:09.99" />
                    <SPLIT distance="350" swimtime="00:07:47.58" />
                    <SPLIT distance="375" swimtime="00:08:20.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-12" firstname="Irena" gender="F" lastname="Filipowska" nation="POL" athleteid="107797">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="107798" heatid="110585" lane="5" entrytime="00:01:53.00" entrycourse="SCM" />
                <RESULT eventid="106294" points="27" reactiontime="+106" swimtime="00:01:25.29" resultid="107799" heatid="110645" lane="4" entrytime="00:01:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="12" swimtime="00:04:28.73" resultid="107800" heatid="110720" lane="4" entrytime="00:03:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:58.99" />
                    <SPLIT distance="50" swimtime="00:02:07.70" />
                    <SPLIT distance="75" swimtime="00:03:20.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="21" reactiontime="+107" swimtime="00:03:17.14" resultid="107801" heatid="110753" lane="8" entrytime="00:03:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:45.82" />
                    <SPLIT distance="75" swimtime="00:02:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="22" swimtime="00:07:03.97" resultid="107802" heatid="110806" lane="8" entrytime="00:06:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:48.48" />
                    <SPLIT distance="50" swimtime="00:01:40.86" />
                    <SPLIT distance="75" swimtime="00:02:37.04" />
                    <SPLIT distance="100" swimtime="00:03:34.22" />
                    <SPLIT distance="125" swimtime="00:04:30.85" />
                    <SPLIT distance="150" swimtime="00:05:23.30" />
                    <SPLIT distance="175" swimtime="00:06:16.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="16" swimtime="00:01:52.31" resultid="107803" heatid="110817" lane="2" entrytime="00:01:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:53.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-08-19" firstname="Zofia" gender="F" lastname="Wełk" nation="POL" athleteid="107804">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="107805" heatid="110586" lane="9" entrytime="00:01:24.00" entrycourse="SCM" />
                <RESULT eventid="98940" points="36" swimtime="00:06:47.51" resultid="107806" heatid="110661" lane="8" entrytime="00:06:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:46.98" />
                    <SPLIT distance="50" swimtime="00:01:37.64" />
                    <SPLIT distance="75" swimtime="00:02:29.16" />
                    <SPLIT distance="100" swimtime="00:03:24.05" />
                    <SPLIT distance="125" swimtime="00:04:15.18" />
                    <SPLIT distance="150" swimtime="00:05:07.62" />
                    <SPLIT distance="175" swimtime="00:06:01.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="19" swimtime="00:03:09.82" resultid="107807" heatid="110671" lane="3" entrytime="00:03:46.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:43.42" />
                    <SPLIT distance="50" swimtime="00:01:31.98" />
                    <SPLIT distance="75" swimtime="00:02:22.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="27" swimtime="00:03:26.07" resultid="107808" heatid="110721" lane="0" entrytime="00:03:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:45.13" />
                    <SPLIT distance="50" swimtime="00:01:40.01" />
                    <SPLIT distance="75" swimtime="00:02:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="9" swimtime="00:01:54.40" resultid="107809" heatid="110735" lane="3" entrytime="00:01:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:53.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="27" swimtime="00:01:34.92" resultid="107810" heatid="110817" lane="6" entrytime="00:01:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:45.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-23" firstname="Krystyna" gender="F" lastname="Witkowska" nation="POL" athleteid="107811">
              <RESULTS>
                <RESULT eventid="98777" points="27" reactiontime="+135" swimtime="00:01:16.99" resultid="107812" heatid="110586" lane="0" entrytime="00:01:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="21" reactiontime="+94" swimtime="00:01:32.62" resultid="107813" heatid="110645" lane="5" entrytime="00:01:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="29" reactiontime="+127" swimtime="00:02:44.51" resultid="107814" heatid="110671" lane="5" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.13" />
                    <SPLIT distance="50" swimtime="00:01:17.88" />
                    <SPLIT distance="75" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="20" reactiontime="+95" swimtime="00:03:22.02" resultid="107815" heatid="110752" lane="4" entrytime="00:03:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:45.58" />
                    <SPLIT distance="50" swimtime="00:01:33.77" />
                    <SPLIT distance="75" swimtime="00:02:29.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="27" reactiontime="+141" swimtime="00:06:07.76" resultid="107816" heatid="110764" lane="2" entrytime="00:06:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:40.65" />
                    <SPLIT distance="50" swimtime="00:01:24.88" />
                    <SPLIT distance="75" swimtime="00:02:11.68" />
                    <SPLIT distance="100" swimtime="00:02:58.98" />
                    <SPLIT distance="125" swimtime="00:03:46.70" />
                    <SPLIT distance="150" swimtime="00:04:36.69" />
                    <SPLIT distance="175" swimtime="00:05:23.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="107817" heatid="110817" lane="7" entrytime="00:01:50.00" entrycourse="SCM" />
                <RESULT eventid="99457" points="29" swimtime="00:12:35.94" resultid="107818" heatid="110842" lane="9" entrytime="00:12:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:39.40" />
                    <SPLIT distance="50" swimtime="00:01:23.86" />
                    <SPLIT distance="75" swimtime="00:02:11.04" />
                    <SPLIT distance="100" swimtime="00:02:59.24" />
                    <SPLIT distance="125" swimtime="00:03:48.91" />
                    <SPLIT distance="150" swimtime="00:04:37.07" />
                    <SPLIT distance="175" swimtime="00:05:25.93" />
                    <SPLIT distance="200" swimtime="00:06:13.99" />
                    <SPLIT distance="225" swimtime="00:07:02.35" />
                    <SPLIT distance="250" swimtime="00:07:50.89" />
                    <SPLIT distance="275" swimtime="00:08:39.00" />
                    <SPLIT distance="300" swimtime="00:09:26.37" />
                    <SPLIT distance="325" swimtime="00:10:13.96" />
                    <SPLIT distance="350" swimtime="00:11:02.51" />
                    <SPLIT distance="375" swimtime="00:11:50.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5130" nation="GER" region="17" clubid="107750" name="TG Lage">
          <CONTACT city="Lage" email="tg-schwimmen@gmx.de" name="Lange Ute" state="NO" street="Ringstr. 3" zip="32791" />
          <ATHLETES>
            <ATHLETE birthdate="1968-04-07" firstname="Konstantin" gender="M" lastname="Sklyar" nation="GER" license="321129" athleteid="107751">
              <RESULTS>
                <RESULT eventid="98830" points="321" reactiontime="+78" swimtime="00:02:39.95" resultid="107752" heatid="110623" lane="6" entrytime="00:02:52.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.96" />
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="75" swimtime="00:00:54.73" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="125" swimtime="00:01:39.30" />
                    <SPLIT distance="150" swimtime="00:02:03.10" />
                    <SPLIT distance="175" swimtime="00:02:22.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="363" swimtime="00:10:21.39" resultid="107753" heatid="110635" lane="9" entrytime="00:10:41.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.40" />
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="75" swimtime="00:00:52.90" />
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                    <SPLIT distance="125" swimtime="00:01:30.77" />
                    <SPLIT distance="150" swimtime="00:01:50.12" />
                    <SPLIT distance="175" swimtime="00:02:09.42" />
                    <SPLIT distance="200" swimtime="00:02:28.93" />
                    <SPLIT distance="225" swimtime="00:02:48.27" />
                    <SPLIT distance="250" swimtime="00:03:08.22" />
                    <SPLIT distance="275" swimtime="00:03:27.50" />
                    <SPLIT distance="300" swimtime="00:03:47.21" />
                    <SPLIT distance="325" swimtime="00:04:06.69" />
                    <SPLIT distance="350" swimtime="00:04:26.48" />
                    <SPLIT distance="375" swimtime="00:04:45.93" />
                    <SPLIT distance="400" swimtime="00:05:05.70" />
                    <SPLIT distance="425" swimtime="00:05:25.36" />
                    <SPLIT distance="450" swimtime="00:05:45.71" />
                    <SPLIT distance="475" swimtime="00:06:04.94" />
                    <SPLIT distance="500" swimtime="00:06:25.09" />
                    <SPLIT distance="525" swimtime="00:06:44.49" />
                    <SPLIT distance="550" swimtime="00:07:04.79" />
                    <SPLIT distance="575" swimtime="00:07:24.37" />
                    <SPLIT distance="600" swimtime="00:07:44.33" />
                    <SPLIT distance="625" swimtime="00:08:03.77" />
                    <SPLIT distance="650" swimtime="00:08:23.81" />
                    <SPLIT distance="675" swimtime="00:08:43.64" />
                    <SPLIT distance="700" swimtime="00:09:03.91" />
                    <SPLIT distance="725" swimtime="00:09:23.32" />
                    <SPLIT distance="750" swimtime="00:09:43.28" />
                    <SPLIT distance="775" swimtime="00:10:02.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="292" reactiontime="+94" swimtime="00:03:01.44" resultid="107754" heatid="110669" lane="8" entrytime="00:02:59.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.12" />
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="75" swimtime="00:01:04.07" />
                    <SPLIT distance="100" swimtime="00:01:27.35" />
                    <SPLIT distance="125" swimtime="00:01:50.85" />
                    <SPLIT distance="150" swimtime="00:02:14.74" />
                    <SPLIT distance="175" swimtime="00:02:38.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="268" swimtime="00:02:48.32" resultid="107755" heatid="110712" lane="9" entrytime="00:03:01.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.15" />
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="75" swimtime="00:00:58.47" />
                    <SPLIT distance="100" swimtime="00:01:20.70" />
                    <SPLIT distance="125" swimtime="00:01:43.96" />
                    <SPLIT distance="150" swimtime="00:02:06.05" />
                    <SPLIT distance="175" swimtime="00:02:26.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="315" reactiontime="+92" swimtime="00:01:21.67" resultid="107756" heatid="110731" lane="3" entrytime="00:01:21.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.65" />
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="75" swimtime="00:01:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="295" swimtime="00:05:53.50" resultid="107757" heatid="110790" lane="6" entrytime="00:06:08.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.91" />
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="75" swimtime="00:00:57.92" />
                    <SPLIT distance="100" swimtime="00:01:21.29" />
                    <SPLIT distance="125" swimtime="00:01:44.65" />
                    <SPLIT distance="150" swimtime="00:02:07.83" />
                    <SPLIT distance="175" swimtime="00:02:30.97" />
                    <SPLIT distance="200" swimtime="00:02:54.02" />
                    <SPLIT distance="225" swimtime="00:03:19.38" />
                    <SPLIT distance="250" swimtime="00:03:44.65" />
                    <SPLIT distance="275" swimtime="00:04:10.24" />
                    <SPLIT distance="300" swimtime="00:04:36.02" />
                    <SPLIT distance="325" swimtime="00:04:56.13" />
                    <SPLIT distance="350" swimtime="00:05:16.01" />
                    <SPLIT distance="375" swimtime="00:05:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="107758" heatid="110802" lane="1" entrytime="00:01:12.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="110113" name="TKKF Koszalin Masters">
          <CONTACT city="Koszalin" email="jakubkielar3@gmail.com" name="Kielar Jakub" phone="693193137" />
          <ATHLETES>
            <ATHLETE birthdate="1960-01-01" firstname="Dorota" gender="F" lastname="Gudaniec" nation="POL" athleteid="110169">
              <RESULTS>
                <RESULT eventid="98777" points="216" reactiontime="+97" swimtime="00:00:38.70" resultid="110170" heatid="110587" lane="4" entrytime="00:00:39.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106254" points="251" reactiontime="+72" swimtime="00:24:17.40" resultid="110171" heatid="110640" lane="7" entrytime="00:24:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.09" />
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                    <SPLIT distance="75" swimtime="00:01:04.69" />
                    <SPLIT distance="100" swimtime="00:01:28.37" />
                    <SPLIT distance="125" swimtime="00:01:52.11" />
                    <SPLIT distance="150" swimtime="00:02:16.07" />
                    <SPLIT distance="175" swimtime="00:02:40.78" />
                    <SPLIT distance="200" swimtime="00:03:04.98" />
                    <SPLIT distance="225" swimtime="00:03:29.33" />
                    <SPLIT distance="250" swimtime="00:03:53.47" />
                    <SPLIT distance="275" swimtime="00:04:17.65" />
                    <SPLIT distance="300" swimtime="00:04:41.93" />
                    <SPLIT distance="325" swimtime="00:05:06.37" />
                    <SPLIT distance="350" swimtime="00:05:31.04" />
                    <SPLIT distance="375" swimtime="00:05:55.60" />
                    <SPLIT distance="400" swimtime="00:06:20.10" />
                    <SPLIT distance="425" swimtime="00:06:44.19" />
                    <SPLIT distance="450" swimtime="00:07:08.61" />
                    <SPLIT distance="475" swimtime="00:07:33.23" />
                    <SPLIT distance="500" swimtime="00:07:58.04" />
                    <SPLIT distance="525" swimtime="00:08:22.52" />
                    <SPLIT distance="550" swimtime="00:08:46.92" />
                    <SPLIT distance="575" swimtime="00:09:11.73" />
                    <SPLIT distance="600" swimtime="00:09:36.21" />
                    <SPLIT distance="625" swimtime="00:10:00.80" />
                    <SPLIT distance="650" swimtime="00:10:25.35" />
                    <SPLIT distance="675" swimtime="00:10:49.97" />
                    <SPLIT distance="700" swimtime="00:11:14.75" />
                    <SPLIT distance="725" swimtime="00:11:39.32" />
                    <SPLIT distance="750" swimtime="00:12:03.82" />
                    <SPLIT distance="775" swimtime="00:12:28.38" />
                    <SPLIT distance="800" swimtime="00:12:52.75" />
                    <SPLIT distance="825" swimtime="00:13:17.35" />
                    <SPLIT distance="850" swimtime="00:13:42.10" />
                    <SPLIT distance="875" swimtime="00:14:07.10" />
                    <SPLIT distance="900" swimtime="00:14:31.57" />
                    <SPLIT distance="925" swimtime="00:14:55.97" />
                    <SPLIT distance="950" swimtime="00:15:20.78" />
                    <SPLIT distance="975" swimtime="00:15:45.27" />
                    <SPLIT distance="1000" swimtime="00:16:09.71" />
                    <SPLIT distance="1025" swimtime="00:16:34.08" />
                    <SPLIT distance="1050" swimtime="00:16:58.54" />
                    <SPLIT distance="1075" swimtime="00:17:23.23" />
                    <SPLIT distance="1100" swimtime="00:17:47.99" />
                    <SPLIT distance="1125" swimtime="00:18:12.38" />
                    <SPLIT distance="1150" swimtime="00:18:37.26" />
                    <SPLIT distance="1175" swimtime="00:19:01.62" />
                    <SPLIT distance="1200" swimtime="00:19:26.20" />
                    <SPLIT distance="1225" swimtime="00:19:50.82" />
                    <SPLIT distance="1250" swimtime="00:20:15.28" />
                    <SPLIT distance="1275" swimtime="00:20:39.42" />
                    <SPLIT distance="1300" swimtime="00:21:04.26" />
                    <SPLIT distance="1325" swimtime="00:21:28.63" />
                    <SPLIT distance="1350" swimtime="00:21:53.21" />
                    <SPLIT distance="1375" swimtime="00:22:17.49" />
                    <SPLIT distance="1400" swimtime="00:22:41.76" />
                    <SPLIT distance="1425" swimtime="00:23:06.14" />
                    <SPLIT distance="1450" swimtime="00:23:30.75" />
                    <SPLIT distance="1475" swimtime="00:23:54.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="186" reactiontime="+105" swimtime="00:03:55.51" resultid="110172" heatid="110663" lane="1" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.66" />
                    <SPLIT distance="50" swimtime="00:00:52.00" />
                    <SPLIT distance="75" swimtime="00:01:21.12" />
                    <SPLIT distance="100" swimtime="00:01:51.67" />
                    <SPLIT distance="125" swimtime="00:02:21.84" />
                    <SPLIT distance="150" swimtime="00:02:53.50" />
                    <SPLIT distance="175" swimtime="00:03:24.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="200" swimtime="00:01:36.86" resultid="110173" heatid="110692" lane="0" entrytime="00:01:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.93" />
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="75" swimtime="00:01:13.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="212" reactiontime="+99" swimtime="00:01:44.54" resultid="110174" heatid="110722" lane="3" entrytime="00:01:42.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.49" />
                    <SPLIT distance="50" swimtime="00:00:49.72" />
                    <SPLIT distance="75" swimtime="00:01:17.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="200" reactiontime="+99" swimtime="00:07:23.21" resultid="110175" heatid="110786" lane="7" entrytime="00:07:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.10" />
                    <SPLIT distance="50" swimtime="00:00:49.05" />
                    <SPLIT distance="75" swimtime="00:01:18.11" />
                    <SPLIT distance="100" swimtime="00:01:47.83" />
                    <SPLIT distance="125" swimtime="00:02:16.38" />
                    <SPLIT distance="150" swimtime="00:02:43.46" />
                    <SPLIT distance="175" swimtime="00:03:11.20" />
                    <SPLIT distance="200" swimtime="00:03:39.50" />
                    <SPLIT distance="225" swimtime="00:04:10.01" />
                    <SPLIT distance="250" swimtime="00:04:40.97" />
                    <SPLIT distance="275" swimtime="00:05:12.46" />
                    <SPLIT distance="300" swimtime="00:05:43.10" />
                    <SPLIT distance="325" swimtime="00:06:08.69" />
                    <SPLIT distance="350" swimtime="00:06:34.00" />
                    <SPLIT distance="375" swimtime="00:06:59.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="180" reactiontime="+81" swimtime="00:03:30.79" resultid="110176" heatid="110808" lane="4" entrytime="00:03:04.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.67" />
                    <SPLIT distance="50" swimtime="00:00:48.92" />
                    <SPLIT distance="75" swimtime="00:01:15.13" />
                    <SPLIT distance="100" swimtime="00:01:42.48" />
                    <SPLIT distance="125" swimtime="00:02:09.87" />
                    <SPLIT distance="150" swimtime="00:02:37.63" />
                    <SPLIT distance="175" swimtime="00:03:04.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="210" reactiontime="+109" swimtime="00:06:34.30" resultid="110177" heatid="110841" lane="2" entrytime="00:06:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.94" />
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                    <SPLIT distance="75" swimtime="00:01:07.66" />
                    <SPLIT distance="100" swimtime="00:01:32.10" />
                    <SPLIT distance="125" swimtime="00:01:56.82" />
                    <SPLIT distance="150" swimtime="00:02:22.22" />
                    <SPLIT distance="175" swimtime="00:02:47.55" />
                    <SPLIT distance="200" swimtime="00:03:13.25" />
                    <SPLIT distance="225" swimtime="00:03:38.63" />
                    <SPLIT distance="250" swimtime="00:04:04.15" />
                    <SPLIT distance="275" swimtime="00:04:29.86" />
                    <SPLIT distance="300" swimtime="00:04:55.54" />
                    <SPLIT distance="325" swimtime="00:05:20.77" />
                    <SPLIT distance="350" swimtime="00:05:45.67" />
                    <SPLIT distance="375" swimtime="00:06:10.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-24" firstname="Wioletta" gender="F" lastname="Pawliczek" nation="POL" athleteid="110178">
              <RESULTS>
                <RESULT eventid="98777" points="268" reactiontime="+87" swimtime="00:00:36.03" resultid="110179" heatid="110588" lane="4" entrytime="00:00:36.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="266" reactiontime="+74" swimtime="00:00:39.90" resultid="110180" heatid="110649" lane="9" entrytime="00:00:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="265" reactiontime="+90" swimtime="00:01:19.18" resultid="110181" heatid="110673" lane="3" entrytime="00:01:19.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.29" />
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="75" swimtime="00:00:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="251" reactiontime="+80" swimtime="00:01:27.23" resultid="110182" heatid="110755" lane="2" entrytime="00:01:27.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.33" />
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                    <SPLIT distance="75" swimtime="00:01:05.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="215" reactiontime="+82" swimtime="00:03:18.88" resultid="110183" heatid="110808" lane="5" entrytime="00:03:07.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.89" />
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                    <SPLIT distance="75" swimtime="00:01:09.77" />
                    <SPLIT distance="100" swimtime="00:02:26.96" />
                    <SPLIT distance="125" swimtime="00:02:00.82" />
                    <SPLIT distance="175" swimtime="00:02:53.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Michał" gender="M" lastname="Pieślak" nation="POL" athleteid="110191">
              <RESULTS>
                <RESULT eventid="98798" points="320" reactiontime="+81" swimtime="00:00:29.59" resultid="110192" heatid="110605" lane="6" entrytime="00:00:28.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="315" reactiontime="+79" swimtime="00:01:05.98" resultid="110193" heatid="110684" lane="8" entrytime="00:01:04.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.83" />
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="75" swimtime="00:00:48.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-22" firstname="Grzegorz" gender="M" lastname="Ćwikła" nation="POL" athleteid="110153">
              <RESULTS>
                <RESULT eventid="98830" points="248" reactiontime="+90" swimtime="00:02:54.42" resultid="110154" heatid="110625" lane="0" entrytime="00:02:41.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.76" />
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="75" swimtime="00:00:56.89" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                    <SPLIT distance="125" swimtime="00:01:48.23" />
                    <SPLIT distance="150" swimtime="00:02:14.55" />
                    <SPLIT distance="175" swimtime="00:02:34.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="246" reactiontime="+79" swimtime="00:11:46.99" resultid="110155" heatid="110637" lane="4" entrytime="00:11:29.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.40" />
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                    <SPLIT distance="75" swimtime="00:00:55.67" />
                    <SPLIT distance="100" swimtime="00:01:17.23" />
                    <SPLIT distance="125" swimtime="00:01:39.04" />
                    <SPLIT distance="150" swimtime="00:02:01.23" />
                    <SPLIT distance="175" swimtime="00:02:23.45" />
                    <SPLIT distance="200" swimtime="00:02:45.85" />
                    <SPLIT distance="225" swimtime="00:03:08.12" />
                    <SPLIT distance="250" swimtime="00:03:30.37" />
                    <SPLIT distance="275" swimtime="00:03:52.77" />
                    <SPLIT distance="300" swimtime="00:04:14.99" />
                    <SPLIT distance="325" swimtime="00:04:37.34" />
                    <SPLIT distance="350" swimtime="00:05:00.02" />
                    <SPLIT distance="375" swimtime="00:05:22.55" />
                    <SPLIT distance="400" swimtime="00:05:44.77" />
                    <SPLIT distance="425" swimtime="00:06:07.85" />
                    <SPLIT distance="450" swimtime="00:06:30.14" />
                    <SPLIT distance="475" swimtime="00:06:52.46" />
                    <SPLIT distance="500" swimtime="00:07:15.38" />
                    <SPLIT distance="525" swimtime="00:07:38.29" />
                    <SPLIT distance="550" swimtime="00:08:01.30" />
                    <SPLIT distance="575" swimtime="00:08:24.32" />
                    <SPLIT distance="600" swimtime="00:08:47.38" />
                    <SPLIT distance="625" swimtime="00:09:10.64" />
                    <SPLIT distance="650" swimtime="00:09:33.55" />
                    <SPLIT distance="675" swimtime="00:09:56.97" />
                    <SPLIT distance="700" swimtime="00:10:20.09" />
                    <SPLIT distance="725" swimtime="00:10:42.65" />
                    <SPLIT distance="750" swimtime="00:11:05.60" />
                    <SPLIT distance="775" swimtime="00:11:27.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="288" reactiontime="+67" swimtime="00:01:16.69" resultid="110156" heatid="110700" lane="2" entrytime="00:01:16.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.36" />
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="75" swimtime="00:00:58.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="216" reactiontime="+91" swimtime="00:01:21.52" resultid="110157" heatid="110761" lane="2" entrytime="00:01:14.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.38" />
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="75" swimtime="00:01:00.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="244" reactiontime="+68" swimtime="00:06:16.66" resultid="110158" heatid="110790" lane="8" entrytime="00:06:18.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.94" />
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="75" swimtime="00:00:59.51" />
                    <SPLIT distance="100" swimtime="00:01:21.28" />
                    <SPLIT distance="125" swimtime="00:01:48.37" />
                    <SPLIT distance="150" swimtime="00:02:14.66" />
                    <SPLIT distance="175" swimtime="00:02:39.89" />
                    <SPLIT distance="200" swimtime="00:03:05.22" />
                    <SPLIT distance="225" swimtime="00:03:32.59" />
                    <SPLIT distance="250" swimtime="00:03:59.95" />
                    <SPLIT distance="275" swimtime="00:04:26.93" />
                    <SPLIT distance="300" swimtime="00:04:53.85" />
                    <SPLIT distance="325" swimtime="00:05:14.34" />
                    <SPLIT distance="350" swimtime="00:05:35.53" />
                    <SPLIT distance="375" swimtime="00:05:57.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="224" reactiontime="+86" swimtime="00:02:53.82" resultid="110159" heatid="110815" lane="2" entrytime="00:02:34.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.58" />
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="75" swimtime="00:01:01.64" />
                    <SPLIT distance="100" swimtime="00:01:24.06" />
                    <SPLIT distance="125" swimtime="00:01:46.81" />
                    <SPLIT distance="150" swimtime="00:02:09.89" />
                    <SPLIT distance="175" swimtime="00:02:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="246" reactiontime="+87" swimtime="00:05:38.49" resultid="110160" heatid="110847" lane="1" entrytime="00:05:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.31" />
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="75" swimtime="00:00:57.49" />
                    <SPLIT distance="100" swimtime="00:01:18.85" />
                    <SPLIT distance="125" swimtime="00:01:40.69" />
                    <SPLIT distance="150" swimtime="00:02:02.73" />
                    <SPLIT distance="175" swimtime="00:02:25.51" />
                    <SPLIT distance="200" swimtime="00:02:48.28" />
                    <SPLIT distance="225" swimtime="00:03:10.18" />
                    <SPLIT distance="250" swimtime="00:03:32.47" />
                    <SPLIT distance="275" swimtime="00:03:55.25" />
                    <SPLIT distance="300" swimtime="00:04:17.10" />
                    <SPLIT distance="325" swimtime="00:04:38.87" />
                    <SPLIT distance="350" swimtime="00:04:59.36" />
                    <SPLIT distance="375" swimtime="00:05:19.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-12-01" firstname="Łukasz" gender="M" lastname="Pańczyszyn" nation="POL" athleteid="110141">
              <RESULTS>
                <RESULT eventid="98798" points="511" reactiontime="+99" swimtime="00:00:25.34" resultid="110142" heatid="110613" lane="0" entrytime="00:00:24.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="110143" heatid="110706" lane="9" entrytime="00:01:04.50" entrycourse="SCM" />
                <RESULT eventid="99170" points="538" swimtime="00:00:26.80" resultid="110144" heatid="110751" lane="0" entrytime="00:00:26.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="110145" heatid="110834" lane="8" entrytime="00:00:31.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-08" firstname="Dawid" gender="M" lastname="Borus" nation="POL" athleteid="110161">
              <RESULTS>
                <RESULT eventid="98798" points="355" reactiontime="+81" swimtime="00:00:28.61" resultid="110162" heatid="110606" lane="1" entrytime="00:00:28.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="110163" heatid="110624" lane="4" entrytime="00:02:43.00" entrycourse="SCM" />
                <RESULT eventid="98924" points="320" reactiontime="+68" swimtime="00:00:32.47" resultid="110164" heatid="110658" lane="7" entrytime="00:00:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="110165" heatid="110703" lane="8" entrytime="00:01:10.00" entrycourse="SCM" />
                <RESULT eventid="99186" points="343" reactiontime="+71" swimtime="00:01:09.87" resultid="110166" heatid="110762" lane="7" entrytime="00:01:09.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="75" swimtime="00:00:51.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="321" reactiontime="+79" swimtime="00:02:34.19" resultid="110167" heatid="110815" lane="0" entrytime="00:02:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.23" />
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="75" swimtime="00:00:54.93" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="125" swimtime="00:01:34.87" />
                    <SPLIT distance="150" swimtime="00:01:55.25" />
                    <SPLIT distance="175" swimtime="00:02:15.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="334" reactiontime="+75" swimtime="00:00:36.36" resultid="110168" heatid="110832" lane="8" entrytime="00:00:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-21" firstname="Jakub" gender="M" lastname="Kielar" nation="POL" athleteid="110119">
              <RESULTS>
                <RESULT eventid="98798" points="433" reactiontime="+71" swimtime="00:00:26.77" resultid="110120" heatid="110609" lane="6" entrytime="00:00:26.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="310" reactiontime="+87" swimtime="00:00:32.82" resultid="110121" heatid="110658" lane="1" entrytime="00:00:32.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="401" swimtime="00:01:08.67" resultid="110122" heatid="110705" lane="0" entrytime="00:01:06.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.35" />
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="75" swimtime="00:00:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="450" swimtime="00:00:28.44" resultid="110123" heatid="110750" lane="9" entrytime="00:00:27.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="309" reactiontime="+80" swimtime="00:01:12.36" resultid="110124" heatid="110762" lane="2" entrytime="00:01:09.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.92" />
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="75" swimtime="00:00:53.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="381" reactiontime="+82" swimtime="00:01:06.79" resultid="110125" heatid="110804" lane="8" entrytime="00:01:07.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="75" swimtime="00:00:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="363" swimtime="00:00:35.37" resultid="110126" heatid="110833" lane="9" entrytime="00:00:34.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-05" firstname="Agnieszka" gender="F" lastname="Paziewska" nation="POL" athleteid="110127">
              <RESULTS>
                <RESULT eventid="98777" points="328" reactiontime="+115" swimtime="00:00:33.67" resultid="110128" heatid="110591" lane="6" entrytime="00:00:31.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="190" swimtime="00:00:44.60" resultid="110129" heatid="110648" lane="3" entrytime="00:00:39.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="293" swimtime="00:01:16.63" resultid="110130" heatid="110675" lane="0" entrytime="00:01:12.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.45" />
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="75" swimtime="00:00:55.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="219" reactiontime="+117" swimtime="00:01:43.34" resultid="110131" heatid="110723" lane="7" entrytime="00:01:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.69" />
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                    <SPLIT distance="75" swimtime="00:01:14.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="257" reactiontime="+124" swimtime="00:02:54.16" resultid="110132" heatid="110767" lane="1" entrytime="00:02:42.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.51" />
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="75" swimtime="00:00:57.29" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="125" swimtime="00:01:42.79" />
                    <SPLIT distance="150" swimtime="00:02:07.01" />
                    <SPLIT distance="175" swimtime="00:02:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="257" reactiontime="+119" swimtime="00:00:45.27" resultid="110133" heatid="110820" lane="5" entrytime="00:00:43.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Janusz" gender="M" lastname="Dudziński" nation="POL" athleteid="110184">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="110185" heatid="110604" lane="7" entrytime="00:00:29.80" entrycourse="SCM" />
                <RESULT eventid="98956" status="WDR" swimtime="00:00:00.00" resultid="110186" heatid="110668" lane="7" entrytime="00:03:07.00" entrycourse="SCM" />
                <RESULT eventid="98988" status="WDR" swimtime="00:00:00.00" resultid="110187" heatid="110699" lane="2" entrytime="00:01:19.60" entrycourse="SCM" />
                <RESULT eventid="99282" status="WDR" swimtime="00:00:00.00" resultid="110189" heatid="110791" lane="9" entrytime="00:05:59.00" entrycourse="SCM" />
                <RESULT eventid="99425" status="WDR" swimtime="00:00:00.00" resultid="110190" heatid="110829" lane="3" entrytime="00:00:37.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-03-02" firstname="Andrzej" gender="M" lastname="Michałkowski" nation="POL" athleteid="110146">
              <RESULTS>
                <RESULT eventid="98798" points="108" reactiontime="+92" swimtime="00:00:42.42" resultid="110147" heatid="110596" lane="1" entrytime="00:00:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="87" reactiontime="+92" swimtime="00:04:06.65" resultid="110148" heatid="110620" lane="8" entrytime="00:03:58.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.56" />
                    <SPLIT distance="50" swimtime="00:00:50.78" />
                    <SPLIT distance="75" swimtime="00:01:28.61" />
                    <SPLIT distance="100" swimtime="00:02:06.72" />
                    <SPLIT distance="125" swimtime="00:02:38.67" />
                    <SPLIT distance="150" swimtime="00:03:10.89" />
                    <SPLIT distance="175" swimtime="00:03:39.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="123" reactiontime="+103" swimtime="00:04:01.93" resultid="110149" heatid="110666" lane="7" entrytime="00:03:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.96" />
                    <SPLIT distance="50" swimtime="00:00:51.09" />
                    <SPLIT distance="75" swimtime="00:01:20.57" />
                    <SPLIT distance="100" swimtime="00:01:52.16" />
                    <SPLIT distance="125" swimtime="00:02:24.52" />
                    <SPLIT distance="150" swimtime="00:02:57.51" />
                    <SPLIT distance="175" swimtime="00:03:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="110" reactiontime="+83" swimtime="00:01:45.48" resultid="110150" heatid="110697" lane="8" entrytime="00:01:45.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.98" />
                    <SPLIT distance="50" swimtime="00:00:52.97" />
                    <SPLIT distance="75" swimtime="00:01:20.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="161" reactiontime="+91" swimtime="00:01:42.07" resultid="110151" heatid="110728" lane="4" entrytime="00:01:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.09" />
                    <SPLIT distance="50" swimtime="00:00:46.19" />
                    <SPLIT distance="75" swimtime="00:01:13.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="210" reactiontime="+96" swimtime="00:00:42.42" resultid="110152" heatid="110826" lane="4" entrytime="00:00:42.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-06" firstname="Joanna" gender="F" lastname="Stankiewicz - Majkowska" nation="POL" athleteid="110134">
              <RESULTS>
                <RESULT eventid="98814" points="193" reactiontime="+98" swimtime="00:03:30.68" resultid="110135" heatid="110615" lane="2" entrytime="00:03:29.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.57" />
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                    <SPLIT distance="75" swimtime="00:01:12.98" />
                    <SPLIT distance="100" swimtime="00:01:39.00" />
                    <SPLIT distance="125" swimtime="00:02:07.34" />
                    <SPLIT distance="150" swimtime="00:02:36.64" />
                    <SPLIT distance="175" swimtime="00:03:04.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="110136" heatid="110691" lane="4" entrytime="00:01:35.50" entrycourse="SCM" />
                <RESULT eventid="99004" points="146" swimtime="00:03:47.02" resultid="110137" heatid="110708" lane="9" entrytime="00:03:44.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.61" />
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                    <SPLIT distance="75" swimtime="00:01:20.20" />
                    <SPLIT distance="100" swimtime="00:01:49.03" />
                    <SPLIT distance="125" swimtime="00:02:17.61" />
                    <SPLIT distance="150" swimtime="00:02:47.80" />
                    <SPLIT distance="175" swimtime="00:03:16.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="206" swimtime="00:01:45.49" resultid="110138" heatid="110722" lane="0" entrytime="00:01:48.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.78" />
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                    <SPLIT distance="75" swimtime="00:01:16.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="200" reactiontime="+112" swimtime="00:07:23.34" resultid="110139" heatid="110786" lane="1" entrytime="00:07:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.51" />
                    <SPLIT distance="50" swimtime="00:00:51.98" />
                    <SPLIT distance="75" swimtime="00:01:21.22" />
                    <SPLIT distance="100" swimtime="00:01:51.23" />
                    <SPLIT distance="125" swimtime="00:02:20.62" />
                    <SPLIT distance="150" swimtime="00:02:47.91" />
                    <SPLIT distance="175" swimtime="00:03:15.59" />
                    <SPLIT distance="200" swimtime="00:03:42.78" />
                    <SPLIT distance="225" swimtime="00:04:11.04" />
                    <SPLIT distance="250" swimtime="00:04:39.32" />
                    <SPLIT distance="275" swimtime="00:05:08.55" />
                    <SPLIT distance="300" swimtime="00:05:38.56" />
                    <SPLIT distance="325" swimtime="00:06:05.18" />
                    <SPLIT distance="350" swimtime="00:06:32.30" />
                    <SPLIT distance="375" swimtime="00:06:57.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="207" reactiontime="+81" swimtime="00:00:48.61" resultid="110140" heatid="110820" lane="1" entrytime="00:00:45.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="399" reactiontime="+70" swimtime="00:02:02.86" resultid="110194" heatid="110719" lane="7" entrytime="00:01:59.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.11" />
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="75" swimtime="00:00:47.82" />
                    <SPLIT distance="100" swimtime="00:01:05.51" />
                    <SPLIT distance="125" swimtime="00:01:18.44" />
                    <SPLIT distance="150" swimtime="00:01:33.70" />
                    <SPLIT distance="175" swimtime="00:01:47.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110161" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="110141" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="110119" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="110191" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="434" swimtime="00:01:49.03" resultid="110195" heatid="110784" lane="0" entrytime="00:01:48.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:24.89" />
                    <SPLIT distance="75" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:00:54.42" />
                    <SPLIT distance="125" swimtime="00:01:07.40" />
                    <SPLIT distance="150" swimtime="00:01:22.04" />
                    <SPLIT distance="175" swimtime="00:01:34.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110119" number="1" />
                    <RELAYPOSITION athleteid="110161" number="2" />
                    <RELAYPOSITION athleteid="110191" number="3" />
                    <RELAYPOSITION athleteid="110141" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99234" points="253" reactiontime="+103" swimtime="00:02:28.89" resultid="110200" heatid="110779" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.91" />
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="75" swimtime="00:00:57.83" />
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="125" swimtime="00:01:36.46" />
                    <SPLIT distance="150" swimtime="00:01:54.71" />
                    <SPLIT distance="175" swimtime="00:02:10.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110169" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="110134" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="110178" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="110127" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99036" points="257" reactiontime="+81" swimtime="00:02:43.44" resultid="110201" heatid="110714" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.37" />
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="75" swimtime="00:01:00.50" />
                    <SPLIT distance="100" swimtime="00:01:25.90" />
                    <SPLIT distance="125" swimtime="00:01:45.93" />
                    <SPLIT distance="150" swimtime="00:02:10.22" />
                    <SPLIT distance="175" swimtime="00:02:25.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110178" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="110134" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="110169" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="110127" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="299" reactiontime="+67" swimtime="00:02:03.48" resultid="110196" heatid="110631" lane="6" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.07" />
                    <SPLIT distance="50" swimtime="00:00:25.07" />
                    <SPLIT distance="75" swimtime="00:00:43.63" />
                    <SPLIT distance="100" swimtime="00:01:03.55" />
                    <SPLIT distance="125" swimtime="00:01:19.20" />
                    <SPLIT distance="150" swimtime="00:01:36.85" />
                    <SPLIT distance="175" swimtime="00:01:49.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110119" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="110169" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="110127" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="110141" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="99441" points="253" reactiontime="+72" swimtime="00:02:22.99" resultid="110199" heatid="110838" lane="9" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.72" />
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                    <SPLIT distance="75" swimtime="00:00:59.82" />
                    <SPLIT distance="100" swimtime="00:01:25.01" />
                    <SPLIT distance="125" swimtime="00:01:38.01" />
                    <SPLIT distance="150" swimtime="00:01:53.79" />
                    <SPLIT distance="175" swimtime="00:02:07.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110178" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="110141" number="2" />
                    <RELAYPOSITION athleteid="110119" number="3" />
                    <RELAYPOSITION athleteid="110127" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="217" reactiontime="+59" swimtime="00:02:17.43" resultid="110197" heatid="110630" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.53" />
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                    <SPLIT distance="75" swimtime="00:00:47.55" />
                    <SPLIT distance="100" swimtime="00:01:06.61" />
                    <SPLIT distance="125" swimtime="00:01:26.08" />
                    <SPLIT distance="150" swimtime="00:01:47.82" />
                    <SPLIT distance="175" swimtime="00:02:01.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110153" number="1" reactiontime="+59" />
                    <RELAYPOSITION athleteid="110178" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="110134" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="110191" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="192" reactiontime="+79" swimtime="00:02:36.74" resultid="110198" heatid="110836" lane="5" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.94" />
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                    <SPLIT distance="75" swimtime="00:01:03.36" />
                    <SPLIT distance="100" swimtime="00:01:23.68" />
                    <SPLIT distance="125" swimtime="00:01:39.07" />
                    <SPLIT distance="150" swimtime="00:01:57.57" />
                    <SPLIT distance="175" swimtime="00:02:16.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110134" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="110161" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="110153" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="110169" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="107057" name="Torpedos">
          <CONTACT email="vilmantasenator@gmail.com" name="Vilmantas Krasauskas" phone="+37068746068" street="Jukneviciaus 78-10" zip="68198" />
          <ATHLETES>
            <ATHLETE birthdate="1956-02-07" firstname="Margarita" gender="F" lastname="Cineliene" nation="LTU" athleteid="107083">
              <RESULTS>
                <RESULT eventid="98972" points="144" reactiontime="+98" swimtime="00:01:47.99" resultid="107084" heatid="110691" lane="8" entrytime="00:01:47.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.46" />
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                    <SPLIT distance="75" swimtime="00:01:19.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="204" reactiontime="+103" swimtime="00:01:45.93" resultid="107085" heatid="110723" lane="2" entrytime="00:01:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.86" />
                    <SPLIT distance="50" swimtime="00:00:49.36" />
                    <SPLIT distance="75" swimtime="00:01:17.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="239" reactiontime="+103" swimtime="00:00:46.39" resultid="107086" heatid="110819" lane="4" entrytime="00:00:46.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-04" firstname="Jurate" gender="F" lastname="Pranckeviciene" nation="LTU" athleteid="107065">
              <RESULTS>
                <RESULT eventid="98907" points="313" reactiontime="+92" swimtime="00:01:14.94" resultid="107066" heatid="110674" lane="1" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="75" swimtime="00:00:55.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="255" reactiontime="+80" swimtime="00:00:38.44" resultid="107067" heatid="110737" lane="5" entrytime="00:00:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="200" reactiontime="+89" swimtime="00:03:23.64" resultid="107068" heatid="110807" lane="3" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.78" />
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                    <SPLIT distance="75" swimtime="00:01:13.41" />
                    <SPLIT distance="100" swimtime="00:01:39.95" />
                    <SPLIT distance="125" swimtime="00:02:06.86" />
                    <SPLIT distance="150" swimtime="00:02:33.68" />
                    <SPLIT distance="175" swimtime="00:02:59.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-07-31" firstname="Vilmantas" gender="M" lastname="Krasauskas" nation="LTU" athleteid="107076">
              <RESULTS>
                <RESULT eventid="106277" points="387" reactiontime="+86" swimtime="00:01:01.66" resultid="107077" heatid="110684" lane="3" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.29" />
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="75" swimtime="00:00:45.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="387" reactiontime="+78" swimtime="00:02:16.31" resultid="107078" heatid="110775" lane="7" entrytime="00:02:21.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.04" />
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="75" swimtime="00:00:48.57" />
                    <SPLIT distance="100" swimtime="00:01:05.87" />
                    <SPLIT distance="125" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:01:41.23" />
                    <SPLIT distance="175" swimtime="00:01:59.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="360" reactiontime="+82" swimtime="00:04:58.11" resultid="107079" heatid="110845" lane="7" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.09" />
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="75" swimtime="00:00:52.03" />
                    <SPLIT distance="100" swimtime="00:01:10.32" />
                    <SPLIT distance="125" swimtime="00:01:28.33" />
                    <SPLIT distance="150" swimtime="00:01:46.85" />
                    <SPLIT distance="175" swimtime="00:02:05.31" />
                    <SPLIT distance="200" swimtime="00:02:24.13" />
                    <SPLIT distance="225" swimtime="00:02:43.01" />
                    <SPLIT distance="250" swimtime="00:03:01.94" />
                    <SPLIT distance="275" swimtime="00:03:21.18" />
                    <SPLIT distance="300" swimtime="00:03:40.63" />
                    <SPLIT distance="325" swimtime="00:03:59.91" />
                    <SPLIT distance="350" swimtime="00:04:19.67" />
                    <SPLIT distance="375" swimtime="00:04:39.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-03-14" firstname="Stasys" gender="M" lastname="Grigas" nation="LTU" athleteid="107069">
              <RESULTS>
                <RESULT eventid="98924" points="41" reactiontime="+114" swimtime="00:01:04.25" resultid="107070" heatid="110651" lane="2" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="33" reactiontime="+116" swimtime="00:02:19.03" resultid="107071" heatid="110678" lane="7" entrytime="00:02:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.17" />
                    <SPLIT distance="50" swimtime="00:01:04.44" />
                    <SPLIT distance="75" swimtime="00:01:41.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="39" reactiontime="+123" swimtime="00:02:43.37" resultid="107072" heatid="110727" lane="8" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.56" />
                    <SPLIT distance="50" swimtime="00:01:19.69" />
                    <SPLIT distance="75" swimtime="00:02:02.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="39" reactiontime="+111" swimtime="00:02:23.91" resultid="107073" heatid="110757" lane="2" entrytime="00:02:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.41" />
                    <SPLIT distance="50" swimtime="00:01:08.90" />
                    <SPLIT distance="75" swimtime="00:01:46.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="37" reactiontime="+121" swimtime="00:05:16.12" resultid="107074" heatid="110810" lane="6" entrytime="00:05:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.95" />
                    <SPLIT distance="50" swimtime="00:01:12.94" />
                    <SPLIT distance="75" swimtime="00:01:51.16" />
                    <SPLIT distance="100" swimtime="00:02:32.93" />
                    <SPLIT distance="125" swimtime="00:03:15.50" />
                    <SPLIT distance="150" swimtime="00:03:57.17" />
                    <SPLIT distance="175" swimtime="00:04:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="67" swimtime="00:01:02.04" resultid="107075" heatid="110824" lane="6" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-11-15" firstname="Aldona" gender="F" lastname="Mazetiene" nation="LTU" athleteid="107080">
              <RESULTS>
                <RESULT eventid="106294" points="103" reactiontime="+103" swimtime="00:00:54.66" resultid="107081" heatid="110647" lane="0" entrytime="00:00:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="115" swimtime="00:00:59.10" resultid="107082" heatid="110818" lane="2" entrytime="00:00:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="KUJ" clubid="107426" name="Toruń Multisport Team">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="107489">
              <RESULTS>
                <RESULT eventid="98798" points="240" reactiontime="+82" swimtime="00:00:32.57" resultid="107490" heatid="110600" lane="6" entrytime="00:00:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="148" reactiontime="+83" swimtime="00:03:27.02" resultid="107491" heatid="110621" lane="3" entrytime="00:03:18.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.43" />
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="75" swimtime="00:01:12.16" />
                    <SPLIT distance="100" swimtime="00:01:40.74" />
                    <SPLIT distance="125" swimtime="00:02:12.71" />
                    <SPLIT distance="150" swimtime="00:02:43.12" />
                    <SPLIT distance="175" swimtime="00:03:06.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="215" reactiontime="+92" swimtime="00:01:24.45" resultid="107492" heatid="110698" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.93" />
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="75" swimtime="00:01:05.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="213" swimtime="00:00:36.47" resultid="107493" heatid="110744" lane="9" entrytime="00:00:35.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="199" reactiontime="+69" swimtime="00:02:49.98" resultid="107494" heatid="110771" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.90" />
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                    <SPLIT distance="75" swimtime="00:01:00.71" />
                    <SPLIT distance="100" swimtime="00:01:22.97" />
                    <SPLIT distance="125" swimtime="00:01:45.54" />
                    <SPLIT distance="150" swimtime="00:02:08.39" />
                    <SPLIT distance="175" swimtime="00:02:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="168" reactiontime="+92" swimtime="00:06:23.96" resultid="107495" heatid="110849" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.81" />
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="75" swimtime="00:01:02.86" />
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                    <SPLIT distance="125" swimtime="00:01:47.93" />
                    <SPLIT distance="150" swimtime="00:02:11.17" />
                    <SPLIT distance="175" swimtime="00:02:34.74" />
                    <SPLIT distance="200" swimtime="00:03:00.10" />
                    <SPLIT distance="225" swimtime="00:03:25.43" />
                    <SPLIT distance="250" swimtime="00:03:51.32" />
                    <SPLIT distance="275" swimtime="00:04:17.58" />
                    <SPLIT distance="300" swimtime="00:04:42.05" />
                    <SPLIT distance="325" swimtime="00:05:07.32" />
                    <SPLIT distance="350" swimtime="00:05:32.56" />
                    <SPLIT distance="375" swimtime="00:05:59.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-23" firstname="Marcin" gender="M" lastname="Mykowski" nation="POL" athleteid="107432">
              <RESULTS>
                <RESULT eventid="98891" points="343" reactiontime="+100" swimtime="00:10:33.35" resultid="107433" heatid="110636" lane="2" entrytime="00:10:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.78" />
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                    <SPLIT distance="75" swimtime="00:00:56.20" />
                    <SPLIT distance="100" swimtime="00:01:16.78" />
                    <SPLIT distance="125" swimtime="00:01:37.13" />
                    <SPLIT distance="150" swimtime="00:01:57.32" />
                    <SPLIT distance="175" swimtime="00:02:17.85" />
                    <SPLIT distance="200" swimtime="00:02:38.03" />
                    <SPLIT distance="225" swimtime="00:02:58.80" />
                    <SPLIT distance="250" swimtime="00:03:19.58" />
                    <SPLIT distance="275" swimtime="00:03:40.23" />
                    <SPLIT distance="300" swimtime="00:04:00.69" />
                    <SPLIT distance="325" swimtime="00:04:21.29" />
                    <SPLIT distance="350" swimtime="00:04:41.98" />
                    <SPLIT distance="375" swimtime="00:05:02.17" />
                    <SPLIT distance="400" swimtime="00:05:22.43" />
                    <SPLIT distance="425" swimtime="00:05:42.34" />
                    <SPLIT distance="450" swimtime="00:06:02.13" />
                    <SPLIT distance="475" swimtime="00:06:22.24" />
                    <SPLIT distance="500" swimtime="00:06:42.14" />
                    <SPLIT distance="525" swimtime="00:07:02.15" />
                    <SPLIT distance="550" swimtime="00:07:22.15" />
                    <SPLIT distance="575" swimtime="00:07:42.60" />
                    <SPLIT distance="600" swimtime="00:08:02.99" />
                    <SPLIT distance="625" swimtime="00:08:21.80" />
                    <SPLIT distance="650" swimtime="00:08:40.81" />
                    <SPLIT distance="675" swimtime="00:09:00.27" />
                    <SPLIT distance="700" swimtime="00:09:19.72" />
                    <SPLIT distance="725" swimtime="00:09:38.60" />
                    <SPLIT distance="750" swimtime="00:09:57.23" />
                    <SPLIT distance="775" swimtime="00:10:15.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="468" reactiontime="+75" swimtime="00:00:57.85" resultid="107434" heatid="110687" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                    <SPLIT distance="75" swimtime="00:00:42.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="107439">
              <RESULTS>
                <RESULT eventid="98830" points="52" reactiontime="+140" swimtime="00:04:53.71" resultid="107440" heatid="110619" lane="5" entrytime="00:04:31.78">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.29" />
                    <SPLIT distance="50" swimtime="00:01:07.23" />
                    <SPLIT distance="75" swimtime="00:01:52.72" />
                    <SPLIT distance="100" swimtime="00:02:33.87" />
                    <SPLIT distance="125" swimtime="00:03:17.27" />
                    <SPLIT distance="150" swimtime="00:03:58.20" />
                    <SPLIT distance="175" swimtime="00:04:25.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="62" reactiontime="+126" swimtime="00:05:04.12" resultid="107441" heatid="110665" lane="4" entrytime="00:04:37.51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.16" />
                    <SPLIT distance="50" swimtime="00:01:13.29" />
                    <SPLIT distance="75" swimtime="00:01:52.48" />
                    <SPLIT distance="100" swimtime="00:02:32.66" />
                    <SPLIT distance="125" swimtime="00:03:11.94" />
                    <SPLIT distance="150" swimtime="00:03:50.69" />
                    <SPLIT distance="175" swimtime="00:04:28.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="33" swimtime="00:05:37.82" resultid="107442" heatid="110710" lane="0" entrytime="00:05:08.04">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.67" />
                    <SPLIT distance="50" swimtime="00:01:14.37" />
                    <SPLIT distance="75" swimtime="00:01:55.48" />
                    <SPLIT distance="100" swimtime="00:02:37.89" />
                    <SPLIT distance="125" swimtime="00:03:21.40" />
                    <SPLIT distance="150" swimtime="00:04:07.88" />
                    <SPLIT distance="175" swimtime="00:04:52.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="65" swimtime="00:04:07.00" resultid="107443" heatid="110770" lane="0" entrytime="00:03:42.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.90" />
                    <SPLIT distance="50" swimtime="00:00:54.29" />
                    <SPLIT distance="75" swimtime="00:01:25.51" />
                    <SPLIT distance="100" swimtime="00:01:57.43" />
                    <SPLIT distance="125" swimtime="00:02:30.37" />
                    <SPLIT distance="150" swimtime="00:03:03.65" />
                    <SPLIT distance="175" swimtime="00:03:37.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="45" reactiontime="+129" swimtime="00:10:59.09" resultid="107444" heatid="110788" lane="8" entrytime="00:09:58.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.71" />
                    <SPLIT distance="50" swimtime="00:01:16.29" />
                    <SPLIT distance="75" swimtime="00:01:59.42" />
                    <SPLIT distance="100" swimtime="00:02:45.12" />
                    <SPLIT distance="125" swimtime="00:03:33.26" />
                    <SPLIT distance="150" swimtime="00:04:19.58" />
                    <SPLIT distance="175" swimtime="00:05:05.32" />
                    <SPLIT distance="200" swimtime="00:05:47.88" />
                    <SPLIT distance="225" swimtime="00:06:35.57" />
                    <SPLIT distance="250" swimtime="00:07:21.02" />
                    <SPLIT distance="275" swimtime="00:08:06.59" />
                    <SPLIT distance="300" swimtime="00:08:53.17" />
                    <SPLIT distance="325" swimtime="00:09:25.54" />
                    <SPLIT distance="350" swimtime="00:09:59.44" />
                    <SPLIT distance="375" swimtime="00:10:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="28" reactiontime="+128" swimtime="00:02:38.25" resultid="107445" heatid="110798" lane="8" entrytime="00:02:15.98">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.78" />
                    <SPLIT distance="50" swimtime="00:01:13.29" />
                    <SPLIT distance="75" swimtime="00:01:55.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="29" reactiontime="+103" swimtime="00:05:41.53" resultid="107446" heatid="110810" lane="5" entrytime="00:05:10.41">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:38.11" />
                    <SPLIT distance="50" swimtime="00:01:24.05" />
                    <SPLIT distance="75" swimtime="00:02:05.22" />
                    <SPLIT distance="100" swimtime="00:02:48.87" />
                    <SPLIT distance="125" swimtime="00:03:31.96" />
                    <SPLIT distance="150" swimtime="00:04:16.86" />
                    <SPLIT distance="175" swimtime="00:05:00.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="107481">
              <RESULTS>
                <RESULT eventid="98814" points="444" reactiontime="+87" swimtime="00:02:39.67" resultid="107482" heatid="110618" lane="1" entrytime="00:02:41.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.20" />
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="75" swimtime="00:00:54.53" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="125" swimtime="00:01:37.32" />
                    <SPLIT distance="150" swimtime="00:02:01.07" />
                    <SPLIT distance="175" swimtime="00:02:20.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="447" swimtime="00:02:55.96" resultid="107483" heatid="110664" lane="6" entrytime="00:02:58.97">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.46" />
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="75" swimtime="00:01:01.90" />
                    <SPLIT distance="100" swimtime="00:01:24.18" />
                    <SPLIT distance="125" swimtime="00:01:46.60" />
                    <SPLIT distance="150" swimtime="00:02:09.49" />
                    <SPLIT distance="175" swimtime="00:02:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="460" swimtime="00:01:13.39" resultid="107484" heatid="110695" lane="0" entrytime="00:01:14.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.05" />
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="75" swimtime="00:00:55.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="429" swimtime="00:01:22.65" resultid="107485" heatid="110725" lane="9" entrytime="00:01:23.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.26" />
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                    <SPLIT distance="75" swimtime="00:01:00.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="423" reactiontime="+85" swimtime="00:05:45.59" resultid="107486" heatid="110787" lane="3" entrytime="00:05:54.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.93" />
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="75" swimtime="00:00:56.00" />
                    <SPLIT distance="100" swimtime="00:01:17.81" />
                    <SPLIT distance="125" swimtime="00:01:40.98" />
                    <SPLIT distance="150" swimtime="00:02:02.93" />
                    <SPLIT distance="175" swimtime="00:02:24.79" />
                    <SPLIT distance="200" swimtime="00:02:46.58" />
                    <SPLIT distance="225" swimtime="00:03:10.76" />
                    <SPLIT distance="250" swimtime="00:03:34.72" />
                    <SPLIT distance="275" swimtime="00:03:58.93" />
                    <SPLIT distance="300" swimtime="00:04:23.48" />
                    <SPLIT distance="325" swimtime="00:04:44.54" />
                    <SPLIT distance="350" swimtime="00:05:05.23" />
                    <SPLIT distance="375" swimtime="00:05:25.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="427" reactiontime="+87" swimtime="00:00:38.24" resultid="107487" heatid="110822" lane="3" entrytime="00:00:38.57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="406" reactiontime="+89" swimtime="00:05:16.49" resultid="107488" heatid="110841" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.21" />
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="75" swimtime="00:00:56.85" />
                    <SPLIT distance="100" swimtime="00:01:17.07" />
                    <SPLIT distance="125" swimtime="00:01:37.96" />
                    <SPLIT distance="150" swimtime="00:01:58.59" />
                    <SPLIT distance="175" swimtime="00:02:18.78" />
                    <SPLIT distance="200" swimtime="00:02:39.51" />
                    <SPLIT distance="225" swimtime="00:02:59.69" />
                    <SPLIT distance="250" swimtime="00:03:20.01" />
                    <SPLIT distance="275" swimtime="00:03:40.16" />
                    <SPLIT distance="300" swimtime="00:03:59.96" />
                    <SPLIT distance="325" swimtime="00:04:19.24" />
                    <SPLIT distance="350" swimtime="00:04:39.07" />
                    <SPLIT distance="375" swimtime="00:04:58.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="107447">
              <RESULTS>
                <RESULT eventid="98798" points="119" reactiontime="+112" swimtime="00:00:41.15" resultid="107448" heatid="110596" lane="6" entrytime="00:00:41.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="42" reactiontime="+86" swimtime="00:01:03.68" resultid="107449" heatid="110651" lane="6" entrytime="00:01:06.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="107450" heatid="110678" lane="4" entrytime="00:01:42.10" />
                <RESULT eventid="99186" points="40" reactiontime="+106" swimtime="00:02:22.74" resultid="107451" heatid="110757" lane="3" entrytime="00:02:14.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.20" />
                    <SPLIT distance="50" swimtime="00:01:05.06" />
                    <SPLIT distance="75" swimtime="00:01:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="36" reactiontime="+100" swimtime="00:05:18.00" resultid="107452" heatid="110811" lane="9" entrytime="00:04:40.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.23" />
                    <SPLIT distance="50" swimtime="00:01:14.15" />
                    <SPLIT distance="75" swimtime="00:01:56.72" />
                    <SPLIT distance="100" swimtime="00:02:36.33" />
                    <SPLIT distance="125" swimtime="00:03:19.82" />
                    <SPLIT distance="150" swimtime="00:03:59.76" />
                    <SPLIT distance="175" swimtime="00:04:39.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-15" firstname="Artur" gender="M" lastname="Rybicki" nation="POL" athleteid="107501">
              <RESULTS>
                <RESULT eventid="98798" points="407" reactiontime="+80" swimtime="00:00:27.32" resultid="107502" heatid="110606" lane="5" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="264" reactiontime="+74" swimtime="00:00:34.63" resultid="107503" heatid="110655" lane="5" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="376" reactiontime="+79" swimtime="00:01:02.21" resultid="107504" heatid="110684" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.20" />
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="75" swimtime="00:00:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="273" reactiontime="+81" swimtime="00:00:33.59" resultid="107505" heatid="110745" lane="7" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="241" reactiontime="+84" swimtime="00:02:39.62" resultid="107506" heatid="110771" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.75" />
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="75" swimtime="00:00:55.64" />
                    <SPLIT distance="100" swimtime="00:01:16.77" />
                    <SPLIT distance="125" swimtime="00:01:38.18" />
                    <SPLIT distance="150" swimtime="00:02:00.29" />
                    <SPLIT distance="175" swimtime="00:02:21.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="210" reactiontime="+88" swimtime="00:05:56.58" resultid="107507" heatid="110849" lane="3" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.13" />
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="75" swimtime="00:01:00.63" />
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                    <SPLIT distance="125" swimtime="00:01:45.35" />
                    <SPLIT distance="150" swimtime="00:02:08.03" />
                    <SPLIT distance="175" swimtime="00:02:31.05" />
                    <SPLIT distance="200" swimtime="00:02:54.70" />
                    <SPLIT distance="225" swimtime="00:03:18.40" />
                    <SPLIT distance="250" swimtime="00:03:41.92" />
                    <SPLIT distance="275" swimtime="00:04:05.60" />
                    <SPLIT distance="300" swimtime="00:04:29.59" />
                    <SPLIT distance="325" swimtime="00:04:53.19" />
                    <SPLIT distance="350" swimtime="00:05:16.26" />
                    <SPLIT distance="375" swimtime="00:05:38.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-24" firstname="Anita" gender="F" lastname="Śliwa" nation="POL" athleteid="107463">
              <RESULTS>
                <RESULT eventid="98777" points="224" reactiontime="+119" swimtime="00:00:38.21" resultid="107464" heatid="110588" lane="0" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="205" reactiontime="+99" swimtime="00:00:43.48" resultid="107465" heatid="110648" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="98972" points="175" reactiontime="+97" swimtime="00:01:41.28" resultid="107466" heatid="110691" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.94" />
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                    <SPLIT distance="75" swimtime="00:01:17.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="187" reactiontime="+90" swimtime="00:01:36.23" resultid="107467" heatid="110754" lane="4" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.28" />
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                    <SPLIT distance="75" swimtime="00:01:11.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="107456">
              <RESULTS>
                <RESULT eventid="98798" points="83" reactiontime="+87" swimtime="00:00:46.35" resultid="107457" heatid="110596" lane="8" entrytime="00:00:43.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="79" reactiontime="+80" swimtime="00:00:51.63" resultid="107458" heatid="110651" lane="5" entrytime="00:00:58.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="81" swimtime="00:04:37.78" resultid="107459" heatid="110666" lane="9" entrytime="00:04:22.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.92" />
                    <SPLIT distance="50" swimtime="00:01:00.34" />
                    <SPLIT distance="75" swimtime="00:01:34.71" />
                    <SPLIT distance="100" swimtime="00:02:10.71" />
                    <SPLIT distance="125" swimtime="00:02:47.17" />
                    <SPLIT distance="150" swimtime="00:03:24.65" />
                    <SPLIT distance="175" swimtime="00:04:02.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="95" reactiontime="+107" swimtime="00:02:01.70" resultid="107460" heatid="110727" lane="2" entrytime="00:01:59.03">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.47" />
                    <SPLIT distance="50" swimtime="00:00:55.74" />
                    <SPLIT distance="75" swimtime="00:01:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="107461" heatid="110758" lane="9" entrytime="00:02:05.45" />
                <RESULT eventid="99425" points="127" swimtime="00:00:50.16" resultid="107462" heatid="110825" lane="6" entrytime="00:00:49.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-01" firstname="Adrian" gender="M" lastname="Bilski" nation="POL" athleteid="107474">
              <RESULTS>
                <RESULT eventid="98798" points="226" reactiontime="+84" swimtime="00:00:33.22" resultid="107475" heatid="110599" lane="5" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="202" reactiontime="+87" swimtime="00:01:16.47" resultid="107476" heatid="110681" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.00" />
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="75" swimtime="00:00:55.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="135" reactiontime="+99" swimtime="00:01:38.64" resultid="107477" heatid="110697" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.43" />
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="75" swimtime="00:01:17.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="127" reactiontime="+91" swimtime="00:01:50.42" resultid="107478" heatid="110726" lane="5">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.02" />
                    <SPLIT distance="50" swimtime="00:00:53.61" />
                    <SPLIT distance="75" swimtime="00:01:21.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="168" reactiontime="+101" swimtime="00:02:59.80" resultid="107479" heatid="110771" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.63" />
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="75" swimtime="00:01:03.69" />
                    <SPLIT distance="100" swimtime="00:01:26.93" />
                    <SPLIT distance="125" swimtime="00:01:50.47" />
                    <SPLIT distance="150" swimtime="00:02:14.04" />
                    <SPLIT distance="175" swimtime="00:02:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="165" reactiontime="+111" swimtime="00:06:26.88" resultid="107480" heatid="110850" lane="1" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.30" />
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="75" swimtime="00:01:05.20" />
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                    <SPLIT distance="125" swimtime="00:01:51.82" />
                    <SPLIT distance="150" swimtime="00:02:15.76" />
                    <SPLIT distance="175" swimtime="00:02:40.63" />
                    <SPLIT distance="200" swimtime="00:03:05.19" />
                    <SPLIT distance="225" swimtime="00:03:29.35" />
                    <SPLIT distance="250" swimtime="00:03:54.31" />
                    <SPLIT distance="275" swimtime="00:04:19.46" />
                    <SPLIT distance="300" swimtime="00:04:44.14" />
                    <SPLIT distance="325" swimtime="00:05:09.17" />
                    <SPLIT distance="350" swimtime="00:05:32.76" />
                    <SPLIT distance="375" swimtime="00:06:02.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-16" firstname="Maciej" gender="M" lastname="Kujawa" nation="POL" athleteid="107496">
              <RESULTS>
                <RESULT eventid="98798" points="222" reactiontime="+90" swimtime="00:00:33.45" resultid="107497" heatid="110601" lane="0" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="217" swimtime="00:01:24.21" resultid="107498" heatid="110699" lane="9" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.39" />
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="75" swimtime="00:01:03.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="225" reactiontime="+94" swimtime="00:01:31.37" resultid="107499" heatid="110730" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.42" />
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                    <SPLIT distance="75" swimtime="00:01:06.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="239" reactiontime="+99" swimtime="00:00:40.68" resultid="107500" heatid="110827" lane="4" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="107508">
              <RESULTS>
                <RESULT eventid="106256" points="436" reactiontime="+100" swimtime="00:18:37.87" resultid="107509" heatid="110641" lane="1" entrytime="00:19:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.65" />
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="75" swimtime="00:00:48.66" />
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                    <SPLIT distance="125" swimtime="00:01:24.64" />
                    <SPLIT distance="150" swimtime="00:01:42.89" />
                    <SPLIT distance="175" swimtime="00:02:01.11" />
                    <SPLIT distance="200" swimtime="00:02:19.67" />
                    <SPLIT distance="225" swimtime="00:02:38.02" />
                    <SPLIT distance="250" swimtime="00:02:56.62" />
                    <SPLIT distance="275" swimtime="00:03:15.06" />
                    <SPLIT distance="300" swimtime="00:03:33.52" />
                    <SPLIT distance="325" swimtime="00:03:52.08" />
                    <SPLIT distance="350" swimtime="00:04:10.87" />
                    <SPLIT distance="375" swimtime="00:04:29.53" />
                    <SPLIT distance="400" swimtime="00:04:48.08" />
                    <SPLIT distance="425" swimtime="00:05:06.64" />
                    <SPLIT distance="450" swimtime="00:05:25.27" />
                    <SPLIT distance="475" swimtime="00:05:44.17" />
                    <SPLIT distance="500" swimtime="00:06:02.92" />
                    <SPLIT distance="525" swimtime="00:06:21.81" />
                    <SPLIT distance="550" swimtime="00:06:40.71" />
                    <SPLIT distance="575" swimtime="00:06:59.73" />
                    <SPLIT distance="600" swimtime="00:07:18.73" />
                    <SPLIT distance="625" swimtime="00:07:37.81" />
                    <SPLIT distance="650" swimtime="00:07:56.78" />
                    <SPLIT distance="675" swimtime="00:08:15.72" />
                    <SPLIT distance="700" swimtime="00:08:34.59" />
                    <SPLIT distance="725" swimtime="00:08:53.44" />
                    <SPLIT distance="750" swimtime="00:09:12.35" />
                    <SPLIT distance="775" swimtime="00:09:31.38" />
                    <SPLIT distance="800" swimtime="00:09:50.39" />
                    <SPLIT distance="825" swimtime="00:10:09.48" />
                    <SPLIT distance="850" swimtime="00:10:28.41" />
                    <SPLIT distance="875" swimtime="00:10:47.27" />
                    <SPLIT distance="900" swimtime="00:11:06.23" />
                    <SPLIT distance="925" swimtime="00:11:25.04" />
                    <SPLIT distance="950" swimtime="00:11:43.98" />
                    <SPLIT distance="975" swimtime="00:12:02.98" />
                    <SPLIT distance="1000" swimtime="00:12:22.32" />
                    <SPLIT distance="1025" swimtime="00:12:41.54" />
                    <SPLIT distance="1050" swimtime="00:13:00.92" />
                    <SPLIT distance="1075" swimtime="00:13:20.37" />
                    <SPLIT distance="1100" swimtime="00:13:39.39" />
                    <SPLIT distance="1125" swimtime="00:13:57.83" />
                    <SPLIT distance="1150" swimtime="00:14:16.95" />
                    <SPLIT distance="1175" swimtime="00:14:35.98" />
                    <SPLIT distance="1200" swimtime="00:14:55.17" />
                    <SPLIT distance="1225" swimtime="00:15:14.34" />
                    <SPLIT distance="1250" swimtime="00:15:33.59" />
                    <SPLIT distance="1275" swimtime="00:15:52.68" />
                    <SPLIT distance="1300" swimtime="00:16:11.70" />
                    <SPLIT distance="1325" swimtime="00:16:30.82" />
                    <SPLIT distance="1350" swimtime="00:16:49.69" />
                    <SPLIT distance="1375" swimtime="00:17:08.17" />
                    <SPLIT distance="1400" swimtime="00:17:27.12" />
                    <SPLIT distance="1425" swimtime="00:17:45.27" />
                    <SPLIT distance="1450" swimtime="00:18:03.53" />
                    <SPLIT distance="1475" swimtime="00:18:21.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="401" reactiontime="+95" swimtime="00:02:43.26" resultid="107510" heatid="110670" lane="1" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.38" />
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="75" swimtime="00:00:56.74" />
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                    <SPLIT distance="125" swimtime="00:01:39.18" />
                    <SPLIT distance="150" swimtime="00:02:00.72" />
                    <SPLIT distance="175" swimtime="00:02:22.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="500" reactiontime="+88" swimtime="00:01:10.02" resultid="107511" heatid="110734" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.27" />
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="75" swimtime="00:00:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="487" reactiontime="+83" swimtime="00:02:06.24" resultid="107512" heatid="110777" lane="7" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.98" />
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                    <SPLIT distance="75" swimtime="00:00:45.40" />
                    <SPLIT distance="100" swimtime="00:01:01.38" />
                    <SPLIT distance="125" swimtime="00:01:17.79" />
                    <SPLIT distance="150" swimtime="00:01:34.43" />
                    <SPLIT distance="175" swimtime="00:01:51.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="481" swimtime="00:00:32.21" resultid="107513" heatid="110834" lane="0" entrytime="00:00:32.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="458" reactiontime="+90" swimtime="00:04:35.21" resultid="107514" heatid="110845" lane="4" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.41" />
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                    <SPLIT distance="75" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:03.85" />
                    <SPLIT distance="125" swimtime="00:01:20.98" />
                    <SPLIT distance="150" swimtime="00:01:38.33" />
                    <SPLIT distance="175" swimtime="00:01:55.98" />
                    <SPLIT distance="200" swimtime="00:02:13.72" />
                    <SPLIT distance="225" swimtime="00:02:31.39" />
                    <SPLIT distance="250" swimtime="00:02:49.47" />
                    <SPLIT distance="275" swimtime="00:03:07.85" />
                    <SPLIT distance="300" swimtime="00:03:26.00" />
                    <SPLIT distance="325" swimtime="00:03:43.90" />
                    <SPLIT distance="350" swimtime="00:04:01.90" />
                    <SPLIT distance="375" swimtime="00:04:19.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-02" firstname="Marcin" gender="M" lastname="Stasiak" nation="POL" athleteid="107435">
              <RESULTS>
                <RESULT eventid="98798" points="319" reactiontime="+77" swimtime="00:00:29.64" resultid="107436" heatid="110605" lane="2" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="317" swimtime="00:01:14.26" resultid="107437" heatid="110701" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.32" />
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="75" swimtime="00:00:55.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="333" reactiontime="+88" swimtime="00:00:36.40" resultid="107438" heatid="110827" lane="3" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="Osóbka" nation="POL" athleteid="107453">
              <RESULTS>
                <RESULT eventid="98798" points="28" reactiontime="+98" swimtime="00:01:05.98" resultid="107454" heatid="110595" lane="7" entrytime="00:01:03.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="15" swimtime="00:01:41.82" resultid="107455" heatid="110825" lane="9" entrytime="00:00:59.03">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:46.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-06-29" firstname="Lucyna" gender="F" lastname="Serożyńska" nation="POL" athleteid="107468">
              <RESULTS>
                <RESULT eventid="98777" points="111" reactiontime="+110" swimtime="00:00:48.28" resultid="107469" heatid="110586" lane="6" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="60" reactiontime="+100" swimtime="00:01:05.40" resultid="107470" heatid="110646" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="130" reactiontime="+127" swimtime="00:02:02.96" resultid="107471" heatid="110721" lane="3" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.98" />
                    <SPLIT distance="50" swimtime="00:00:57.70" />
                    <SPLIT distance="75" swimtime="00:01:29.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="54" reactiontime="+89" swimtime="00:02:25.49" resultid="107472" heatid="110753" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.43" />
                    <SPLIT distance="50" swimtime="00:01:11.77" />
                    <SPLIT distance="75" swimtime="00:01:50.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="115" swimtime="00:00:59.09" resultid="107473" heatid="110818" lane="9" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="69" swimtime="00:03:20.51" resultid="107520" heatid="110781" lane="6">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.66" />
                    <SPLIT distance="50" swimtime="00:00:48.87" />
                    <SPLIT distance="75" swimtime="00:01:15.17" />
                    <SPLIT distance="100" swimtime="00:01:51.11" />
                    <SPLIT distance="125" swimtime="00:02:13.41" />
                    <SPLIT distance="150" swimtime="00:02:38.76" />
                    <SPLIT distance="175" swimtime="00:02:57.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107456" number="1" />
                    <RELAYPOSITION athleteid="107453" number="2" />
                    <RELAYPOSITION athleteid="107439" number="3" reactiontime="+85" />
                    <RELAYPOSITION athleteid="107447" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99059" points="46" reactiontime="+65" swimtime="00:04:11.62" resultid="107521" heatid="110716" lane="6">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.63" />
                    <SPLIT distance="50" swimtime="00:00:54.17" />
                    <SPLIT distance="75" swimtime="00:01:33.67" />
                    <SPLIT distance="100" swimtime="00:02:11.60" />
                    <SPLIT distance="125" swimtime="00:02:53.31" />
                    <SPLIT distance="150" swimtime="00:03:30.17" />
                    <SPLIT distance="175" swimtime="00:03:48.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107456" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="107453" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="107439" number="3" />
                    <RELAYPOSITION athleteid="107447" number="4" reactiontime="+89" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="99250" points="322" swimtime="00:02:00.44" resultid="107524" heatid="110783" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.18" />
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="75" swimtime="00:00:48.36" />
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                    <SPLIT distance="125" swimtime="00:01:19.70" />
                    <SPLIT distance="150" swimtime="00:01:34.15" />
                    <SPLIT distance="175" swimtime="00:01:46.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107489" number="1" />
                    <RELAYPOSITION athleteid="107496" number="2" />
                    <RELAYPOSITION athleteid="107501" number="3" />
                    <RELAYPOSITION athleteid="107508" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99059" points="271" reactiontime="+85" swimtime="00:02:19.82" resultid="107525" heatid="110717" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.27" />
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                    <SPLIT distance="75" swimtime="00:00:58.26" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="125" swimtime="00:01:32.62" />
                    <SPLIT distance="150" swimtime="00:01:52.57" />
                    <SPLIT distance="175" swimtime="00:02:05.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107496" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="107508" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="107489" number="3" />
                    <RELAYPOSITION athleteid="107501" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="318" reactiontime="+88" swimtime="00:02:00.89" resultid="107522" heatid="110631" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="75" swimtime="00:00:48.41" />
                    <SPLIT distance="100" swimtime="00:01:08.14" />
                    <SPLIT distance="125" swimtime="00:01:21.11" />
                    <SPLIT distance="150" swimtime="00:01:35.05" />
                    <SPLIT distance="175" swimtime="00:01:47.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107481" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="107463" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="107501" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="107508" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="295" reactiontime="+92" swimtime="00:02:15.89" resultid="107523" heatid="110837" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.35" />
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                    <SPLIT distance="75" swimtime="00:00:58.21" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="125" swimtime="00:01:30.28" />
                    <SPLIT distance="150" swimtime="00:01:48.46" />
                    <SPLIT distance="175" swimtime="00:02:01.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107463" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="107508" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="107481" number="3" />
                    <RELAYPOSITION athleteid="107501" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="110021" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1964-01-01" firstname="Joanna" gender="F" lastname="Bartosiewicz" nation="POL" athleteid="110101">
              <RESULTS>
                <RESULT eventid="98814" status="WDR" swimtime="00:00:00.00" resultid="110102" entrytime="00:03:10.00" />
                <RESULT eventid="98940" points="333" reactiontime="+97" swimtime="00:03:13.99" resultid="110103" heatid="110663" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.82" />
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                    <SPLIT distance="75" swimtime="00:01:09.55" />
                    <SPLIT distance="100" swimtime="00:01:34.53" />
                    <SPLIT distance="125" swimtime="00:01:59.18" />
                    <SPLIT distance="150" swimtime="00:02:24.27" />
                    <SPLIT distance="175" swimtime="00:02:49.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="313" reactiontime="+103" swimtime="00:01:23.40" resultid="110104" heatid="110692" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.32" />
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="75" swimtime="00:01:03.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="346" reactiontime="+76" swimtime="00:01:28.81" resultid="110105" heatid="110722" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.88" />
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                    <SPLIT distance="75" swimtime="00:01:05.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="329" swimtime="00:00:35.29" resultid="110106" heatid="110736" lane="3" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="305" reactiontime="+89" swimtime="00:01:21.08" resultid="110107" heatid="110794" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.88" />
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="75" swimtime="00:01:00.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="332" reactiontime="+91" swimtime="00:00:41.57" resultid="110108" heatid="110819" lane="8" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="110053">
              <RESULTS>
                <RESULT eventid="98798" points="158" reactiontime="+99" swimtime="00:00:37.47" resultid="110054" heatid="110597" lane="7" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="122" reactiontime="+103" swimtime="00:03:40.68" resultid="110055" heatid="110620" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.66" />
                    <SPLIT distance="50" swimtime="00:00:53.66" />
                    <SPLIT distance="75" swimtime="00:01:21.02" />
                    <SPLIT distance="100" swimtime="00:01:49.42" />
                    <SPLIT distance="125" swimtime="00:02:20.92" />
                    <SPLIT distance="150" swimtime="00:02:53.10" />
                    <SPLIT distance="175" swimtime="00:03:17.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="120" reactiontime="+90" swimtime="00:00:44.93" resultid="110056" heatid="110653" lane="2" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="138" reactiontime="+120" swimtime="00:01:26.87" resultid="110057" heatid="110679" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.71" />
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                    <SPLIT distance="75" swimtime="00:01:03.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="112" reactiontime="+81" swimtime="00:01:41.48" resultid="110058" heatid="110758" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.67" />
                    <SPLIT distance="50" swimtime="00:00:48.62" />
                    <SPLIT distance="75" swimtime="00:01:15.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="101" reactiontime="+91" swimtime="00:03:46.11" resultid="110059" heatid="110811" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.09" />
                    <SPLIT distance="50" swimtime="00:00:51.82" />
                    <SPLIT distance="75" swimtime="00:01:20.29" />
                    <SPLIT distance="100" swimtime="00:01:49.66" />
                    <SPLIT distance="125" swimtime="00:02:19.31" />
                    <SPLIT distance="150" swimtime="00:02:49.01" />
                    <SPLIT distance="175" swimtime="00:03:17.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="147" reactiontime="+103" swimtime="00:00:47.76" resultid="110060" heatid="110825" lane="7" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="110084">
              <RESULTS>
                <RESULT eventid="98798" status="WDR" swimtime="00:00:00.00" resultid="110085" entrytime="00:00:28.50" />
                <RESULT eventid="98956" points="262" reactiontime="+85" swimtime="00:03:08.13" resultid="110086" heatid="110668" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.69" />
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="75" swimtime="00:01:04.14" />
                    <SPLIT distance="100" swimtime="00:01:28.67" />
                    <SPLIT distance="125" swimtime="00:01:53.96" />
                    <SPLIT distance="150" swimtime="00:02:20.10" />
                    <SPLIT distance="175" swimtime="00:02:44.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="237" swimtime="00:01:21.80" resultid="110087" heatid="110701" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.05" />
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="75" swimtime="00:01:02.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="314" swimtime="00:01:21.79" resultid="110088" heatid="110732" lane="9" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.42" />
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="75" swimtime="00:00:59.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="268" swimtime="00:02:34.09" resultid="110089" heatid="110775" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.73" />
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="75" swimtime="00:00:52.96" />
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="125" swimtime="00:01:32.84" />
                    <SPLIT distance="150" swimtime="00:01:53.96" />
                    <SPLIT distance="175" swimtime="00:02:14.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="197" reactiontime="+77" swimtime="00:01:23.12" resultid="110090" heatid="110801" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.12" />
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="75" swimtime="00:01:01.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="343" reactiontime="+85" swimtime="00:00:36.05" resultid="110091" heatid="110830" lane="3" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="110066">
              <RESULTS>
                <RESULT eventid="98830" points="197" reactiontime="+110" swimtime="00:03:08.32" resultid="110067" heatid="110622" lane="1" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.52" />
                    <SPLIT distance="50" swimtime="00:00:46.32" />
                    <SPLIT distance="75" swimtime="00:01:10.20" />
                    <SPLIT distance="100" swimtime="00:01:32.65" />
                    <SPLIT distance="125" swimtime="00:01:58.84" />
                    <SPLIT distance="150" swimtime="00:02:25.27" />
                    <SPLIT distance="175" swimtime="00:02:47.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="204" reactiontime="+103" swimtime="00:12:32.27" resultid="110068" heatid="110637" lane="7" entrytime="00:12:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.53" />
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="75" swimtime="00:01:04.76" />
                    <SPLIT distance="100" swimtime="00:01:27.75" />
                    <SPLIT distance="125" swimtime="00:01:51.75" />
                    <SPLIT distance="150" swimtime="00:02:15.43" />
                    <SPLIT distance="175" swimtime="00:02:39.04" />
                    <SPLIT distance="200" swimtime="00:03:02.99" />
                    <SPLIT distance="225" swimtime="00:03:26.70" />
                    <SPLIT distance="250" swimtime="00:03:50.52" />
                    <SPLIT distance="275" swimtime="00:04:14.44" />
                    <SPLIT distance="300" swimtime="00:04:38.59" />
                    <SPLIT distance="325" swimtime="00:05:02.80" />
                    <SPLIT distance="350" swimtime="00:05:26.85" />
                    <SPLIT distance="375" swimtime="00:05:50.80" />
                    <SPLIT distance="400" swimtime="00:06:14.86" />
                    <SPLIT distance="425" swimtime="00:06:38.84" />
                    <SPLIT distance="450" swimtime="00:07:03.10" />
                    <SPLIT distance="475" swimtime="00:07:27.08" />
                    <SPLIT distance="500" swimtime="00:07:51.15" />
                    <SPLIT distance="525" swimtime="00:08:14.90" />
                    <SPLIT distance="550" swimtime="00:08:38.87" />
                    <SPLIT distance="575" swimtime="00:09:02.54" />
                    <SPLIT distance="600" swimtime="00:09:26.40" />
                    <SPLIT distance="625" swimtime="00:09:49.92" />
                    <SPLIT distance="650" swimtime="00:10:13.61" />
                    <SPLIT distance="675" swimtime="00:10:37.34" />
                    <SPLIT distance="700" swimtime="00:11:00.88" />
                    <SPLIT distance="725" swimtime="00:11:23.97" />
                    <SPLIT distance="750" swimtime="00:11:47.16" />
                    <SPLIT distance="775" swimtime="00:12:10.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="156" reactiontime="+84" swimtime="00:00:41.22" resultid="110069" heatid="110654" lane="7" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="199" reactiontime="+79" swimtime="00:01:26.64" resultid="110070" heatid="110698" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.68" />
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="75" swimtime="00:01:06.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="174" reactiontime="+78" swimtime="00:01:27.48" resultid="110071" heatid="110759" lane="5" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.81" />
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="75" swimtime="00:01:05.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="195" reactiontime="+113" swimtime="00:06:45.45" resultid="110072" heatid="110789" lane="3" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.45" />
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                    <SPLIT distance="75" swimtime="00:01:17.67" />
                    <SPLIT distance="100" swimtime="00:01:46.61" />
                    <SPLIT distance="125" swimtime="00:02:10.75" />
                    <SPLIT distance="150" swimtime="00:02:34.55" />
                    <SPLIT distance="175" swimtime="00:02:59.15" />
                    <SPLIT distance="200" swimtime="00:03:23.75" />
                    <SPLIT distance="225" swimtime="00:03:50.94" />
                    <SPLIT distance="250" swimtime="00:04:18.56" />
                    <SPLIT distance="275" swimtime="00:04:46.27" />
                    <SPLIT distance="300" swimtime="00:05:13.92" />
                    <SPLIT distance="325" swimtime="00:05:37.23" />
                    <SPLIT distance="350" swimtime="00:06:00.00" />
                    <SPLIT distance="375" swimtime="00:06:22.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="166" reactiontime="+91" swimtime="00:03:12.14" resultid="110073" heatid="110813" lane="0" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.88" />
                    <SPLIT distance="50" swimtime="00:00:44.61" />
                    <SPLIT distance="75" swimtime="00:01:07.95" />
                    <SPLIT distance="100" swimtime="00:01:32.34" />
                    <SPLIT distance="125" swimtime="00:01:57.58" />
                    <SPLIT distance="150" swimtime="00:02:22.73" />
                    <SPLIT distance="175" swimtime="00:02:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="179" reactiontime="+94" swimtime="00:06:16.12" resultid="110074" heatid="110849" lane="7" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.80" />
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="75" swimtime="00:01:04.42" />
                    <SPLIT distance="100" swimtime="00:01:28.33" />
                    <SPLIT distance="125" swimtime="00:01:52.19" />
                    <SPLIT distance="150" swimtime="00:02:16.12" />
                    <SPLIT distance="175" swimtime="00:02:40.36" />
                    <SPLIT distance="200" swimtime="00:03:04.34" />
                    <SPLIT distance="225" swimtime="00:03:28.25" />
                    <SPLIT distance="250" swimtime="00:03:52.40" />
                    <SPLIT distance="275" swimtime="00:04:16.80" />
                    <SPLIT distance="300" swimtime="00:04:41.22" />
                    <SPLIT distance="325" swimtime="00:05:05.53" />
                    <SPLIT distance="350" swimtime="00:05:29.76" />
                    <SPLIT distance="375" swimtime="00:05:53.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="110092">
              <RESULTS>
                <RESULT eventid="98777" points="205" reactiontime="+97" swimtime="00:00:39.41" resultid="110093" heatid="110588" lane="7" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="124" reactiontime="+106" swimtime="00:04:03.87" resultid="110094" heatid="110614" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.00" />
                    <SPLIT distance="50" swimtime="00:00:54.13" />
                    <SPLIT distance="75" swimtime="00:01:25.96" />
                    <SPLIT distance="100" swimtime="00:01:56.62" />
                    <SPLIT distance="125" swimtime="00:02:32.46" />
                    <SPLIT distance="150" swimtime="00:03:07.88" />
                    <SPLIT distance="175" swimtime="00:03:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="128" reactiontime="+55" swimtime="00:00:50.86" resultid="110095" heatid="110647" lane="8" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="76" reactiontime="+109" swimtime="00:04:41.36" resultid="110096" heatid="110707" lane="6" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.40" />
                    <SPLIT distance="50" swimtime="00:01:00.08" />
                    <SPLIT distance="75" swimtime="00:01:35.24" />
                    <SPLIT distance="100" swimtime="00:02:11.22" />
                    <SPLIT distance="125" swimtime="00:02:49.32" />
                    <SPLIT distance="150" swimtime="00:03:27.41" />
                    <SPLIT distance="175" swimtime="00:04:06.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="127" swimtime="00:00:48.46" resultid="110097" heatid="110736" lane="6" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="129" swimtime="00:08:33.50" resultid="110098" heatid="110786" lane="9" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.00" />
                    <SPLIT distance="50" swimtime="00:01:00.99" />
                    <SPLIT distance="75" swimtime="00:01:36.67" />
                    <SPLIT distance="100" swimtime="00:02:12.62" />
                    <SPLIT distance="125" swimtime="00:02:48.49" />
                    <SPLIT distance="150" swimtime="00:03:22.39" />
                    <SPLIT distance="175" swimtime="00:03:55.92" />
                    <SPLIT distance="200" swimtime="00:04:29.67" />
                    <SPLIT distance="225" swimtime="00:05:04.55" />
                    <SPLIT distance="250" swimtime="00:05:39.27" />
                    <SPLIT distance="275" swimtime="00:06:13.86" />
                    <SPLIT distance="300" swimtime="00:06:50.23" />
                    <SPLIT distance="325" swimtime="00:07:17.09" />
                    <SPLIT distance="350" swimtime="00:07:44.21" />
                    <SPLIT distance="375" swimtime="00:08:09.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="87" swimtime="00:02:02.84" resultid="110099" heatid="110794" lane="9" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.17" />
                    <SPLIT distance="50" swimtime="00:00:55.75" />
                    <SPLIT distance="75" swimtime="00:01:30.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="160" swimtime="00:07:11.42" resultid="110100" heatid="110842" lane="6" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.50" />
                    <SPLIT distance="50" swimtime="00:00:47.39" />
                    <SPLIT distance="75" swimtime="00:01:15.48" />
                    <SPLIT distance="100" swimtime="00:01:45.44" />
                    <SPLIT distance="125" swimtime="00:02:15.00" />
                    <SPLIT distance="150" swimtime="00:02:42.95" />
                    <SPLIT distance="175" swimtime="00:03:10.82" />
                    <SPLIT distance="200" swimtime="00:03:38.31" />
                    <SPLIT distance="225" swimtime="00:04:05.87" />
                    <SPLIT distance="250" swimtime="00:04:32.96" />
                    <SPLIT distance="275" swimtime="00:05:00.48" />
                    <SPLIT distance="300" swimtime="00:05:27.93" />
                    <SPLIT distance="325" swimtime="00:05:54.97" />
                    <SPLIT distance="350" swimtime="00:06:22.36" />
                    <SPLIT distance="375" swimtime="00:06:48.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" athleteid="110075">
              <RESULTS>
                <RESULT eventid="98798" points="254" reactiontime="+76" swimtime="00:00:31.99" resultid="110076" heatid="110600" lane="8" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="220" swimtime="00:03:01.49" resultid="110077" heatid="110621" lane="4" entrytime="00:03:10.41">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.83" />
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                    <SPLIT distance="75" swimtime="00:00:59.42" />
                    <SPLIT distance="100" swimtime="00:01:24.01" />
                    <SPLIT distance="125" swimtime="00:01:50.30" />
                    <SPLIT distance="150" swimtime="00:02:16.92" />
                    <SPLIT distance="175" swimtime="00:02:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="227" reactiontime="+90" swimtime="00:03:17.44" resultid="110078" heatid="110667" lane="1" entrytime="00:03:20.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.20" />
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                    <SPLIT distance="75" swimtime="00:01:06.58" />
                    <SPLIT distance="100" swimtime="00:01:32.07" />
                    <SPLIT distance="125" swimtime="00:01:57.87" />
                    <SPLIT distance="150" swimtime="00:02:24.65" />
                    <SPLIT distance="175" swimtime="00:02:51.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="124" swimtime="00:03:37.61" resultid="110079" heatid="110710" lane="4" entrytime="00:03:53.51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.70" />
                    <SPLIT distance="50" swimtime="00:00:46.99" />
                    <SPLIT distance="75" swimtime="00:01:14.49" />
                    <SPLIT distance="100" swimtime="00:01:42.77" />
                    <SPLIT distance="125" swimtime="00:02:11.38" />
                    <SPLIT distance="150" swimtime="00:02:40.74" />
                    <SPLIT distance="175" swimtime="00:03:11.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="243" swimtime="00:01:29.02" resultid="110080" heatid="110729" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.79" />
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="75" swimtime="00:01:04.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="223" reactiontime="+86" swimtime="00:00:35.91" resultid="110081" heatid="110744" lane="1" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="142" swimtime="00:01:32.77" resultid="110082" heatid="110800" lane="9" entrytime="00:01:32.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="75" swimtime="00:01:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="255" swimtime="00:00:39.78" resultid="110083" heatid="110828" lane="0" entrytime="00:00:39.95">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="110061">
              <RESULTS>
                <RESULT eventid="98891" points="120" reactiontime="+106" swimtime="00:14:57.87" resultid="110062" heatid="110638" lane="6" entrytime="00:15:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.09" />
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                    <SPLIT distance="75" swimtime="00:01:15.26" />
                    <SPLIT distance="100" swimtime="00:01:43.74" />
                    <SPLIT distance="125" swimtime="00:02:12.01" />
                    <SPLIT distance="150" swimtime="00:02:40.17" />
                    <SPLIT distance="175" swimtime="00:03:07.60" />
                    <SPLIT distance="200" swimtime="00:03:35.97" />
                    <SPLIT distance="225" swimtime="00:04:03.90" />
                    <SPLIT distance="250" swimtime="00:04:32.94" />
                    <SPLIT distance="275" swimtime="00:05:01.30" />
                    <SPLIT distance="300" swimtime="00:05:30.51" />
                    <SPLIT distance="325" swimtime="00:05:58.46" />
                    <SPLIT distance="350" swimtime="00:06:27.47" />
                    <SPLIT distance="375" swimtime="00:06:55.80" />
                    <SPLIT distance="400" swimtime="00:07:24.07" />
                    <SPLIT distance="425" swimtime="00:07:51.88" />
                    <SPLIT distance="450" swimtime="00:08:21.06" />
                    <SPLIT distance="475" swimtime="00:08:49.53" />
                    <SPLIT distance="500" swimtime="00:09:18.20" />
                    <SPLIT distance="525" swimtime="00:09:46.61" />
                    <SPLIT distance="550" swimtime="00:10:15.44" />
                    <SPLIT distance="575" swimtime="00:10:42.88" />
                    <SPLIT distance="600" swimtime="00:11:12.40" />
                    <SPLIT distance="625" swimtime="00:11:40.45" />
                    <SPLIT distance="650" swimtime="00:12:09.36" />
                    <SPLIT distance="675" swimtime="00:12:38.65" />
                    <SPLIT distance="700" swimtime="00:13:07.97" />
                    <SPLIT distance="725" swimtime="00:13:36.73" />
                    <SPLIT distance="750" swimtime="00:14:05.49" />
                    <SPLIT distance="775" swimtime="00:14:32.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="125" swimtime="00:00:44.40" resultid="110063" heatid="110653" lane="6" entrytime="00:00:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="108" reactiontime="+84" swimtime="00:01:42.68" resultid="110064" heatid="110759" lane="9" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.73" />
                    <SPLIT distance="50" swimtime="00:00:50.87" />
                    <SPLIT distance="75" swimtime="00:01:17.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="100" reactiontime="+105" swimtime="00:03:46.87" resultid="110065" heatid="110811" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.51" />
                    <SPLIT distance="50" swimtime="00:00:53.55" />
                    <SPLIT distance="75" swimtime="00:01:21.93" />
                    <SPLIT distance="100" swimtime="00:01:51.47" />
                    <SPLIT distance="125" swimtime="00:02:21.25" />
                    <SPLIT distance="150" swimtime="00:02:51.01" />
                    <SPLIT distance="175" swimtime="00:03:20.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="212" reactiontime="+80" swimtime="00:02:31.68" resultid="110111" heatid="110717" lane="8" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.24" />
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                    <SPLIT distance="75" swimtime="00:01:02.65" />
                    <SPLIT distance="100" swimtime="00:01:22.34" />
                    <SPLIT distance="125" swimtime="00:01:38.18" />
                    <SPLIT distance="150" swimtime="00:01:57.65" />
                    <SPLIT distance="175" swimtime="00:02:13.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110061" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="110084" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="110075" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="110066" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="231" reactiontime="+77" swimtime="00:02:14.61" resultid="110112" heatid="110782" lane="7" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="75" swimtime="00:00:48.43" />
                    <SPLIT distance="100" swimtime="00:01:07.64" />
                    <SPLIT distance="125" swimtime="00:01:23.89" />
                    <SPLIT distance="150" swimtime="00:01:42.11" />
                    <SPLIT distance="175" swimtime="00:01:57.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110084" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="110061" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="110066" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="110075" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" status="WDR" swimtime="00:00:00.00" resultid="110109" entrytime="00:02:15.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110084" number="1" />
                    <RELAYPOSITION athleteid="110092" number="2" />
                    <RELAYPOSITION athleteid="110101" number="3" />
                    <RELAYPOSITION athleteid="110075" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" status="WDR" swimtime="00:00:00.00" resultid="110110" entrytime="00:02:32.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110101" number="1" />
                    <RELAYPOSITION athleteid="110075" number="2" />
                    <RELAYPOSITION athleteid="110084" number="3" />
                    <RELAYPOSITION athleteid="110092" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="100413" nation="POL" region="WAR" clubid="109053" name="UKP Jedynka Elbląg">
          <CONTACT city="Elbląg" name="Wysocki" phone="696427414" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1980-03-21" firstname="Tomasz" gender="M" lastname="Wysocki" nation="POL" athleteid="109054">
              <RESULTS>
                <RESULT eventid="98924" points="454" reactiontime="+79" swimtime="00:00:28.90" resultid="109055" heatid="110660" lane="8" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="RZ" clubid="107272" name="UKS Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1970-03-15" firstname="Witold" gender="M" lastname="Flak" nation="POL" athleteid="109008">
              <RESULTS>
                <RESULT eventid="98798" points="361" reactiontime="+86" swimtime="00:00:28.43" resultid="109009" heatid="110606" lane="8" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="225" reactiontime="+78" swimtime="00:00:36.48" resultid="109010" heatid="110655" lane="4" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="366" swimtime="00:01:10.81" resultid="109011" heatid="110702" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="75" swimtime="00:00:53.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="362" reactiontime="+85" swimtime="00:01:17.97" resultid="109012" heatid="110731" lane="7" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="75" swimtime="00:00:57.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="330" swimtime="00:00:31.52" resultid="109013" heatid="110747" lane="9" entrytime="00:00:31.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="371" swimtime="00:00:35.11" resultid="109014" heatid="110831" lane="0" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="108994">
              <RESULTS>
                <RESULT eventid="98798" points="319" reactiontime="+75" swimtime="00:00:29.65" resultid="108995" heatid="110604" lane="8" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="267" reactiontime="+89" swimtime="00:21:55.53" resultid="108996" heatid="110642" lane="1" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.58" />
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="75" swimtime="00:00:54.63" />
                    <SPLIT distance="100" swimtime="00:01:14.04" />
                    <SPLIT distance="125" swimtime="00:01:33.71" />
                    <SPLIT distance="150" swimtime="00:01:54.28" />
                    <SPLIT distance="175" swimtime="00:02:14.68" />
                    <SPLIT distance="200" swimtime="00:02:35.12" />
                    <SPLIT distance="225" swimtime="00:02:55.50" />
                    <SPLIT distance="250" swimtime="00:03:16.39" />
                    <SPLIT distance="275" swimtime="00:03:37.25" />
                    <SPLIT distance="300" swimtime="00:03:58.38" />
                    <SPLIT distance="325" swimtime="00:04:19.52" />
                    <SPLIT distance="350" swimtime="00:04:40.90" />
                    <SPLIT distance="375" swimtime="00:05:02.06" />
                    <SPLIT distance="400" swimtime="00:05:23.63" />
                    <SPLIT distance="425" swimtime="00:05:44.60" />
                    <SPLIT distance="450" swimtime="00:06:07.29" />
                    <SPLIT distance="475" swimtime="00:06:28.84" />
                    <SPLIT distance="500" swimtime="00:06:50.85" />
                    <SPLIT distance="525" swimtime="00:07:12.51" />
                    <SPLIT distance="550" swimtime="00:07:34.57" />
                    <SPLIT distance="575" swimtime="00:07:56.58" />
                    <SPLIT distance="600" swimtime="00:08:18.94" />
                    <SPLIT distance="625" swimtime="00:08:41.07" />
                    <SPLIT distance="650" swimtime="00:09:03.12" />
                    <SPLIT distance="675" swimtime="00:09:26.06" />
                    <SPLIT distance="700" swimtime="00:09:48.56" />
                    <SPLIT distance="725" swimtime="00:10:10.87" />
                    <SPLIT distance="750" swimtime="00:10:33.76" />
                    <SPLIT distance="775" swimtime="00:10:56.58" />
                    <SPLIT distance="800" swimtime="00:11:19.74" />
                    <SPLIT distance="825" swimtime="00:11:42.15" />
                    <SPLIT distance="850" swimtime="00:12:05.49" />
                    <SPLIT distance="875" swimtime="00:12:28.61" />
                    <SPLIT distance="900" swimtime="00:12:52.27" />
                    <SPLIT distance="925" swimtime="00:13:15.43" />
                    <SPLIT distance="950" swimtime="00:13:39.03" />
                    <SPLIT distance="975" swimtime="00:14:01.94" />
                    <SPLIT distance="1000" swimtime="00:14:25.34" />
                    <SPLIT distance="1025" swimtime="00:14:48.06" />
                    <SPLIT distance="1050" swimtime="00:15:11.40" />
                    <SPLIT distance="1075" swimtime="00:15:34.23" />
                    <SPLIT distance="1100" swimtime="00:15:57.61" />
                    <SPLIT distance="1125" swimtime="00:16:20.53" />
                    <SPLIT distance="1150" swimtime="00:16:43.73" />
                    <SPLIT distance="1175" swimtime="00:17:06.46" />
                    <SPLIT distance="1200" swimtime="00:17:29.85" />
                    <SPLIT distance="1225" swimtime="00:17:52.34" />
                    <SPLIT distance="1250" swimtime="00:18:15.48" />
                    <SPLIT distance="1275" swimtime="00:18:37.94" />
                    <SPLIT distance="1300" swimtime="00:19:00.71" />
                    <SPLIT distance="1325" swimtime="00:19:22.95" />
                    <SPLIT distance="1350" swimtime="00:19:45.38" />
                    <SPLIT distance="1375" swimtime="00:20:08.00" />
                    <SPLIT distance="1400" swimtime="00:20:30.42" />
                    <SPLIT distance="1425" swimtime="00:20:52.01" />
                    <SPLIT distance="1450" swimtime="00:21:13.89" />
                    <SPLIT distance="1475" swimtime="00:21:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="317" reactiontime="+55" swimtime="00:01:05.90" resultid="108997" heatid="110683" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="75" swimtime="00:00:49.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="203" reactiontime="+77" swimtime="00:03:04.47" resultid="108998" heatid="110711" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.42" />
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="75" swimtime="00:01:03.55" />
                    <SPLIT distance="100" swimtime="00:01:28.86" />
                    <SPLIT distance="125" swimtime="00:01:54.14" />
                    <SPLIT distance="150" swimtime="00:02:19.73" />
                    <SPLIT distance="175" swimtime="00:02:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="311" reactiontime="+65" swimtime="00:02:26.56" resultid="108999" heatid="110773" lane="7" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.68" />
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="75" swimtime="00:00:51.47" />
                    <SPLIT distance="100" swimtime="00:01:10.09" />
                    <SPLIT distance="125" swimtime="00:01:29.26" />
                    <SPLIT distance="150" swimtime="00:01:48.95" />
                    <SPLIT distance="175" swimtime="00:02:08.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="109000" heatid="110789" lane="5" entrytime="00:06:40.00" />
                <RESULT eventid="99473" points="308" reactiontime="+78" swimtime="00:05:14.13" resultid="109001" heatid="110847" lane="5" entrytime="00:05:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.54" />
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="75" swimtime="00:00:54.43" />
                    <SPLIT distance="100" swimtime="00:01:13.86" />
                    <SPLIT distance="125" swimtime="00:01:33.68" />
                    <SPLIT distance="150" swimtime="00:01:53.64" />
                    <SPLIT distance="175" swimtime="00:02:13.69" />
                    <SPLIT distance="200" swimtime="00:02:34.33" />
                    <SPLIT distance="225" swimtime="00:02:54.80" />
                    <SPLIT distance="250" swimtime="00:03:15.05" />
                    <SPLIT distance="275" swimtime="00:03:35.26" />
                    <SPLIT distance="300" swimtime="00:03:55.15" />
                    <SPLIT distance="325" swimtime="00:04:15.15" />
                    <SPLIT distance="350" swimtime="00:04:35.36" />
                    <SPLIT distance="375" swimtime="00:04:55.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-27" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="109002">
              <RESULTS>
                <RESULT eventid="106256" points="345" reactiontime="+82" swimtime="00:20:09.15" resultid="109003" heatid="110641" lane="2" entrytime="00:19:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.41" />
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="75" swimtime="00:00:51.09" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="125" swimtime="00:01:29.00" />
                    <SPLIT distance="150" swimtime="00:01:48.17" />
                    <SPLIT distance="175" swimtime="00:02:07.48" />
                    <SPLIT distance="200" swimtime="00:02:26.91" />
                    <SPLIT distance="225" swimtime="00:02:47.09" />
                    <SPLIT distance="250" swimtime="00:03:07.19" />
                    <SPLIT distance="275" swimtime="00:03:27.51" />
                    <SPLIT distance="300" swimtime="00:03:48.06" />
                    <SPLIT distance="325" swimtime="00:04:08.91" />
                    <SPLIT distance="350" swimtime="00:04:29.98" />
                    <SPLIT distance="375" swimtime="00:04:51.09" />
                    <SPLIT distance="400" swimtime="00:05:11.91" />
                    <SPLIT distance="425" swimtime="00:05:33.13" />
                    <SPLIT distance="450" swimtime="00:05:53.89" />
                    <SPLIT distance="475" swimtime="00:06:14.77" />
                    <SPLIT distance="500" swimtime="00:06:35.32" />
                    <SPLIT distance="525" swimtime="00:06:55.93" />
                    <SPLIT distance="550" swimtime="00:07:16.90" />
                    <SPLIT distance="575" swimtime="00:07:37.92" />
                    <SPLIT distance="600" swimtime="00:07:58.32" />
                    <SPLIT distance="625" swimtime="00:08:18.73" />
                    <SPLIT distance="650" swimtime="00:08:39.54" />
                    <SPLIT distance="675" swimtime="00:08:59.56" />
                    <SPLIT distance="700" swimtime="00:09:20.20" />
                    <SPLIT distance="725" swimtime="00:09:40.55" />
                    <SPLIT distance="750" swimtime="00:10:01.36" />
                    <SPLIT distance="775" swimtime="00:10:21.63" />
                    <SPLIT distance="800" swimtime="00:10:41.98" />
                    <SPLIT distance="825" swimtime="00:11:02.07" />
                    <SPLIT distance="850" swimtime="00:11:22.62" />
                    <SPLIT distance="875" swimtime="00:11:43.36" />
                    <SPLIT distance="900" swimtime="00:12:03.93" />
                    <SPLIT distance="925" swimtime="00:12:24.28" />
                    <SPLIT distance="950" swimtime="00:12:45.07" />
                    <SPLIT distance="975" swimtime="00:13:05.19" />
                    <SPLIT distance="1000" swimtime="00:13:25.71" />
                    <SPLIT distance="1025" swimtime="00:13:45.61" />
                    <SPLIT distance="1050" swimtime="00:14:05.64" />
                    <SPLIT distance="1075" swimtime="00:14:25.41" />
                    <SPLIT distance="1100" swimtime="00:14:45.48" />
                    <SPLIT distance="1125" swimtime="00:15:05.55" />
                    <SPLIT distance="1150" swimtime="00:15:25.61" />
                    <SPLIT distance="1175" swimtime="00:15:45.56" />
                    <SPLIT distance="1200" swimtime="00:16:06.11" />
                    <SPLIT distance="1225" swimtime="00:16:26.56" />
                    <SPLIT distance="1250" swimtime="00:16:47.25" />
                    <SPLIT distance="1275" swimtime="00:17:07.71" />
                    <SPLIT distance="1300" swimtime="00:17:28.06" />
                    <SPLIT distance="1325" swimtime="00:17:48.36" />
                    <SPLIT distance="1350" swimtime="00:18:08.97" />
                    <SPLIT distance="1375" swimtime="00:18:29.42" />
                    <SPLIT distance="1400" swimtime="00:18:50.16" />
                    <SPLIT distance="1425" swimtime="00:19:10.04" />
                    <SPLIT distance="1450" swimtime="00:19:30.18" />
                    <SPLIT distance="1475" swimtime="00:19:49.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="518" reactiontime="+65" swimtime="00:02:29.95" resultid="109004" heatid="110670" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.41" />
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="75" swimtime="00:00:52.81" />
                    <SPLIT distance="100" swimtime="00:01:11.65" />
                    <SPLIT distance="125" swimtime="00:01:31.03" />
                    <SPLIT distance="150" swimtime="00:01:50.46" />
                    <SPLIT distance="175" swimtime="00:02:10.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="477" reactiontime="+80" swimtime="00:01:11.14" resultid="109005" heatid="110734" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.16" />
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="75" swimtime="00:00:51.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="502" reactiontime="+62" swimtime="00:00:31.76" resultid="109006" heatid="110834" lane="5" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="109007" heatid="110845" lane="2" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="Szklarz" nation="POL" athleteid="108988">
              <RESULTS>
                <RESULT eventid="98798" points="360" reactiontime="+81" swimtime="00:00:28.46" resultid="108989" heatid="110606" lane="2" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="278" reactiontime="+68" swimtime="00:00:34.04" resultid="108990" heatid="110657" lane="7" entrytime="00:00:33.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="108991" heatid="110685" lane="3" entrytime="00:01:02.00" />
                <RESULT eventid="99170" points="349" reactiontime="+76" swimtime="00:00:30.94" resultid="108992" heatid="110747" lane="7" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="351" swimtime="00:00:35.78" resultid="108993" heatid="110831" lane="6" entrytime="00:00:35.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-17" firstname="Sławomir" gender="M" lastname="Kowalski" nation="POL" athleteid="108978">
              <RESULTS>
                <RESULT eventid="98798" points="383" reactiontime="+73" swimtime="00:00:27.89" resultid="108979" heatid="110599" lane="3" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="108980" heatid="110624" lane="6" entrytime="00:02:45.00" />
                <RESULT eventid="98956" points="319" swimtime="00:02:56.19" resultid="108981" heatid="110668" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.64" />
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="75" swimtime="00:00:56.86" />
                    <SPLIT distance="100" swimtime="00:01:19.05" />
                    <SPLIT distance="125" swimtime="00:01:42.50" />
                    <SPLIT distance="150" swimtime="00:02:06.84" />
                    <SPLIT distance="175" swimtime="00:02:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="343" swimtime="00:01:04.19" resultid="108982" heatid="110685" lane="0" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.95" />
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="75" swimtime="00:00:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="371" swimtime="00:01:17.39" resultid="108984" heatid="110733" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.73" />
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="75" swimtime="00:00:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="108985" heatid="110746" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="108986" heatid="110801" lane="5" entrytime="00:01:15.00" />
                <RESULT eventid="99425" points="403" swimtime="00:00:34.16" resultid="108987" heatid="110832" lane="0" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="108969">
              <RESULTS>
                <RESULT eventid="98798" points="480" reactiontime="+79" swimtime="00:00:25.86" resultid="108970" heatid="110606" lane="4" entrytime="00:00:28.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="399" reactiontime="+72" swimtime="00:02:28.83" resultid="108971" heatid="110625" lane="5" entrytime="00:02:36.36">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.53" />
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="75" swimtime="00:00:50.61" />
                    <SPLIT distance="100" swimtime="00:01:10.36" />
                    <SPLIT distance="125" swimtime="00:01:32.61" />
                    <SPLIT distance="150" swimtime="00:01:54.88" />
                    <SPLIT distance="175" swimtime="00:02:13.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="482" reactiontime="+81" swimtime="00:00:57.31" resultid="108972" heatid="110686" lane="7" entrytime="00:01:01.28">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.01" />
                    <SPLIT distance="50" swimtime="00:00:27.34" />
                    <SPLIT distance="75" swimtime="00:00:42.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="430" swimtime="00:01:07.07" resultid="108973" heatid="110704" lane="0" entrytime="00:01:08.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.39" />
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="75" swimtime="00:00:50.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="439" reactiontime="+78" swimtime="00:00:28.67" resultid="108974" heatid="110747" lane="8" entrytime="00:00:31.22">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="476" reactiontime="+86" swimtime="00:02:07.23" resultid="108975" heatid="110777" lane="8" entrytime="00:02:11.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.83" />
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="75" swimtime="00:00:45.19" />
                    <SPLIT distance="100" swimtime="00:01:01.39" />
                    <SPLIT distance="125" swimtime="00:01:17.63" />
                    <SPLIT distance="150" swimtime="00:01:34.54" />
                    <SPLIT distance="175" swimtime="00:01:51.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="409" reactiontime="+79" swimtime="00:01:05.24" resultid="108976" heatid="110802" lane="7" entrytime="00:01:12.38">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.80" />
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="75" swimtime="00:00:47.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="450" swimtime="00:00:32.94" resultid="108977" heatid="110832" lane="6" entrytime="00:00:34.68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-17" firstname="Tomasz" gender="M" lastname="Ostrowski" nation="POL" athleteid="109030">
              <RESULTS>
                <RESULT eventid="98798" points="500" reactiontime="+84" swimtime="00:00:25.51" resultid="109031" heatid="110610" lane="1" entrytime="00:00:26.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="493" reactiontime="+76" swimtime="00:00:56.88" resultid="109032" heatid="110687" lane="7" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.52" />
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                    <SPLIT distance="75" swimtime="00:00:41.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="455" reactiontime="+75" swimtime="00:01:05.83" resultid="109033" heatid="110704" lane="8" entrytime="00:01:08.09">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.74" />
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="75" swimtime="00:00:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="503" reactiontime="+78" swimtime="00:00:27.41" resultid="109034" heatid="110749" lane="3" entrytime="00:00:28.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="419" reactiontime="+87" swimtime="00:00:33.73" resultid="109035" heatid="110832" lane="1" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-14" firstname="Piotr" gender="M" lastname="Darowski" nation="POL" athleteid="109023">
              <RESULTS>
                <RESULT eventid="98830" points="417" reactiontime="+89" swimtime="00:02:26.67" resultid="109024" heatid="110626" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.58" />
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="75" swimtime="00:00:51.50" />
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                    <SPLIT distance="125" swimtime="00:01:30.79" />
                    <SPLIT distance="150" swimtime="00:01:51.51" />
                    <SPLIT distance="175" swimtime="00:02:09.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="455" reactiontime="+76" swimtime="00:02:36.62" resultid="109025" heatid="110670" lane="8" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.82" />
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="75" swimtime="00:00:53.21" />
                    <SPLIT distance="100" swimtime="00:01:13.12" />
                    <SPLIT distance="125" swimtime="00:01:33.21" />
                    <SPLIT distance="150" swimtime="00:01:54.12" />
                    <SPLIT distance="175" swimtime="00:02:15.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="451" reactiontime="+84" swimtime="00:01:12.49" resultid="109026" heatid="110733" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.60" />
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="75" swimtime="00:00:52.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="395" swimtime="00:05:20.73" resultid="109027" heatid="110791" lane="6" entrytime="00:05:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.32" />
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="75" swimtime="00:00:52.05" />
                    <SPLIT distance="100" swimtime="00:01:12.05" />
                    <SPLIT distance="125" swimtime="00:01:33.94" />
                    <SPLIT distance="150" swimtime="00:01:55.58" />
                    <SPLIT distance="175" swimtime="00:02:16.79" />
                    <SPLIT distance="200" swimtime="00:02:38.34" />
                    <SPLIT distance="225" swimtime="00:02:59.86" />
                    <SPLIT distance="250" swimtime="00:03:21.40" />
                    <SPLIT distance="275" swimtime="00:03:42.95" />
                    <SPLIT distance="300" swimtime="00:04:04.89" />
                    <SPLIT distance="325" swimtime="00:04:24.14" />
                    <SPLIT distance="350" swimtime="00:04:43.53" />
                    <SPLIT distance="375" swimtime="00:05:03.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="351" swimtime="00:01:08.65" resultid="109028" heatid="110803" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.47" />
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="75" swimtime="00:00:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="446" reactiontime="+69" swimtime="00:00:33.04" resultid="109029" heatid="110833" lane="7" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="109015">
              <RESULTS>
                <RESULT eventid="98814" points="338" reactiontime="+85" swimtime="00:02:54.87" resultid="109016" heatid="110617" lane="2" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.73" />
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="75" swimtime="00:00:59.07" />
                    <SPLIT distance="100" swimtime="00:01:20.97" />
                    <SPLIT distance="125" swimtime="00:01:46.63" />
                    <SPLIT distance="150" swimtime="00:02:13.26" />
                    <SPLIT distance="175" swimtime="00:02:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="341" swimtime="00:03:12.57" resultid="109017" heatid="110663" lane="6" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.88" />
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                    <SPLIT distance="75" swimtime="00:01:08.64" />
                    <SPLIT distance="100" swimtime="00:01:33.53" />
                    <SPLIT distance="125" swimtime="00:01:58.12" />
                    <SPLIT distance="150" swimtime="00:02:23.54" />
                    <SPLIT distance="175" swimtime="00:02:48.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="353" swimtime="00:01:20.11" resultid="109018" heatid="110694" lane="9" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.76" />
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="75" swimtime="00:01:01.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="352" swimtime="00:01:28.29" resultid="109019" heatid="110724" lane="9" entrytime="00:01:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.80" />
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="75" swimtime="00:01:05.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="285" swimtime="00:00:37.03" resultid="109020" heatid="110739" lane="0" entrytime="00:00:35.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="109021" heatid="110794" lane="5" entrytime="00:01:30.00" />
                <RESULT eventid="99409" points="346" reactiontime="+47" swimtime="00:00:41.00" resultid="109022" heatid="110821" lane="2" entrytime="00:00:40.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="108962">
              <RESULTS>
                <RESULT eventid="98777" points="378" reactiontime="+96" swimtime="00:00:32.12" resultid="108963" heatid="110591" lane="2" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="370" reactiontime="+83" swimtime="00:01:10.90" resultid="108964" heatid="110675" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.91" />
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="75" swimtime="00:00:51.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="329" reactiontime="+77" swimtime="00:01:22.07" resultid="108965" heatid="110693" lane="5" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.97" />
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="75" swimtime="00:01:03.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="292" reactiontime="+96" swimtime="00:00:36.74" resultid="108966" heatid="110738" lane="1" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="339" reactiontime="+82" swimtime="00:02:38.79" resultid="108967" heatid="110766" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.07" />
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="75" swimtime="00:00:56.59" />
                    <SPLIT distance="100" swimtime="00:01:17.16" />
                    <SPLIT distance="125" swimtime="00:01:37.73" />
                    <SPLIT distance="150" swimtime="00:01:58.81" />
                    <SPLIT distance="175" swimtime="00:02:19.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="252" reactiontime="+89" swimtime="00:01:26.45" resultid="108968" heatid="110795" lane="7" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.01" />
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="75" swimtime="00:01:01.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="447" reactiontime="+74" swimtime="00:01:58.36" resultid="109038" heatid="110719" lane="2" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.43" />
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="75" swimtime="00:00:48.19" />
                    <SPLIT distance="100" swimtime="00:01:05.57" />
                    <SPLIT distance="125" swimtime="00:01:18.10" />
                    <SPLIT distance="150" swimtime="00:01:32.74" />
                    <SPLIT distance="175" swimtime="00:01:45.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108988" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="109002" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="109030" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="108969" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="459" reactiontime="+75" swimtime="00:01:47.07" resultid="109040" heatid="110784" lane="7" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.51" />
                    <SPLIT distance="50" swimtime="00:00:25.39" />
                    <SPLIT distance="75" swimtime="00:00:38.66" />
                    <SPLIT distance="100" swimtime="00:00:53.23" />
                    <SPLIT distance="125" swimtime="00:01:06.50" />
                    <SPLIT distance="150" swimtime="00:01:21.27" />
                    <SPLIT distance="175" swimtime="00:01:33.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109030" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="108988" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="108978" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="108969" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT comment="S4/ IV ZMIANA" eventid="99059" reactiontime="+70" status="DSQ" swimtime="00:00:00.00" resultid="109039" heatid="110718" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.54" />
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="75" swimtime="00:00:48.87" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="125" swimtime="00:01:21.56" />
                    <SPLIT distance="150" swimtime="00:01:38.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109023" number="1" reactiontime="+70" status="DSQ" />
                    <RELAYPOSITION athleteid="108978" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="109008" number="3" reactiontime="+46" status="DSQ" />
                    <RELAYPOSITION athleteid="108994" number="4" reactiontime="-8" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="390" reactiontime="+77" swimtime="00:01:53.00" resultid="109041" heatid="110783" lane="4" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.65" />
                    <SPLIT distance="50" swimtime="00:00:28.27" />
                    <SPLIT distance="75" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:00:57.58" />
                    <SPLIT distance="125" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:25.50" />
                    <SPLIT distance="175" swimtime="00:01:38.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109023" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="108994" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="109008" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="109002" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="372" swimtime="00:01:54.83" resultid="109036" heatid="110632" lane="9" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.29" />
                    <SPLIT distance="50" swimtime="00:00:25.35" />
                    <SPLIT distance="75" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:00:56.91" />
                    <SPLIT distance="125" swimtime="00:01:11.94" />
                    <SPLIT distance="150" swimtime="00:01:28.65" />
                    <SPLIT distance="175" swimtime="00:01:41.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109030" number="1" />
                    <RELAYPOSITION athleteid="108962" number="2" />
                    <RELAYPOSITION athleteid="109015" number="3" />
                    <RELAYPOSITION athleteid="108969" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="99441" points="305" reactiontime="+67" swimtime="00:02:14.38" resultid="109037" heatid="110838" lane="0" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.81" />
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="75" swimtime="00:00:48.88" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="125" swimtime="00:01:22.86" />
                    <SPLIT distance="150" swimtime="00:01:42.47" />
                    <SPLIT distance="175" swimtime="00:01:57.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108988" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="109002" number="2" />
                    <RELAYPOSITION athleteid="109015" number="3" />
                    <RELAYPOSITION athleteid="108962" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="DOL" clubid="108358" name="UKS Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www.plywanie-zgorzelec.pl" name="Kondracki Łukasz" phone="693852488" state="DOL" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="108359">
              <RESULTS>
                <RESULT eventid="98798" points="105" reactiontime="+86" swimtime="00:00:42.92" resultid="108360" heatid="110597" lane="8" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="92" reactiontime="+96" swimtime="00:16:19.74" resultid="108361" heatid="110638" lane="8" entrytime="00:16:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.35" />
                    <SPLIT distance="50" swimtime="00:00:50.53" />
                    <SPLIT distance="75" swimtime="00:01:18.50" />
                    <SPLIT distance="100" swimtime="00:01:47.82" />
                    <SPLIT distance="125" swimtime="00:02:18.29" />
                    <SPLIT distance="150" swimtime="00:02:49.29" />
                    <SPLIT distance="175" swimtime="00:03:18.20" />
                    <SPLIT distance="200" swimtime="00:03:48.47" />
                    <SPLIT distance="225" swimtime="00:04:17.99" />
                    <SPLIT distance="250" swimtime="00:04:48.83" />
                    <SPLIT distance="275" swimtime="00:05:19.57" />
                    <SPLIT distance="300" swimtime="00:05:50.04" />
                    <SPLIT distance="325" swimtime="00:06:20.83" />
                    <SPLIT distance="350" swimtime="00:06:52.95" />
                    <SPLIT distance="375" swimtime="00:07:24.98" />
                    <SPLIT distance="400" swimtime="00:07:57.40" />
                    <SPLIT distance="425" swimtime="00:08:29.17" />
                    <SPLIT distance="450" swimtime="00:09:01.71" />
                    <SPLIT distance="475" swimtime="00:09:33.98" />
                    <SPLIT distance="500" swimtime="00:10:06.26" />
                    <SPLIT distance="525" swimtime="00:10:37.61" />
                    <SPLIT distance="550" swimtime="00:11:08.92" />
                    <SPLIT distance="575" swimtime="00:11:41.29" />
                    <SPLIT distance="600" swimtime="00:12:12.48" />
                    <SPLIT distance="625" swimtime="00:12:43.90" />
                    <SPLIT distance="650" swimtime="00:13:15.19" />
                    <SPLIT distance="675" swimtime="00:13:47.42" />
                    <SPLIT distance="700" swimtime="00:14:19.01" />
                    <SPLIT distance="725" swimtime="00:14:50.11" />
                    <SPLIT distance="750" swimtime="00:15:22.35" />
                    <SPLIT distance="775" swimtime="00:15:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="78" reactiontime="+87" swimtime="00:04:40.88" resultid="108362" heatid="110665" lane="5" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.96" />
                    <SPLIT distance="50" swimtime="00:01:03.51" />
                    <SPLIT distance="75" swimtime="00:01:38.66" />
                    <SPLIT distance="100" swimtime="00:02:15.09" />
                    <SPLIT distance="125" swimtime="00:02:51.53" />
                    <SPLIT distance="150" swimtime="00:03:27.91" />
                    <SPLIT distance="175" swimtime="00:04:03.61" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z2G3" eventid="98988" reactiontime="+93" status="DSQ" swimtime="00:00:00.00" resultid="108363" heatid="110696" lane="5" entrytime="00:01:58.00" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="108364" heatid="110758" lane="6" entrytime="00:01:50.00" />
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="108365" heatid="110788" lane="2" entrytime="00:09:15.00" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="108366" heatid="110811" lane="6" entrytime="00:03:50.00" />
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="108367" heatid="110851" lane="9" entrytime="00:08:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAL" clubid="107759" name="UKS SP 8 Chrzanów">
          <CONTACT city="Chrzanów" email="abalp@poczta.onet.pl" name="Zabrzański Alfred" phone="692076808" state="MAL" street="Niepodległości 7/46" zip="32-500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="107760">
              <RESULTS>
                <RESULT eventid="98798" points="273" reactiontime="+85" swimtime="00:00:31.20" resultid="107761" heatid="110602" lane="6" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="107762" heatid="110639" lane="4" entrytime="00:12:45.00" />
                <RESULT eventid="98924" points="168" reactiontime="+87" swimtime="00:00:40.22" resultid="107763" heatid="110654" lane="1" entrytime="00:00:41.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="256" reactiontime="+90" swimtime="00:01:10.76" resultid="107764" heatid="110682" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.80" />
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="75" swimtime="00:00:51.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="192" reactiontime="+102" swimtime="00:01:36.31" resultid="107765" heatid="110729" lane="1" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.42" />
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                    <SPLIT distance="75" swimtime="00:01:10.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="225" reactiontime="+89" swimtime="00:02:43.33" resultid="107766" heatid="110772" lane="7" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="75" swimtime="00:00:55.74" />
                    <SPLIT distance="100" swimtime="00:01:16.26" />
                    <SPLIT distance="125" swimtime="00:01:37.62" />
                    <SPLIT distance="150" swimtime="00:01:59.07" />
                    <SPLIT distance="175" swimtime="00:02:21.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="184" reactiontime="+90" swimtime="00:00:44.35" resultid="107767" heatid="110826" lane="5" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="107768" heatid="110849" lane="0" entrytime="00:06:16.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" region="KA" clubid="106995" name="UKS Wodnik 29 Katowice">
          <CONTACT email="skoczyt@gmail.com" name="Skoczylas Tomasz" />
          <ATHLETES>
            <ATHLETE birthdate="1983-05-05" firstname="Marek" gender="M" lastname="Mróz" nation="POL" athleteid="107020">
              <RESULTS>
                <RESULT eventid="98798" status="WDR" swimtime="00:00:00.00" resultid="107021" entrytime="00:00:26.00" />
                <RESULT eventid="106277" status="WDR" swimtime="00:00:00.00" resultid="107022" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-09" firstname="Krystyna" gender="F" lastname="Nicpoń" nation="POL" athleteid="107011">
              <RESULTS>
                <RESULT eventid="98814" points="85" reactiontime="+119" swimtime="00:04:36.94" resultid="107012" heatid="110614" lane="2" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.17" />
                    <SPLIT distance="50" swimtime="00:01:14.52" />
                    <SPLIT distance="75" swimtime="00:01:45.62" />
                    <SPLIT distance="100" swimtime="00:02:16.22" />
                    <SPLIT distance="125" swimtime="00:02:54.02" />
                    <SPLIT distance="150" swimtime="00:03:32.78" />
                    <SPLIT distance="175" swimtime="00:04:04.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106254" points="93" reactiontime="+102" swimtime="00:33:44.99" resultid="107013" heatid="110640" lane="0" entrytime="00:36:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.73" />
                    <SPLIT distance="50" swimtime="00:00:53.40" />
                    <SPLIT distance="75" swimtime="00:01:25.31" />
                    <SPLIT distance="100" swimtime="00:01:58.33" />
                    <SPLIT distance="125" swimtime="00:02:31.56" />
                    <SPLIT distance="150" swimtime="00:03:05.23" />
                    <SPLIT distance="175" swimtime="00:03:38.42" />
                    <SPLIT distance="200" swimtime="00:04:12.20" />
                    <SPLIT distance="225" swimtime="00:04:46.78" />
                    <SPLIT distance="250" swimtime="00:05:20.83" />
                    <SPLIT distance="275" swimtime="00:05:54.50" />
                    <SPLIT distance="300" swimtime="00:06:27.98" />
                    <SPLIT distance="325" swimtime="00:07:01.94" />
                    <SPLIT distance="350" swimtime="00:07:35.59" />
                    <SPLIT distance="375" swimtime="00:08:09.57" />
                    <SPLIT distance="400" swimtime="00:08:42.91" />
                    <SPLIT distance="425" swimtime="00:09:16.84" />
                    <SPLIT distance="450" swimtime="00:09:50.99" />
                    <SPLIT distance="475" swimtime="00:10:24.86" />
                    <SPLIT distance="500" swimtime="00:10:58.50" />
                    <SPLIT distance="525" swimtime="00:11:31.81" />
                    <SPLIT distance="550" swimtime="00:12:05.48" />
                    <SPLIT distance="575" swimtime="00:12:39.18" />
                    <SPLIT distance="600" swimtime="00:13:13.21" />
                    <SPLIT distance="625" swimtime="00:13:47.17" />
                    <SPLIT distance="650" swimtime="00:14:21.21" />
                    <SPLIT distance="675" swimtime="00:14:55.33" />
                    <SPLIT distance="700" swimtime="00:15:29.41" />
                    <SPLIT distance="725" swimtime="00:16:03.17" />
                    <SPLIT distance="750" swimtime="00:16:37.09" />
                    <SPLIT distance="775" swimtime="00:17:09.80" />
                    <SPLIT distance="800" swimtime="00:17:43.77" />
                    <SPLIT distance="825" swimtime="00:18:17.86" />
                    <SPLIT distance="850" swimtime="00:18:52.39" />
                    <SPLIT distance="875" swimtime="00:19:26.10" />
                    <SPLIT distance="900" swimtime="00:20:00.29" />
                    <SPLIT distance="925" swimtime="00:20:34.28" />
                    <SPLIT distance="950" swimtime="00:21:08.82" />
                    <SPLIT distance="975" swimtime="00:21:42.78" />
                    <SPLIT distance="1000" swimtime="00:22:17.49" />
                    <SPLIT distance="1025" swimtime="00:22:51.55" />
                    <SPLIT distance="1050" swimtime="00:23:26.04" />
                    <SPLIT distance="1075" swimtime="00:23:59.87" />
                    <SPLIT distance="1100" swimtime="00:24:34.69" />
                    <SPLIT distance="1125" swimtime="00:25:08.83" />
                    <SPLIT distance="1150" swimtime="00:25:42.90" />
                    <SPLIT distance="1175" swimtime="00:26:17.60" />
                    <SPLIT distance="1200" swimtime="00:26:52.79" />
                    <SPLIT distance="1225" swimtime="00:27:26.66" />
                    <SPLIT distance="1250" swimtime="00:28:01.71" />
                    <SPLIT distance="1275" swimtime="00:28:35.48" />
                    <SPLIT distance="1300" swimtime="00:29:10.74" />
                    <SPLIT distance="1325" swimtime="00:29:44.75" />
                    <SPLIT distance="1350" swimtime="00:30:19.61" />
                    <SPLIT distance="1375" swimtime="00:30:54.85" />
                    <SPLIT distance="1400" swimtime="00:31:29.44" />
                    <SPLIT distance="1425" swimtime="00:32:03.84" />
                    <SPLIT distance="1450" swimtime="00:32:38.00" />
                    <SPLIT distance="1475" swimtime="00:33:11.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="106" reactiontime="+100" swimtime="00:00:54.10" resultid="107014" heatid="110646" lane="4" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="83" swimtime="00:02:09.52" resultid="107015" heatid="110690" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.02" />
                    <SPLIT distance="50" swimtime="00:01:03.23" />
                    <SPLIT distance="75" swimtime="00:01:39.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="35" reactiontime="+100" swimtime="00:01:14.47" resultid="107016" heatid="110735" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="95" reactiontime="+92" swimtime="00:02:00.28" resultid="107017" heatid="110753" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.20" />
                    <SPLIT distance="50" swimtime="00:00:57.54" />
                    <SPLIT distance="75" swimtime="00:01:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="112" reactiontime="+91" swimtime="00:04:07.28" resultid="107018" heatid="110806" lane="4" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.81" />
                    <SPLIT distance="50" swimtime="00:00:56.76" />
                    <SPLIT distance="75" swimtime="00:01:27.20" />
                    <SPLIT distance="100" swimtime="00:01:59.08" />
                    <SPLIT distance="125" swimtime="00:02:31.23" />
                    <SPLIT distance="150" swimtime="00:03:04.24" />
                    <SPLIT distance="175" swimtime="00:03:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="94" reactiontime="+116" swimtime="00:08:34.69" resultid="107019" heatid="110842" lane="8" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.17" />
                    <SPLIT distance="50" swimtime="00:00:54.25" />
                    <SPLIT distance="75" swimtime="00:01:26.08" />
                    <SPLIT distance="100" swimtime="00:01:58.41" />
                    <SPLIT distance="125" swimtime="00:02:30.79" />
                    <SPLIT distance="150" swimtime="00:03:04.51" />
                    <SPLIT distance="175" swimtime="00:03:35.87" />
                    <SPLIT distance="200" swimtime="00:04:09.47" />
                    <SPLIT distance="225" swimtime="00:04:42.49" />
                    <SPLIT distance="250" swimtime="00:05:15.88" />
                    <SPLIT distance="275" swimtime="00:05:49.79" />
                    <SPLIT distance="300" swimtime="00:06:22.99" />
                    <SPLIT distance="325" swimtime="00:06:56.52" />
                    <SPLIT distance="350" swimtime="00:07:31.05" />
                    <SPLIT distance="375" swimtime="00:08:03.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="106996">
              <RESULTS>
                <RESULT eventid="98798" points="364" reactiontime="+88" swimtime="00:00:28.35" resultid="106997" heatid="110607" lane="7" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="356" reactiontime="+100" swimtime="00:19:56.16" resultid="106998" heatid="110641" lane="8" entrytime="00:20:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.18" />
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="75" swimtime="00:00:52.57" />
                    <SPLIT distance="100" swimtime="00:01:11.85" />
                    <SPLIT distance="125" swimtime="00:01:30.97" />
                    <SPLIT distance="150" swimtime="00:01:50.42" />
                    <SPLIT distance="175" swimtime="00:02:09.89" />
                    <SPLIT distance="200" swimtime="00:02:29.47" />
                    <SPLIT distance="225" swimtime="00:02:49.00" />
                    <SPLIT distance="250" swimtime="00:03:08.74" />
                    <SPLIT distance="275" swimtime="00:03:28.41" />
                    <SPLIT distance="300" swimtime="00:03:47.96" />
                    <SPLIT distance="325" swimtime="00:04:07.59" />
                    <SPLIT distance="350" swimtime="00:04:27.36" />
                    <SPLIT distance="375" swimtime="00:04:47.26" />
                    <SPLIT distance="400" swimtime="00:05:07.02" />
                    <SPLIT distance="425" swimtime="00:05:26.95" />
                    <SPLIT distance="450" swimtime="00:05:47.29" />
                    <SPLIT distance="475" swimtime="00:06:07.28" />
                    <SPLIT distance="500" swimtime="00:06:27.37" />
                    <SPLIT distance="525" swimtime="00:06:47.38" />
                    <SPLIT distance="550" swimtime="00:07:07.65" />
                    <SPLIT distance="575" swimtime="00:07:27.74" />
                    <SPLIT distance="600" swimtime="00:07:47.91" />
                    <SPLIT distance="625" swimtime="00:08:07.99" />
                    <SPLIT distance="650" swimtime="00:08:28.09" />
                    <SPLIT distance="675" swimtime="00:08:48.66" />
                    <SPLIT distance="700" swimtime="00:09:09.02" />
                    <SPLIT distance="725" swimtime="00:09:29.19" />
                    <SPLIT distance="750" swimtime="00:09:49.44" />
                    <SPLIT distance="775" swimtime="00:10:09.68" />
                    <SPLIT distance="800" swimtime="00:10:29.62" />
                    <SPLIT distance="825" swimtime="00:10:49.75" />
                    <SPLIT distance="850" swimtime="00:11:09.88" />
                    <SPLIT distance="875" swimtime="00:11:30.20" />
                    <SPLIT distance="900" swimtime="00:11:50.52" />
                    <SPLIT distance="925" swimtime="00:12:10.93" />
                    <SPLIT distance="950" swimtime="00:12:31.12" />
                    <SPLIT distance="975" swimtime="00:12:51.43" />
                    <SPLIT distance="1000" swimtime="00:13:11.89" />
                    <SPLIT distance="1025" swimtime="00:13:32.24" />
                    <SPLIT distance="1050" swimtime="00:13:52.44" />
                    <SPLIT distance="1075" swimtime="00:14:12.77" />
                    <SPLIT distance="1100" swimtime="00:14:32.83" />
                    <SPLIT distance="1125" swimtime="00:14:53.17" />
                    <SPLIT distance="1150" swimtime="00:15:13.50" />
                    <SPLIT distance="1175" swimtime="00:15:33.79" />
                    <SPLIT distance="1200" swimtime="00:15:54.11" />
                    <SPLIT distance="1225" swimtime="00:16:14.48" />
                    <SPLIT distance="1250" swimtime="00:16:34.84" />
                    <SPLIT distance="1275" swimtime="00:16:55.31" />
                    <SPLIT distance="1300" swimtime="00:17:15.74" />
                    <SPLIT distance="1325" swimtime="00:17:35.79" />
                    <SPLIT distance="1350" swimtime="00:17:56.14" />
                    <SPLIT distance="1375" swimtime="00:18:16.19" />
                    <SPLIT distance="1400" swimtime="00:18:36.20" />
                    <SPLIT distance="1425" swimtime="00:18:56.25" />
                    <SPLIT distance="1450" swimtime="00:19:16.56" />
                    <SPLIT distance="1475" swimtime="00:19:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="357" reactiontime="+90" swimtime="00:01:03.30" resultid="106999" heatid="110685" lane="8" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.72" />
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="75" swimtime="00:00:46.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="225" reactiontime="+110" swimtime="00:02:58.34" resultid="107000" heatid="110712" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.05" />
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="75" swimtime="00:00:59.99" />
                    <SPLIT distance="100" swimtime="00:01:22.65" />
                    <SPLIT distance="125" swimtime="00:01:45.85" />
                    <SPLIT distance="150" swimtime="00:02:09.58" />
                    <SPLIT distance="175" swimtime="00:02:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="273" reactiontime="+97" swimtime="00:01:15.35" resultid="107001" heatid="110760" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.01" />
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="75" swimtime="00:00:56.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="350" reactiontime="+77" swimtime="00:02:20.92" resultid="107002" heatid="110774" lane="7" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="75" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                    <SPLIT distance="125" swimtime="00:01:27.07" />
                    <SPLIT distance="150" swimtime="00:01:45.42" />
                    <SPLIT distance="175" swimtime="00:02:03.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="219" reactiontime="+78" swimtime="00:01:20.29" resultid="107003" heatid="110801" lane="7" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.38" />
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="75" swimtime="00:00:58.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="350" reactiontime="+85" swimtime="00:05:01.05" resultid="107004" heatid="110846" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.20" />
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="75" swimtime="00:00:52.15" />
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                    <SPLIT distance="125" swimtime="00:01:29.63" />
                    <SPLIT distance="150" swimtime="00:01:49.21" />
                    <SPLIT distance="175" swimtime="00:02:08.89" />
                    <SPLIT distance="200" swimtime="00:02:28.65" />
                    <SPLIT distance="225" swimtime="00:02:48.03" />
                    <SPLIT distance="250" swimtime="00:03:07.68" />
                    <SPLIT distance="275" swimtime="00:03:26.98" />
                    <SPLIT distance="300" swimtime="00:03:46.69" />
                    <SPLIT distance="325" swimtime="00:04:05.70" />
                    <SPLIT distance="350" swimtime="00:04:24.69" />
                    <SPLIT distance="375" swimtime="00:04:43.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="107005">
              <RESULTS>
                <RESULT eventid="98798" points="276" reactiontime="+90" swimtime="00:00:31.09" resultid="107006" heatid="110601" lane="2" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="305" swimtime="00:02:58.92" resultid="107007" heatid="110669" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.04" />
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="75" swimtime="00:01:02.51" />
                    <SPLIT distance="100" swimtime="00:01:25.88" />
                    <SPLIT distance="125" swimtime="00:01:49.08" />
                    <SPLIT distance="150" swimtime="00:02:12.82" />
                    <SPLIT distance="175" swimtime="00:02:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="313" reactiontime="+79" swimtime="00:01:14.55" resultid="107008" heatid="110700" lane="7" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="75" swimtime="00:00:55.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="346" reactiontime="+69" swimtime="00:01:19.18" resultid="107009" heatid="110732" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.70" />
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="75" swimtime="00:00:57.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="365" reactiontime="+83" swimtime="00:00:35.30" resultid="107010" heatid="110830" lane="4" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" nation="POL" region="WAR" clubid="107125" name="Ursynów Masters">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1968-06-01" firstname="Robert" gender="M" lastname="Zieliński" nation="POL" athleteid="107148">
              <RESULTS>
                <RESULT eventid="98798" points="232" reactiontime="+74" swimtime="00:00:32.96" resultid="107149" heatid="110601" lane="7" entrytime="00:00:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="160" reactiontime="+89" swimtime="00:03:21.62" resultid="107150" heatid="110621" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.25" />
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="75" swimtime="00:02:06.39" />
                    <SPLIT distance="100" swimtime="00:01:36.28" />
                    <SPLIT distance="125" swimtime="00:03:00.38" />
                    <SPLIT distance="150" swimtime="00:02:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="168" reactiontime="+76" swimtime="00:00:40.26" resultid="107151" heatid="110654" lane="9" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="175" reactiontime="+74" swimtime="00:01:30.48" resultid="107152" heatid="110697" lane="6" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="75" swimtime="00:01:09.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="172" reactiontime="+82" swimtime="00:01:39.94" resultid="107153" heatid="110728" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.82" />
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                    <SPLIT distance="75" swimtime="00:01:14.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="193" reactiontime="+78" swimtime="00:02:51.67" resultid="107154" heatid="110771" lane="7" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.80" />
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="75" swimtime="00:00:58.37" />
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="125" swimtime="00:01:41.77" />
                    <SPLIT distance="150" swimtime="00:02:04.61" />
                    <SPLIT distance="175" swimtime="00:02:29.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="107155" heatid="110812" lane="1" entrytime="00:03:30.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="107156" heatid="110826" lane="9" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="Rybarczyk" nation="POL" athleteid="107134">
              <RESULTS>
                <RESULT eventid="98798" points="346" swimtime="00:00:28.84" resultid="107135" heatid="110605" lane="9" entrytime="00:00:29.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="128" reactiontime="+69" swimtime="00:00:43.99" resultid="107136" heatid="110654" lane="6" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="318" reactiontime="+74" swimtime="00:01:05.78" resultid="107137" heatid="110683" lane="5" entrytime="00:01:05.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.95" />
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="75" swimtime="00:00:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="275" reactiontime="+91" swimtime="00:00:33.49" resultid="107138" heatid="110745" lane="1" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="276" reactiontime="+66" swimtime="00:02:32.50" resultid="107139" heatid="110773" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.51" />
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="75" swimtime="00:00:52.13" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="125" swimtime="00:01:31.71" />
                    <SPLIT distance="150" swimtime="00:01:52.40" />
                    <SPLIT distance="175" swimtime="00:02:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="107140" heatid="110800" lane="3" entrytime="00:01:23.00" />
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="107141" heatid="110848" lane="3" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="Nowak" nation="POL" athleteid="107126">
              <RESULTS>
                <RESULT eventid="98830" points="218" reactiontime="+87" swimtime="00:03:01.95" resultid="107127" heatid="110622" lane="3" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.88" />
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="75" swimtime="00:01:04.96" />
                    <SPLIT distance="100" swimtime="00:01:28.59" />
                    <SPLIT distance="125" swimtime="00:01:53.24" />
                    <SPLIT distance="150" swimtime="00:02:18.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="256" reactiontime="+66" swimtime="00:03:09.73" resultid="107128" heatid="110668" lane="2" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.14" />
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                    <SPLIT distance="75" swimtime="00:01:05.21" />
                    <SPLIT distance="100" swimtime="00:01:29.17" />
                    <SPLIT distance="125" swimtime="00:01:53.54" />
                    <SPLIT distance="150" swimtime="00:02:18.60" />
                    <SPLIT distance="175" swimtime="00:02:44.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="281" reactiontime="+81" swimtime="00:01:17.27" resultid="107129" heatid="110699" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.53" />
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="75" swimtime="00:00:58.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="295" reactiontime="+70" swimtime="00:01:23.45" resultid="107130" heatid="110731" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.58" />
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="75" swimtime="00:01:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="185" reactiontime="+73" swimtime="00:06:53.18" resultid="107131" heatid="110789" lane="2" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.31" />
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="75" swimtime="00:01:13.73" />
                    <SPLIT distance="100" swimtime="00:01:42.44" />
                    <SPLIT distance="125" swimtime="00:03:03.52" />
                    <SPLIT distance="150" swimtime="00:03:30.68" />
                    <SPLIT distance="175" swimtime="00:03:57.06" />
                    <SPLIT distance="200" swimtime="00:04:23.48" />
                    <SPLIT distance="225" swimtime="00:04:49.96" />
                    <SPLIT distance="250" swimtime="00:05:17.40" />
                    <SPLIT distance="275" swimtime="00:06:31.13" />
                    <SPLIT distance="300" swimtime="00:06:53.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="133" swimtime="00:01:34.71" resultid="107132" heatid="110800" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.67" />
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                    <SPLIT distance="75" swimtime="00:01:07.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="324" reactiontime="+84" swimtime="00:00:36.76" resultid="107133" heatid="110830" lane="1" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-03-23" firstname="Ryszard" gender="M" lastname="Rybarczyk" nation="POL" athleteid="107142">
              <RESULTS>
                <RESULT eventid="98798" points="84" reactiontime="+103" swimtime="00:00:46.23" resultid="107143" heatid="110596" lane="3" entrytime="00:00:41.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="55" reactiontime="+102" swimtime="00:00:58.42" resultid="107144" heatid="110652" lane="7" entrytime="00:00:56.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="113" reactiontime="+109" swimtime="00:01:54.97" resultid="107145" heatid="110727" lane="3" entrytime="00:01:58.93">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.65" />
                    <SPLIT distance="50" swimtime="00:00:54.43" />
                    <SPLIT distance="75" swimtime="00:01:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="107146" heatid="110757" lane="4" entrytime="00:02:12.00" />
                <RESULT eventid="99425" points="125" reactiontime="+100" swimtime="00:00:50.46" resultid="107147" heatid="110825" lane="5" entrytime="00:00:48.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="199" reactiontime="+67" swimtime="00:02:34.77" resultid="107157" heatid="110717" lane="0" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.26" />
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="75" swimtime="00:00:57.61" />
                    <SPLIT distance="100" swimtime="00:01:16.74" />
                    <SPLIT distance="125" swimtime="00:01:31.93" />
                    <SPLIT distance="150" swimtime="00:01:50.49" />
                    <SPLIT distance="175" swimtime="00:02:11.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107148" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="107126" number="2" />
                    <RELAYPOSITION athleteid="107134" number="3" />
                    <RELAYPOSITION athleteid="107142" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="214" reactiontime="+74" swimtime="00:02:17.94" resultid="107158" heatid="110782" lane="8" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.86" />
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="75" swimtime="00:00:52.90" />
                    <SPLIT distance="100" swimtime="00:01:15.59" />
                    <SPLIT distance="125" swimtime="00:01:31.56" />
                    <SPLIT distance="150" swimtime="00:01:48.89" />
                    <SPLIT distance="175" swimtime="00:02:02.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107126" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="107142" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="107148" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="107134" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="031" nation="POL" region="LOD" clubid="108002" name="UTW Masters Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="108012">
              <RESULTS>
                <RESULT eventid="98777" points="354" reactiontime="+86" swimtime="00:00:32.84" resultid="108013" heatid="110590" lane="8" entrytime="00:00:33.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="302" reactiontime="+82" swimtime="00:00:38.23" resultid="108014" heatid="110649" lane="6" entrytime="00:00:37.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="210" reactiontime="+94" swimtime="00:03:21.20" resultid="108015" heatid="110708" lane="7" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.23" />
                    <SPLIT distance="50" swimtime="00:00:21.53" />
                    <SPLIT distance="75" swimtime="00:01:08.73" />
                    <SPLIT distance="100" swimtime="00:00:43.84" />
                    <SPLIT distance="125" swimtime="00:02:00.86" />
                    <SPLIT distance="150" swimtime="00:02:27.52" />
                    <SPLIT distance="175" swimtime="00:02:55.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="354" reactiontime="+91" swimtime="00:00:34.45" resultid="108016" heatid="110739" lane="8" entrytime="00:00:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="237" reactiontime="+95" swimtime="00:01:28.85" resultid="108017" heatid="110755" lane="3" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.64" />
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="75" swimtime="00:01:06.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="245" swimtime="00:01:27.16" resultid="108018" heatid="110795" lane="9" entrytime="00:01:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.29" />
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="75" swimtime="00:01:02.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" status="DNS" swimtime="00:00:00.00" resultid="108019" heatid="110808" lane="3" entrytime="00:03:10.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-25" firstname="Michał" gender="M" lastname="Wożniak" nation="POL" license="503105700039" athleteid="108056">
              <RESULTS>
                <RESULT eventid="98924" points="357" reactiontime="+75" swimtime="00:00:31.32" resultid="108057" heatid="110659" lane="7" entrytime="00:00:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="108058" heatid="110703" lane="0" entrytime="00:01:10.50" entrycourse="SCM" />
                <RESULT eventid="99186" points="387" reactiontime="+64" swimtime="00:01:07.10" resultid="108059" heatid="110762" lane="5" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.55" />
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="75" swimtime="00:00:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="374" reactiontime="+70" swimtime="00:02:26.55" resultid="108060" heatid="110815" lane="7" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.71" />
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="75" swimtime="00:00:50.95" />
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                    <SPLIT distance="125" swimtime="00:01:28.91" />
                    <SPLIT distance="150" swimtime="00:01:48.36" />
                    <SPLIT distance="175" swimtime="00:02:07.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105600018" athleteid="108082">
              <RESULTS>
                <RESULT eventid="98777" points="486" reactiontime="+86" swimtime="00:00:29.55" resultid="108083" heatid="110592" lane="5" entrytime="00:00:28.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="419" reactiontime="+99" swimtime="00:02:42.82" resultid="108084" heatid="110616" lane="0" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.28" />
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="75" swimtime="00:00:53.72" />
                    <SPLIT distance="100" swimtime="00:01:13.62" />
                    <SPLIT distance="125" swimtime="00:01:37.26" />
                    <SPLIT distance="150" swimtime="00:02:01.47" />
                    <SPLIT distance="175" swimtime="00:02:22.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="460" reactiontime="+85" swimtime="00:00:33.25" resultid="108085" heatid="110650" lane="3" entrytime="00:00:31.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="438" reactiontime="+88" swimtime="00:01:14.57" resultid="108086" heatid="110694" lane="2" entrytime="00:01:19.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="75" swimtime="00:00:56.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="395" reactiontime="+86" swimtime="00:00:33.22" resultid="108087" heatid="110740" lane="7" entrytime="00:00:30.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="416" reactiontime="+82" swimtime="00:01:13.67" resultid="108088" heatid="110756" lane="3" entrytime="00:01:11.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="75" swimtime="00:00:53.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="369" reactiontime="+70" swimtime="00:02:46.13" resultid="108089" heatid="110807" lane="6" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.67" />
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="75" swimtime="00:00:56.97" />
                    <SPLIT distance="100" swimtime="00:01:18.19" />
                    <SPLIT distance="125" swimtime="00:01:40.36" />
                    <SPLIT distance="150" swimtime="00:02:02.61" />
                    <SPLIT distance="175" swimtime="00:02:24.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700034" athleteid="108007">
              <RESULTS>
                <RESULT eventid="98798" points="152" reactiontime="+99" swimtime="00:00:37.90" resultid="108008" heatid="110598" lane="3" entrytime="00:00:37.50" entrycourse="SCM" />
                <RESULT eventid="98956" points="189" reactiontime="+90" swimtime="00:03:29.88" resultid="108009" heatid="110666" lane="5" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.35" />
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                    <SPLIT distance="75" swimtime="00:01:13.08" />
                    <SPLIT distance="100" swimtime="00:01:40.55" />
                    <SPLIT distance="125" swimtime="00:02:07.95" />
                    <SPLIT distance="150" swimtime="00:02:35.83" />
                    <SPLIT distance="175" swimtime="00:03:03.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="204" swimtime="00:01:34.34" resultid="108010" heatid="110730" lane="9" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.59" />
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                    <SPLIT distance="75" swimtime="00:01:09.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="242" reactiontime="+86" swimtime="00:00:40.51" resultid="108011" heatid="110827" lane="5" entrytime="00:00:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700027" athleteid="108020">
              <RESULTS>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="108021" heatid="110623" lane="1" entrytime="00:02:57.00" entrycourse="SCM" />
                <RESULT eventid="106256" points="244" swimtime="00:22:36.47" resultid="108022" heatid="110642" lane="9" entrytime="00:23:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="75" swimtime="00:00:57.87" />
                    <SPLIT distance="100" swimtime="00:01:19.37" />
                    <SPLIT distance="125" swimtime="00:01:41.48" />
                    <SPLIT distance="150" swimtime="00:02:04.18" />
                    <SPLIT distance="175" swimtime="00:02:26.37" />
                    <SPLIT distance="200" swimtime="00:02:49.12" />
                    <SPLIT distance="225" swimtime="00:03:11.30" />
                    <SPLIT distance="250" swimtime="00:03:33.86" />
                    <SPLIT distance="275" swimtime="00:03:56.32" />
                    <SPLIT distance="300" swimtime="00:04:18.69" />
                    <SPLIT distance="325" swimtime="00:04:41.30" />
                    <SPLIT distance="350" swimtime="00:05:03.97" />
                    <SPLIT distance="375" swimtime="00:05:26.61" />
                    <SPLIT distance="400" swimtime="00:05:49.75" />
                    <SPLIT distance="425" swimtime="00:06:12.69" />
                    <SPLIT distance="450" swimtime="00:06:35.66" />
                    <SPLIT distance="475" swimtime="00:06:58.24" />
                    <SPLIT distance="500" swimtime="00:07:21.36" />
                    <SPLIT distance="525" swimtime="00:07:44.39" />
                    <SPLIT distance="550" swimtime="00:08:07.40" />
                    <SPLIT distance="575" swimtime="00:08:29.98" />
                    <SPLIT distance="600" swimtime="00:08:53.27" />
                    <SPLIT distance="625" swimtime="00:09:16.17" />
                    <SPLIT distance="650" swimtime="00:09:39.67" />
                    <SPLIT distance="675" swimtime="00:10:02.19" />
                    <SPLIT distance="700" swimtime="00:10:25.34" />
                    <SPLIT distance="725" swimtime="00:10:48.08" />
                    <SPLIT distance="750" swimtime="00:11:11.38" />
                    <SPLIT distance="775" swimtime="00:11:34.21" />
                    <SPLIT distance="800" swimtime="00:11:57.77" />
                    <SPLIT distance="825" swimtime="00:12:20.69" />
                    <SPLIT distance="850" swimtime="00:12:44.07" />
                    <SPLIT distance="875" swimtime="00:13:06.99" />
                    <SPLIT distance="900" swimtime="00:13:30.59" />
                    <SPLIT distance="925" swimtime="00:13:53.93" />
                    <SPLIT distance="950" swimtime="00:14:17.24" />
                    <SPLIT distance="975" swimtime="00:14:39.86" />
                    <SPLIT distance="1000" swimtime="00:15:03.27" />
                    <SPLIT distance="1025" swimtime="00:15:25.85" />
                    <SPLIT distance="1050" swimtime="00:15:49.05" />
                    <SPLIT distance="1075" swimtime="00:16:11.80" />
                    <SPLIT distance="1100" swimtime="00:16:35.24" />
                    <SPLIT distance="1125" swimtime="00:16:58.31" />
                    <SPLIT distance="1150" swimtime="00:17:21.40" />
                    <SPLIT distance="1175" swimtime="00:17:44.06" />
                    <SPLIT distance="1200" swimtime="00:18:07.83" />
                    <SPLIT distance="1225" swimtime="00:18:30.35" />
                    <SPLIT distance="1250" swimtime="00:18:53.57" />
                    <SPLIT distance="1275" swimtime="00:19:15.85" />
                    <SPLIT distance="1300" swimtime="00:19:38.94" />
                    <SPLIT distance="1325" swimtime="00:20:01.66" />
                    <SPLIT distance="1350" swimtime="00:20:24.68" />
                    <SPLIT distance="1375" swimtime="00:20:47.40" />
                    <SPLIT distance="1400" swimtime="00:21:10.13" />
                    <SPLIT distance="1425" swimtime="00:21:32.37" />
                    <SPLIT distance="1450" swimtime="00:21:54.87" />
                    <SPLIT distance="1475" swimtime="00:22:16.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="236" reactiontime="+83" swimtime="00:00:35.95" resultid="108023" heatid="110655" lane="3" entrytime="00:00:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="303" swimtime="00:01:06.87" resultid="108024" heatid="110683" lane="0" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="75" swimtime="00:00:49.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="293" reactiontime="+86" swimtime="00:00:32.81" resultid="108025" heatid="110745" lane="3" entrytime="00:00:32.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="299" reactiontime="+85" swimtime="00:02:28.45" resultid="108026" heatid="110773" lane="4" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.13" />
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="75" swimtime="00:00:52.14" />
                    <SPLIT distance="100" swimtime="00:01:10.61" />
                    <SPLIT distance="125" swimtime="00:01:30.11" />
                    <SPLIT distance="150" swimtime="00:01:49.56" />
                    <SPLIT distance="175" swimtime="00:02:09.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="228" reactiontime="+89" swimtime="00:01:19.20" resultid="108027" heatid="110800" lane="4" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.39" />
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="75" swimtime="00:00:56.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="108028" heatid="110813" lane="1" entrytime="00:03:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="108029">
              <RESULTS>
                <RESULT eventid="98798" points="226" reactiontime="+93" swimtime="00:00:33.22" resultid="108030" heatid="110600" lane="4" entrytime="00:00:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="123" reactiontime="+109" swimtime="00:03:40.11" resultid="108031" heatid="110620" lane="3" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.44" />
                    <SPLIT distance="50" swimtime="00:00:54.43" />
                    <SPLIT distance="75" swimtime="00:01:22.02" />
                    <SPLIT distance="100" swimtime="00:01:51.38" />
                    <SPLIT distance="125" swimtime="00:02:23.85" />
                    <SPLIT distance="150" swimtime="00:02:58.05" />
                    <SPLIT distance="175" swimtime="00:03:20.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="149" reactiontime="+103" swimtime="00:01:35.50" resultid="108032" heatid="110697" lane="3" entrytime="00:01:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.61" />
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                    <SPLIT distance="75" swimtime="00:01:15.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="108033" heatid="110710" lane="6" entrytime="00:04:08.00" entrycourse="SCM" />
                <RESULT eventid="99170" points="210" swimtime="00:00:36.62" resultid="108034" heatid="110743" lane="6" entrytime="00:00:36.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="108035" heatid="110758" lane="1" entrytime="00:01:52.00" entrycourse="SCM" />
                <RESULT eventid="99361" points="102" swimtime="00:01:43.45" resultid="108036" heatid="110799" lane="2" entrytime="00:01:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.62" />
                    <SPLIT distance="50" swimtime="00:00:52.17" />
                    <SPLIT distance="75" swimtime="00:01:22.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="108037" heatid="110850" lane="3" entrytime="00:06:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1922-01-04" firstname="Kazimierz" gender="M" lastname="Mrówczyński" nation="POL" license="503105700021" athleteid="108003">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="108004" heatid="110595" lane="2" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="108005" heatid="110678" lane="2" entrytime="00:02:10.00" entrycourse="SCM" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="108006" heatid="110824" lane="3" entrytime="00:01:11.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-16" firstname="Krzysztof" gender="M" lastname="Gawłowicz" nation="POL" athleteid="106439">
              <RESULTS>
                <RESULT eventid="98798" points="534" reactiontime="+70" swimtime="00:00:24.97" resultid="106440" heatid="110612" lane="4" entrytime="00:00:24.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="544" reactiontime="+68" swimtime="00:00:26.70" resultid="106441" heatid="110751" lane="7" entrytime="00:00:25.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-08" firstname="Ewa" gender="F" lastname="Zimna-Walendzik" nation="POL" license="03105600019" athleteid="108090">
              <RESULTS>
                <RESULT eventid="98777" points="167" reactiontime="+101" swimtime="00:00:42.16" resultid="108091" heatid="110587" lane="2" entrytime="00:00:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="141" swimtime="00:03:54.09" resultid="108092" heatid="110614" lane="4" entrytime="00:03:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.20" />
                    <SPLIT distance="50" swimtime="00:00:53.44" />
                    <SPLIT distance="75" swimtime="00:01:23.77" />
                    <SPLIT distance="100" swimtime="00:01:55.32" />
                    <SPLIT distance="125" swimtime="00:02:27.76" />
                    <SPLIT distance="150" swimtime="00:02:59.54" />
                    <SPLIT distance="175" swimtime="00:03:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="139" swimtime="00:01:49.25" resultid="108093" heatid="110691" lane="0" entrytime="00:01:49.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.93" />
                    <SPLIT distance="50" swimtime="00:00:52.36" />
                    <SPLIT distance="75" swimtime="00:01:23.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="90" swimtime="00:04:26.06" resultid="108094" heatid="110707" lane="4" entrytime="00:04:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.96" />
                    <SPLIT distance="50" swimtime="00:00:56.16" />
                    <SPLIT distance="75" swimtime="00:01:29.13" />
                    <SPLIT distance="100" swimtime="00:02:02.73" />
                    <SPLIT distance="125" swimtime="00:02:38.75" />
                    <SPLIT distance="150" swimtime="00:03:15.96" />
                    <SPLIT distance="175" swimtime="00:03:53.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="112" reactiontime="+83" swimtime="00:00:50.45" resultid="108095" heatid="110736" lane="7" entrytime="00:00:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="130" swimtime="00:03:38.39" resultid="108096" heatid="110764" lane="3" entrytime="00:03:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.04" />
                    <SPLIT distance="50" swimtime="00:00:49.21" />
                    <SPLIT distance="75" swimtime="00:01:16.62" />
                    <SPLIT distance="100" swimtime="00:01:44.62" />
                    <SPLIT distance="125" swimtime="00:02:13.73" />
                    <SPLIT distance="150" swimtime="00:02:42.09" />
                    <SPLIT distance="175" swimtime="00:03:10.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-09-13" firstname="Mirosława" gender="F" lastname="Rajtar" nation="POL" license="503105600020" athleteid="108061">
              <RESULTS>
                <RESULT eventid="98777" points="218" reactiontime="+106" swimtime="00:00:38.58" resultid="108062" heatid="110588" lane="2" entrytime="00:00:38.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="167" swimtime="00:00:46.53" resultid="108063" heatid="110647" lane="3" entrytime="00:00:47.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="193" reactiontime="+106" swimtime="00:01:37.94" resultid="108064" heatid="110691" lane="3" entrytime="00:01:39.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.25" />
                    <SPLIT distance="50" swimtime="00:00:46.32" />
                    <SPLIT distance="75" swimtime="00:01:14.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="162" swimtime="00:00:44.72" resultid="108065" heatid="110737" lane="9" entrytime="00:00:46.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="170" reactiontime="+108" swimtime="00:03:19.69" resultid="108066" heatid="110765" lane="1" entrytime="00:03:21.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.37" />
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                    <SPLIT distance="75" swimtime="00:01:06.15" />
                    <SPLIT distance="100" swimtime="00:01:31.60" />
                    <SPLIT distance="125" swimtime="00:01:58.40" />
                    <SPLIT distance="150" swimtime="00:02:25.74" />
                    <SPLIT distance="175" swimtime="00:02:53.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="180" swimtime="00:00:50.92" resultid="108067" heatid="110818" lane="4" entrytime="00:00:54.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" license="503105600029" athleteid="108038">
              <RESULTS>
                <RESULT eventid="98777" points="330" reactiontime="+76" swimtime="00:00:33.61" resultid="108039" heatid="110590" lane="0" entrytime="00:00:33.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="272" swimtime="00:03:07.92" resultid="108040" heatid="110616" lane="4" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.44" />
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="75" swimtime="00:01:04.36" />
                    <SPLIT distance="100" swimtime="00:01:29.14" />
                    <SPLIT distance="125" swimtime="00:01:54.63" />
                    <SPLIT distance="150" swimtime="00:02:20.92" />
                    <SPLIT distance="175" swimtime="00:02:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="329" swimtime="00:01:13.73" resultid="108041" heatid="110675" lane="9" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.75" />
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="75" swimtime="00:00:54.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="324" reactiontime="+66" swimtime="00:01:22.47" resultid="108042" heatid="110693" lane="7" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.09" />
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="75" swimtime="00:01:02.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="317" reactiontime="+87" swimtime="00:01:31.38" resultid="108043" heatid="110724" lane="2" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.91" />
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                    <SPLIT distance="75" swimtime="00:01:06.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="284" swimtime="00:02:48.52" resultid="108044" heatid="110766" lane="9" entrytime="00:02:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.11" />
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="75" swimtime="00:00:58.67" />
                    <SPLIT distance="100" swimtime="00:01:20.38" />
                    <SPLIT distance="125" swimtime="00:01:42.61" />
                    <SPLIT distance="150" swimtime="00:02:05.19" />
                    <SPLIT distance="175" swimtime="00:02:27.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="368" swimtime="00:00:40.16" resultid="108045" heatid="110822" lane="9" entrytime="00:00:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" status="DNS" swimtime="00:00:00.00" resultid="108046" heatid="110840" lane="4" entrytime="00:05:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="503105700036" athleteid="108047">
              <RESULTS>
                <RESULT eventid="98798" points="500" reactiontime="+95" swimtime="00:00:25.52" resultid="108048" heatid="110607" lane="3" entrytime="00:00:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="400" swimtime="00:02:28.73" resultid="108049" heatid="110627" lane="9" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="75" swimtime="00:00:50.25" />
                    <SPLIT distance="100" swimtime="00:01:09.01" />
                    <SPLIT distance="125" swimtime="00:01:30.79" />
                    <SPLIT distance="150" swimtime="00:01:53.18" />
                    <SPLIT distance="175" swimtime="00:02:12.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="403" reactiontime="+79" swimtime="00:00:30.08" resultid="108050" heatid="110658" lane="4" entrytime="00:00:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="476" reactiontime="+82" swimtime="00:01:04.86" resultid="108051" heatid="110704" lane="5" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.10" />
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="75" swimtime="00:00:47.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="444" reactiontime="+89" swimtime="00:00:28.56" resultid="108052" heatid="110747" lane="3" entrytime="00:00:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="371" reactiontime="+82" swimtime="00:01:08.05" resultid="108053" heatid="110762" lane="3" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.92" />
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="75" swimtime="00:00:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="400" reactiontime="+84" swimtime="00:01:05.71" resultid="108054" heatid="110803" lane="8" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="75" swimtime="00:00:46.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="485" swimtime="00:00:32.12" resultid="108055" heatid="110833" lane="6" entrytime="00:00:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="108077">
              <RESULTS>
                <RESULT eventid="98814" points="415" reactiontime="+85" swimtime="00:02:43.27" resultid="108078" heatid="110617" lane="5" entrytime="00:02:49.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.51" />
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="75" swimtime="00:00:54.30" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="125" swimtime="00:01:38.59" />
                    <SPLIT distance="150" swimtime="00:02:02.84" />
                    <SPLIT distance="175" swimtime="00:02:23.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="432" reactiontime="+85" swimtime="00:01:14.96" resultid="108079" heatid="110695" lane="7" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="75" swimtime="00:00:56.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="423" swimtime="00:00:32.47" resultid="108080" heatid="110740" lane="9" entrytime="00:00:32.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="413" swimtime="00:01:13.30" resultid="108081" heatid="110796" lane="2" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.77" />
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="75" swimtime="00:00:53.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" license="503105700050" athleteid="108068">
              <RESULTS>
                <RESULT eventid="98798" points="146" swimtime="00:00:38.45" resultid="108069" heatid="110597" lane="9" entrytime="00:00:40.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="74" swimtime="00:04:20.97" resultid="108070" heatid="110620" lane="9" entrytime="00:04:11.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.90" />
                    <SPLIT distance="50" swimtime="00:00:55.07" />
                    <SPLIT distance="75" swimtime="00:01:30.29" />
                    <SPLIT distance="100" swimtime="00:02:07.23" />
                    <SPLIT distance="125" swimtime="00:02:45.42" />
                    <SPLIT distance="150" swimtime="00:03:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="122" reactiontime="+88" swimtime="00:01:30.54" resultid="108071" heatid="110679" lane="3" entrytime="00:01:30.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                    <SPLIT distance="75" swimtime="00:01:08.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="55" reactiontime="+104" swimtime="00:04:43.91" resultid="108072" heatid="110710" lane="8" entrytime="00:04:54.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.79" />
                    <SPLIT distance="50" swimtime="00:00:59.21" />
                    <SPLIT distance="75" swimtime="00:01:35.27" />
                    <SPLIT distance="100" swimtime="00:02:12.67" />
                    <SPLIT distance="125" swimtime="00:02:50.61" />
                    <SPLIT distance="150" swimtime="00:03:29.05" />
                    <SPLIT distance="175" swimtime="00:04:07.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="99" reactiontime="+94" swimtime="00:03:34.77" resultid="108073" heatid="110770" lane="1" entrytime="00:03:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.72" />
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="79" reactiontime="+81" swimtime="00:09:08.62" resultid="108074" heatid="110788" lane="7" entrytime="00:09:24.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.12" />
                    <SPLIT distance="50" swimtime="00:00:59.07" />
                    <SPLIT distance="75" swimtime="00:01:35.25" />
                    <SPLIT distance="100" swimtime="00:02:13.24" />
                    <SPLIT distance="125" swimtime="00:02:52.15" />
                    <SPLIT distance="150" swimtime="00:03:28.42" />
                    <SPLIT distance="175" swimtime="00:05:21.07" />
                    <SPLIT distance="200" swimtime="00:04:40.29" />
                    <SPLIT distance="225" swimtime="00:06:37.86" />
                    <SPLIT distance="250" swimtime="00:05:59.50" />
                    <SPLIT distance="275" swimtime="00:07:46.06" />
                    <SPLIT distance="300" swimtime="00:07:16.03" />
                    <SPLIT distance="325" swimtime="00:08:45.49" />
                    <SPLIT distance="350" swimtime="00:09:08.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="50" swimtime="00:02:11.12" resultid="108075" heatid="110798" lane="2" entrytime="00:02:05.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.15" />
                    <SPLIT distance="50" swimtime="00:00:58.74" />
                    <SPLIT distance="75" swimtime="00:01:35.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="90" reactiontime="+93" swimtime="00:07:52.97" resultid="108076" heatid="110851" lane="8" entrytime="00:07:54.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                    <SPLIT distance="75" swimtime="00:01:21.48" />
                    <SPLIT distance="100" swimtime="00:01:51.77" />
                    <SPLIT distance="125" swimtime="00:02:22.45" />
                    <SPLIT distance="225" swimtime="00:04:26.22" />
                    <SPLIT distance="325" swimtime="00:06:30.45" />
                    <SPLIT distance="375" swimtime="00:07:29.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="344" reactiontime="+66" swimtime="00:02:09.14" resultid="108105" heatid="110718" lane="8" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                    <SPLIT distance="75" swimtime="00:00:45.81" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="125" swimtime="00:01:18.30" />
                    <SPLIT distance="150" swimtime="00:01:35.69" />
                    <SPLIT distance="175" swimtime="00:01:51.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108056" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="108047" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="108020" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="108029" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="336" swimtime="00:01:58.74" resultid="108106" heatid="110783" lane="0" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="75" swimtime="00:00:43.75" />
                    <SPLIT distance="100" swimtime="00:01:01.85" />
                    <SPLIT distance="125" swimtime="00:01:17.04" />
                    <SPLIT distance="150" swimtime="00:01:33.63" />
                    <SPLIT distance="175" swimtime="00:01:45.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108047" number="1" />
                    <RELAYPOSITION athleteid="108056" number="2" />
                    <RELAYPOSITION athleteid="108029" number="3" />
                    <RELAYPOSITION athleteid="108020" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="412" reactiontime="+75" swimtime="00:02:19.74" resultid="108103" heatid="110715" lane="5" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.57" />
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                    <SPLIT distance="75" swimtime="00:00:51.81" />
                    <SPLIT distance="100" swimtime="00:01:13.54" />
                    <SPLIT distance="125" swimtime="00:01:28.70" />
                    <SPLIT distance="150" swimtime="00:01:46.55" />
                    <SPLIT distance="175" swimtime="00:02:02.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108082" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="108038" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="108077" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="108012" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99234" points="408" reactiontime="+83" swimtime="00:02:07.01" resultid="108104" heatid="110780" lane="5" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.00" />
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="75" swimtime="00:00:46.83" />
                    <SPLIT distance="100" swimtime="00:01:03.78" />
                    <SPLIT distance="125" swimtime="00:01:19.70" />
                    <SPLIT distance="150" swimtime="00:01:36.86" />
                    <SPLIT distance="175" swimtime="00:01:51.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108077" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="108012" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="108038" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="108082" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="361" reactiontime="+58" swimtime="00:01:55.93" resultid="108097" heatid="110631" lane="4" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.10" />
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                    <SPLIT distance="75" swimtime="00:00:42.34" />
                    <SPLIT distance="100" swimtime="00:00:58.54" />
                    <SPLIT distance="125" swimtime="00:01:12.49" />
                    <SPLIT distance="150" swimtime="00:01:28.60" />
                    <SPLIT distance="175" swimtime="00:01:41.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108056" number="1" reactiontime="+58" />
                    <RELAYPOSITION athleteid="108077" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="108082" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="108047" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="367" reactiontime="+66" swimtime="00:02:06.36" resultid="108098" heatid="110838" lane="7" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.14" />
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="75" swimtime="00:00:45.89" />
                    <SPLIT distance="100" swimtime="00:01:03.12" />
                    <SPLIT distance="125" swimtime="00:01:18.49" />
                    <SPLIT distance="150" swimtime="00:01:36.14" />
                    <SPLIT distance="175" swimtime="00:01:50.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108056" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="108047" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="108077" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="108082" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="282" reactiontime="+75" swimtime="00:02:05.87" resultid="108099" heatid="110630" lane="4" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                    <SPLIT distance="50" swimtime="00:00:25.56" />
                    <SPLIT distance="75" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:00:58.88" />
                    <SPLIT distance="125" swimtime="00:01:15.30" />
                    <SPLIT distance="150" swimtime="00:01:33.00" />
                    <SPLIT distance="175" swimtime="00:01:49.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106439" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="108012" number="2" />
                    <RELAYPOSITION athleteid="108029" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="108038" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="232" reactiontime="+82" swimtime="00:02:27.12" resultid="108100" heatid="110836" lane="4" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.53" />
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                    <SPLIT distance="75" swimtime="00:00:58.10" />
                    <SPLIT distance="100" swimtime="00:01:20.16" />
                    <SPLIT distance="125" swimtime="00:01:35.63" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                    <SPLIT distance="175" swimtime="00:02:09.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108012" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="108038" number="2" />
                    <RELAYPOSITION athleteid="108020" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="108029" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="98846" points="168" reactiontime="+118" swimtime="00:02:29.61" resultid="108101" heatid="110630" lane="0" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.17" />
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="75" swimtime="00:00:56.53" />
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="125" swimtime="00:01:36.24" />
                    <SPLIT distance="150" swimtime="00:01:58.77" />
                    <SPLIT distance="175" swimtime="00:02:13.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108061" number="1" reactiontime="+118" />
                    <RELAYPOSITION athleteid="108007" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="108090" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="108020" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="137" reactiontime="+77" swimtime="00:02:55.55" resultid="108102" heatid="110836" lane="7" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.48" />
                    <SPLIT distance="50" swimtime="00:00:46.03" />
                    <SPLIT distance="75" swimtime="00:01:04.52" />
                    <SPLIT distance="100" swimtime="00:01:25.75" />
                    <SPLIT distance="125" swimtime="00:01:49.13" />
                    <SPLIT distance="150" swimtime="00:02:17.07" />
                    <SPLIT distance="175" swimtime="00:02:35.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108061" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="108007" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="108090" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="108068" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="108188" name="Vandenynas">
          <CONTACT city="KOWNO" email="audrius.maske@gmail.com" name="Audrius Kiauke" phone="+37068697440" street="Taikos pr.61-39" zip="LT-50433" />
          <ATHLETES>
            <ATHLETE birthdate="1962-08-11" firstname="Kiauke" gender="M" lastname="Audrius" nation="LTU" athleteid="108189">
              <RESULTS>
                <RESULT eventid="98798" points="231" reactiontime="+85" swimtime="00:00:33.00" resultid="108918" heatid="110600" lane="5" entrytime="00:00:33.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="203" reactiontime="+72" swimtime="00:02:48.92" resultid="108919" heatid="110772" lane="2" entrytime="00:02:47.16">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.90" />
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="75" swimtime="00:00:57.65" />
                    <SPLIT distance="100" swimtime="00:01:19.14" />
                    <SPLIT distance="125" swimtime="00:01:41.84" />
                    <SPLIT distance="150" swimtime="00:02:04.72" />
                    <SPLIT distance="175" swimtime="00:02:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="230" reactiontime="+101" swimtime="00:01:13.25" resultid="108920" heatid="110681" lane="3" entrytime="00:01:14.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.36" />
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="75" swimtime="00:00:53.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="192" reactiontime="+81" swimtime="00:06:07.66" resultid="108921" heatid="110848" lane="8" entrytime="00:05:58.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.17" />
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="75" swimtime="00:01:00.97" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="125" swimtime="00:01:46.69" />
                    <SPLIT distance="150" swimtime="00:02:10.17" />
                    <SPLIT distance="175" swimtime="00:02:34.07" />
                    <SPLIT distance="200" swimtime="00:02:57.50" />
                    <SPLIT distance="225" swimtime="00:03:21.38" />
                    <SPLIT distance="250" swimtime="00:03:45.76" />
                    <SPLIT distance="275" swimtime="00:04:09.55" />
                    <SPLIT distance="300" swimtime="00:04:33.43" />
                    <SPLIT distance="325" swimtime="00:04:57.65" />
                    <SPLIT distance="350" swimtime="00:05:21.97" />
                    <SPLIT distance="375" swimtime="00:05:45.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="109056" name="Victory Masters Elbląg">
          <CONTACT city="Elbląg" email="lateccy@o2.pl" name="Latecki Grzegorz" phone="606147184" state="WARM-" street="Łokietka 45" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner-Mateusiak" nation="POL" athleteid="109083">
              <RESULTS>
                <RESULT eventid="98863" points="60" reactiontime="+128" swimtime="00:20:18.90" resultid="109591" heatid="110634" lane="8" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.94" />
                    <SPLIT distance="50" swimtime="00:01:00.47" />
                    <SPLIT distance="75" swimtime="00:01:36.78" />
                    <SPLIT distance="100" swimtime="00:02:13.88" />
                    <SPLIT distance="125" swimtime="00:02:51.32" />
                    <SPLIT distance="150" swimtime="00:03:29.43" />
                    <SPLIT distance="175" swimtime="00:04:07.17" />
                    <SPLIT distance="225" swimtime="00:05:23.67" />
                    <SPLIT distance="275" swimtime="00:06:42.93" />
                    <SPLIT distance="300" swimtime="00:07:22.50" />
                    <SPLIT distance="325" swimtime="00:08:01.90" />
                    <SPLIT distance="375" swimtime="00:09:20.45" />
                    <SPLIT distance="400" swimtime="00:09:59.93" />
                    <SPLIT distance="425" swimtime="00:10:38.76" />
                    <SPLIT distance="450" swimtime="00:11:16.51" />
                    <SPLIT distance="475" swimtime="00:11:55.80" />
                    <SPLIT distance="500" swimtime="00:12:34.93" />
                    <SPLIT distance="525" swimtime="00:13:12.92" />
                    <SPLIT distance="575" swimtime="00:14:31.38" />
                    <SPLIT distance="600" swimtime="00:15:10.87" />
                    <SPLIT distance="625" swimtime="00:15:49.56" />
                    <SPLIT distance="675" swimtime="00:17:06.82" />
                    <SPLIT distance="700" swimtime="00:17:45.67" />
                    <SPLIT distance="725" swimtime="00:18:23.11" />
                    <SPLIT distance="750" swimtime="00:19:01.35" />
                    <SPLIT distance="775" swimtime="00:19:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="53" swimtime="00:10:21.91" resultid="109592" heatid="110842" lane="0" entrytime="00:09:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.62" />
                    <SPLIT distance="50" swimtime="00:01:02.62" />
                    <SPLIT distance="75" swimtime="00:01:38.09" />
                    <SPLIT distance="100" swimtime="00:02:16.39" />
                    <SPLIT distance="125" swimtime="00:02:53.71" />
                    <SPLIT distance="150" swimtime="00:03:31.81" />
                    <SPLIT distance="175" swimtime="00:04:09.25" />
                    <SPLIT distance="200" swimtime="00:04:49.05" />
                    <SPLIT distance="225" swimtime="00:05:26.48" />
                    <SPLIT distance="250" swimtime="00:06:06.03" />
                    <SPLIT distance="275" swimtime="00:06:45.14" />
                    <SPLIT distance="300" swimtime="00:07:25.34" />
                    <SPLIT distance="325" swimtime="00:08:06.46" />
                    <SPLIT distance="350" swimtime="00:08:50.49" />
                    <SPLIT distance="375" swimtime="00:09:39.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98777" points="76" reactiontime="+113" swimtime="00:00:54.81" resultid="110354" heatid="110586" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="55" reactiontime="+88" swimtime="00:01:07.33" resultid="110355" heatid="110646" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="61" reactiontime="+126" swimtime="00:05:40.32" resultid="110356" heatid="110661" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.44" />
                    <SPLIT distance="50" swimtime="00:01:18.05" />
                    <SPLIT distance="75" swimtime="00:01:59.53" />
                    <SPLIT distance="100" swimtime="00:02:42.60" />
                    <SPLIT distance="125" swimtime="00:03:31.69" />
                    <SPLIT distance="150" swimtime="00:04:15.66" />
                    <SPLIT distance="175" swimtime="00:04:58.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="59" reactiontime="+117" swimtime="00:02:39.44" resultid="110357" heatid="110721" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.83" />
                    <SPLIT distance="50" swimtime="00:01:18.07" />
                    <SPLIT distance="75" swimtime="00:01:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="52" reactiontime="+92" swimtime="00:02:27.34" resultid="110358" heatid="110753" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.52" />
                    <SPLIT distance="50" swimtime="00:01:10.20" />
                    <SPLIT distance="75" swimtime="00:01:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="54" reactiontime="+86" swimtime="00:05:14.88" resultid="110359" heatid="110806" lane="1" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.06" />
                    <SPLIT distance="50" swimtime="00:01:13.06" />
                    <SPLIT distance="75" swimtime="00:01:51.47" />
                    <SPLIT distance="100" swimtime="00:02:32.31" />
                    <SPLIT distance="125" swimtime="00:03:12.10" />
                    <SPLIT distance="150" swimtime="00:03:52.98" />
                    <SPLIT distance="175" swimtime="00:04:33.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-12" firstname="Grzegorz" gender="M" lastname="Latecki" nation="POL" athleteid="109057">
              <RESULTS>
                <RESULT eventid="98798" points="419" swimtime="00:00:27.07" resultid="109058" heatid="110606" lane="9" entrytime="00:00:28.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="367" reactiontime="+84" swimtime="00:02:33.04" resultid="109059" heatid="110624" lane="5" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.32" />
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="75" swimtime="00:00:52.12" />
                    <SPLIT distance="100" swimtime="00:01:11.24" />
                    <SPLIT distance="125" swimtime="00:01:33.96" />
                    <SPLIT distance="150" swimtime="00:01:56.93" />
                    <SPLIT distance="175" swimtime="00:02:16.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="340" reactiontime="+72" swimtime="00:00:31.83" resultid="109060" heatid="110657" lane="0" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="397" reactiontime="+90" swimtime="00:01:08.92" resultid="109061" heatid="110702" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.74" />
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="75" swimtime="00:00:51.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="391" swimtime="00:00:29.80" resultid="109062" heatid="110748" lane="0" entrytime="00:00:30.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="324" reactiontime="+95" swimtime="00:05:42.75" resultid="109063" heatid="110790" lane="3" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.54" />
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="75" swimtime="00:00:57.54" />
                    <SPLIT distance="100" swimtime="00:01:19.59" />
                    <SPLIT distance="125" swimtime="00:01:41.40" />
                    <SPLIT distance="150" swimtime="00:02:03.70" />
                    <SPLIT distance="175" swimtime="00:02:25.95" />
                    <SPLIT distance="200" swimtime="00:02:47.73" />
                    <SPLIT distance="225" swimtime="00:03:11.54" />
                    <SPLIT distance="250" swimtime="00:03:36.31" />
                    <SPLIT distance="275" swimtime="00:04:00.84" />
                    <SPLIT distance="300" swimtime="00:04:26.25" />
                    <SPLIT distance="325" swimtime="00:04:45.90" />
                    <SPLIT distance="350" swimtime="00:05:05.46" />
                    <SPLIT distance="375" swimtime="00:05:24.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="348" reactiontime="+89" swimtime="00:01:08.85" resultid="109064" heatid="110802" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.29" />
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="75" swimtime="00:00:50.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="354" swimtime="00:00:35.67" resultid="109065" heatid="110829" lane="2" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="109079">
              <RESULTS>
                <RESULT eventid="98907" points="163" reactiontime="+106" swimtime="00:01:33.08" resultid="109080" heatid="110672" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.88" />
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                    <SPLIT distance="75" swimtime="00:01:09.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="149" reactiontime="+102" swimtime="00:03:28.71" resultid="109081" heatid="110765" lane="8" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.53" />
                    <SPLIT distance="50" swimtime="00:00:50.23" />
                    <SPLIT distance="75" swimtime="00:01:17.09" />
                    <SPLIT distance="100" swimtime="00:01:44.34" />
                    <SPLIT distance="125" swimtime="00:02:10.97" />
                    <SPLIT distance="150" swimtime="00:02:37.42" />
                    <SPLIT distance="175" swimtime="00:03:03.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="163" reactiontime="+115" swimtime="00:07:09.10" resultid="109082" heatid="110842" lane="2" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.82" />
                    <SPLIT distance="50" swimtime="00:00:49.81" />
                    <SPLIT distance="75" swimtime="00:01:16.82" />
                    <SPLIT distance="100" swimtime="00:01:44.32" />
                    <SPLIT distance="125" swimtime="00:02:12.06" />
                    <SPLIT distance="150" swimtime="00:02:39.48" />
                    <SPLIT distance="175" swimtime="00:03:06.85" />
                    <SPLIT distance="200" swimtime="00:03:34.88" />
                    <SPLIT distance="225" swimtime="00:04:02.64" />
                    <SPLIT distance="250" swimtime="00:04:30.19" />
                    <SPLIT distance="275" swimtime="00:04:57.16" />
                    <SPLIT distance="300" swimtime="00:05:24.30" />
                    <SPLIT distance="325" swimtime="00:05:50.92" />
                    <SPLIT distance="350" swimtime="00:06:18.23" />
                    <SPLIT distance="375" swimtime="00:06:44.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-06" firstname="Andrzej" gender="M" lastname="Pasieczny" nation="POL" athleteid="109066">
              <RESULTS>
                <RESULT eventid="98798" points="377" reactiontime="+90" swimtime="00:00:28.04" resultid="109067" heatid="110606" lane="3" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="415" reactiontime="+81" swimtime="00:02:25.45" resultid="109068" heatid="110713" lane="7" entrytime="00:02:27.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.32" />
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="75" swimtime="00:00:49.60" />
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                    <SPLIT distance="125" swimtime="00:01:26.80" />
                    <SPLIT distance="150" swimtime="00:01:46.03" />
                    <SPLIT distance="175" swimtime="00:02:05.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="464" swimtime="00:02:08.32" resultid="109069" heatid="110777" lane="9" entrytime="00:02:12.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.36" />
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="75" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:02.85" />
                    <SPLIT distance="125" swimtime="00:01:19.35" />
                    <SPLIT distance="150" swimtime="00:01:36.00" />
                    <SPLIT distance="175" swimtime="00:01:52.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="429" reactiontime="+88" swimtime="00:01:04.19" resultid="109070" heatid="110804" lane="3" entrytime="00:01:03.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="75" swimtime="00:00:46.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" reactiontime="+90" status="DNF" swimtime="00:00:00.00" resultid="109071" heatid="110843" lane="7" entrytime="00:04:31.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.92" />
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="75" swimtime="00:00:47.99" />
                    <SPLIT distance="100" swimtime="00:01:04.74" />
                    <SPLIT distance="125" swimtime="00:01:21.93" />
                    <SPLIT distance="150" swimtime="00:01:39.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-04" firstname="Karol" gender="M" lastname="Sosna" nation="POL" athleteid="109072">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="109073" heatid="110602" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="109074" heatid="110668" lane="0" entrytime="00:03:15.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="109075" heatid="110700" lane="8" entrytime="00:01:18.00" />
                <RESULT eventid="99091" points="293" swimtime="00:01:23.65" resultid="109076" heatid="110731" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.32" />
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="75" swimtime="00:01:01.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="219" reactiontime="+94" swimtime="00:00:36.12" resultid="109077" heatid="110744" lane="5" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="340" swimtime="00:00:36.17" resultid="109078" heatid="110831" lane="9" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WMT" nation="POL" region="MAZ" clubid="108724" name="Warsaw Masters Team">
          <CONTACT city="Warszawa" email="wojciech.kaluzynski@gmail.com" name="Wojciech Kałużyński" phone="607454444" state="MAZ" />
          <ATHLETES>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="109361">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="109362" heatid="110608" lane="5" entrytime="00:00:27.11" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="109363" heatid="110626" lane="9" entrytime="00:02:35.56" />
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="109364" heatid="110688" lane="8" entrytime="00:00:58.31" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="109365" heatid="110704" lane="9" entrytime="00:01:08.34" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="109366" heatid="110733" lane="8" entrytime="00:01:16.72" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="109367" heatid="110777" lane="0" entrytime="00:02:11.72" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="109368" heatid="110833" lane="8" entrytime="00:00:34.12" />
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="109369" heatid="110844" lane="8" entrytime="00:04:51.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="109344">
              <RESULTS>
                <RESULT eventid="98830" status="WDR" swimtime="00:00:00.00" resultid="109345" heatid="110619" lane="7" />
                <RESULT eventid="98956" status="WDR" swimtime="00:00:00.00" resultid="109346" heatid="110665" lane="6" />
                <RESULT eventid="98988" status="WDR" swimtime="00:00:00.00" resultid="109347" heatid="110696" lane="7" />
                <RESULT eventid="99091" status="WDR" swimtime="00:00:00.00" resultid="109348" heatid="110726" lane="4" />
                <RESULT eventid="99393" status="WDR" swimtime="00:00:00.00" resultid="109350" heatid="110810" lane="2" />
                <RESULT eventid="99425" status="WDR" swimtime="00:00:00.00" resultid="109351" heatid="110824" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-10-19" firstname="Emilia" gender="F" lastname="Sączyńska" nation="POL" athleteid="109421">
              <RESULTS>
                <RESULT eventid="106294" points="345" reactiontime="+84" swimtime="00:00:36.57" resultid="109422" heatid="110649" lane="3" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="343" reactiontime="+89" swimtime="00:01:20.90" resultid="109423" heatid="110694" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.37" />
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="75" swimtime="00:01:01.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="319" reactiontime="+82" swimtime="00:00:35.66" resultid="109424" heatid="110738" lane="5" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="347" reactiontime="+74" swimtime="00:01:18.30" resultid="109425" heatid="110756" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="75" swimtime="00:00:57.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="109426" heatid="110795" lane="5" entrytime="00:01:24.00" />
                <RESULT eventid="99377" status="DNS" swimtime="00:00:00.00" resultid="109427" heatid="110809" lane="7" entrytime="00:02:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-06" firstname="Mateusz" gender="M" lastname="Bednarz" nation="POL" athleteid="109352">
              <RESULTS>
                <RESULT eventid="98798" points="328" reactiontime="+89" swimtime="00:00:29.37" resultid="109353" heatid="110604" lane="6" entrytime="00:00:29.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="293" reactiontime="+86" swimtime="00:02:45.03" resultid="109354" heatid="110624" lane="8" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.57" />
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="75" swimtime="00:00:59.06" />
                    <SPLIT distance="100" swimtime="00:01:20.63" />
                    <SPLIT distance="125" swimtime="00:01:44.57" />
                    <SPLIT distance="150" swimtime="00:02:08.89" />
                    <SPLIT distance="175" swimtime="00:02:28.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="203" reactiontime="+92" swimtime="00:00:37.75" resultid="109355" heatid="110655" lane="0" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="322" reactiontime="+74" swimtime="00:01:13.84" resultid="109356" heatid="110700" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.90" />
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="75" swimtime="00:00:56.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="312" swimtime="00:00:32.13" resultid="109357" heatid="110745" lane="6" entrytime="00:00:32.84">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="349" reactiontime="+93" swimtime="00:02:21.13" resultid="109358" heatid="110774" lane="3" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.47" />
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="75" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:08.81" />
                    <SPLIT distance="125" swimtime="00:01:27.25" />
                    <SPLIT distance="150" swimtime="00:01:45.95" />
                    <SPLIT distance="175" swimtime="00:02:04.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="109359" heatid="110801" lane="0" entrytime="00:01:18.00" />
                <RESULT eventid="99473" points="350" reactiontime="+102" swimtime="00:05:01.02" resultid="109360" heatid="110846" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.61" />
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="75" swimtime="00:00:51.40" />
                    <SPLIT distance="100" swimtime="00:01:10.13" />
                    <SPLIT distance="125" swimtime="00:01:29.13" />
                    <SPLIT distance="150" swimtime="00:01:48.73" />
                    <SPLIT distance="175" swimtime="00:02:08.29" />
                    <SPLIT distance="200" swimtime="00:02:27.79" />
                    <SPLIT distance="225" swimtime="00:02:47.32" />
                    <SPLIT distance="250" swimtime="00:03:06.78" />
                    <SPLIT distance="275" swimtime="00:03:26.08" />
                    <SPLIT distance="300" swimtime="00:03:45.61" />
                    <SPLIT distance="325" swimtime="00:04:04.90" />
                    <SPLIT distance="350" swimtime="00:04:24.51" />
                    <SPLIT distance="375" swimtime="00:04:43.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-04-14" firstname="Wiesław" gender="M" lastname="Załuski" nation="POL" athleteid="109370">
              <RESULTS>
                <RESULT eventid="98830" points="241" reactiontime="+122" swimtime="00:02:56.14" resultid="109371" heatid="110622" lane="4" entrytime="00:03:00.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.82" />
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="75" swimtime="00:00:58.60" />
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="125" swimtime="00:01:47.27" />
                    <SPLIT distance="150" swimtime="00:02:13.89" />
                    <SPLIT distance="175" swimtime="00:02:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="247" reactiontime="+80" swimtime="00:00:35.38" resultid="109372" heatid="110655" lane="9" entrytime="00:00:38.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="276" swimtime="00:01:17.72" resultid="109373" heatid="110699" lane="0" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.31" />
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="75" swimtime="00:00:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="245" reactiontime="+73" swimtime="00:01:18.17" resultid="109374" heatid="110760" lane="9" entrytime="00:01:25.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.98" />
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="75" swimtime="00:00:57.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="214" reactiontime="+75" swimtime="00:02:56.51" resultid="109375" heatid="110813" lane="9" entrytime="00:03:07.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.93" />
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                    <SPLIT distance="75" swimtime="00:00:59.54" />
                    <SPLIT distance="100" swimtime="00:01:21.40" />
                    <SPLIT distance="125" swimtime="00:01:44.06" />
                    <SPLIT distance="150" swimtime="00:02:08.10" />
                    <SPLIT distance="175" swimtime="00:02:32.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="109433">
              <RESULTS>
                <RESULT eventid="98956" points="203" reactiontime="+100" swimtime="00:03:24.85" resultid="109434" heatid="110667" lane="8" entrytime="00:03:22.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.21" />
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="75" swimtime="00:01:09.70" />
                    <SPLIT distance="100" swimtime="00:01:35.74" />
                    <SPLIT distance="125" swimtime="00:02:02.07" />
                    <SPLIT distance="150" swimtime="00:02:29.41" />
                    <SPLIT distance="175" swimtime="00:02:57.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="109435" heatid="110710" lane="5" entrytime="00:03:54.45" />
                <RESULT eventid="99091" points="186" reactiontime="+105" swimtime="00:01:37.25" resultid="109436" heatid="110729" lane="3" entrytime="00:01:33.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.47" />
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="75" swimtime="00:01:10.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="117" reactiontime="+119" swimtime="00:01:39.02" resultid="109437" heatid="110799" lane="3" entrytime="00:01:38.46">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.30" />
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="75" swimtime="00:01:12.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="216" swimtime="00:00:42.04" resultid="109438" heatid="110827" lane="9" entrytime="00:00:42.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-18" firstname="Barbara" gender="F" lastname="Łowkis" nation="POL" athleteid="109451">
              <RESULTS>
                <RESULT eventid="98777" points="193" swimtime="00:00:40.19" resultid="109452" heatid="110588" lane="9" entrytime="00:00:39.69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="166" reactiontime="+78" swimtime="00:00:46.69" resultid="109453" heatid="110647" lane="6" entrytime="00:00:47.31">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="157" reactiontime="+107" swimtime="00:01:34.30" resultid="109454" heatid="110672" lane="7" entrytime="00:01:43.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="135" reactiontime="+84" swimtime="00:01:47.25" resultid="109455" heatid="110754" lane="0" entrytime="00:01:50.66" />
                <RESULT eventid="99377" points="121" reactiontime="+98" swimtime="00:04:00.55" resultid="109456" heatid="110807" lane="0" entrytime="00:04:02.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="109397">
              <RESULTS>
                <RESULT eventid="98798" points="374" reactiontime="+91" swimtime="00:00:28.10" resultid="109398" heatid="110602" lane="3" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="369" reactiontime="+82" swimtime="00:02:32.74" resultid="109399" heatid="110626" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.27" />
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="75" swimtime="00:00:52.61" />
                    <SPLIT distance="100" swimtime="00:01:11.75" />
                    <SPLIT distance="125" swimtime="00:01:34.95" />
                    <SPLIT distance="150" swimtime="00:01:58.09" />
                    <SPLIT distance="175" swimtime="00:02:16.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="375" reactiontime="+83" swimtime="00:00:30.79" resultid="109400" heatid="110659" lane="9" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="436" reactiontime="+87" swimtime="00:01:06.76" resultid="109401" heatid="110703" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.47" />
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="75" swimtime="00:00:51.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="379" reactiontime="+87" swimtime="00:01:07.56" resultid="109402" heatid="110762" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.81" />
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="75" swimtime="00:00:50.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="403" reactiontime="+63" swimtime="00:02:14.43" resultid="109403" heatid="110776" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.63" />
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="75" swimtime="00:00:48.40" />
                    <SPLIT distance="100" swimtime="00:01:05.77" />
                    <SPLIT distance="125" swimtime="00:01:23.11" />
                    <SPLIT distance="150" swimtime="00:01:40.85" />
                    <SPLIT distance="175" swimtime="00:01:58.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="376" swimtime="00:01:07.11" resultid="109404" heatid="110798" lane="0">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.06" />
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="75" swimtime="00:00:49.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="330" reactiontime="+84" swimtime="00:02:32.84" resultid="109405" heatid="110815" lane="3" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.90" />
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="75" swimtime="00:00:54.35" />
                    <SPLIT distance="100" swimtime="00:01:13.91" />
                    <SPLIT distance="125" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:01:53.98" />
                    <SPLIT distance="175" swimtime="00:02:13.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="109389">
              <RESULTS>
                <RESULT eventid="98798" points="137" reactiontime="+119" swimtime="00:00:39.24" resultid="109390" heatid="110597" lane="0" entrytime="00:00:40.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="142" swimtime="00:14:08.71" resultid="109391" heatid="110638" lane="4" entrytime="00:13:59.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.94" />
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                    <SPLIT distance="75" swimtime="00:01:10.22" />
                    <SPLIT distance="100" swimtime="00:01:36.23" />
                    <SPLIT distance="125" swimtime="00:02:02.85" />
                    <SPLIT distance="150" swimtime="00:02:29.75" />
                    <SPLIT distance="175" swimtime="00:02:57.08" />
                    <SPLIT distance="200" swimtime="00:03:23.85" />
                    <SPLIT distance="225" swimtime="00:03:51.88" />
                    <SPLIT distance="250" swimtime="00:04:18.57" />
                    <SPLIT distance="275" swimtime="00:04:45.98" />
                    <SPLIT distance="300" swimtime="00:05:12.39" />
                    <SPLIT distance="325" swimtime="00:05:39.67" />
                    <SPLIT distance="350" swimtime="00:06:06.12" />
                    <SPLIT distance="375" swimtime="00:06:32.92" />
                    <SPLIT distance="400" swimtime="00:06:59.41" />
                    <SPLIT distance="425" swimtime="00:07:26.26" />
                    <SPLIT distance="450" swimtime="00:07:53.10" />
                    <SPLIT distance="475" swimtime="00:09:14.68" />
                    <SPLIT distance="500" swimtime="00:08:47.22" />
                    <SPLIT distance="525" swimtime="00:10:10.42" />
                    <SPLIT distance="550" swimtime="00:09:42.99" />
                    <SPLIT distance="575" swimtime="00:11:04.76" />
                    <SPLIT distance="600" swimtime="00:10:37.51" />
                    <SPLIT distance="625" swimtime="00:11:59.00" />
                    <SPLIT distance="650" swimtime="00:11:31.57" />
                    <SPLIT distance="675" swimtime="00:12:52.93" />
                    <SPLIT distance="700" swimtime="00:12:25.73" />
                    <SPLIT distance="725" swimtime="00:13:45.43" />
                    <SPLIT distance="750" swimtime="00:13:19.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="66" reactiontime="+102" swimtime="00:00:54.96" resultid="109392" heatid="110652" lane="1" entrytime="00:00:56.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="137" reactiontime="+113" swimtime="00:01:27.00" resultid="109393" heatid="110680" lane="8" entrytime="00:01:27.19">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.90" />
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                    <SPLIT distance="75" swimtime="00:01:05.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="92" swimtime="00:00:48.23" resultid="109394" heatid="110742" lane="6" entrytime="00:00:48.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="146" reactiontime="+97" swimtime="00:03:08.32" resultid="109395" heatid="110770" lane="4" entrytime="00:03:08.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.97" />
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                    <SPLIT distance="75" swimtime="00:01:06.80" />
                    <SPLIT distance="100" swimtime="00:01:31.29" />
                    <SPLIT distance="125" swimtime="00:01:56.71" />
                    <SPLIT distance="150" swimtime="00:02:21.30" />
                    <SPLIT distance="175" swimtime="00:02:46.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="153" reactiontime="+114" swimtime="00:06:36.25" resultid="109396" heatid="110850" lane="5" entrytime="00:06:27.39">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.95" />
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                    <SPLIT distance="75" swimtime="00:01:10.76" />
                    <SPLIT distance="100" swimtime="00:01:36.52" />
                    <SPLIT distance="125" swimtime="00:03:45.75" />
                    <SPLIT distance="150" swimtime="00:02:28.25" />
                    <SPLIT distance="175" swimtime="00:06:14.88" />
                    <SPLIT distance="200" swimtime="00:03:19.92" />
                    <SPLIT distance="250" swimtime="00:05:00.56" />
                    <SPLIT distance="300" swimtime="00:05:50.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-22" firstname="Karol" gender="M" lastname="Dzięcioł" nation="POL" athleteid="109439">
              <RESULTS>
                <RESULT eventid="98798" points="500" reactiontime="+80" swimtime="00:00:25.52" resultid="109440" heatid="110611" lane="2" entrytime="00:00:25.64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="495" reactiontime="+79" swimtime="00:00:56.81" resultid="109441" heatid="110688" lane="3" entrytime="00:00:56.85">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.68" />
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                    <SPLIT distance="75" swimtime="00:00:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="449" reactiontime="+73" swimtime="00:01:06.13" resultid="109442" heatid="110705" lane="7" entrytime="00:01:05.85">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.60" />
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="75" swimtime="00:00:50.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="436" reactiontime="+79" swimtime="00:02:11.00" resultid="109443" heatid="110776" lane="3" entrytime="00:02:14.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="75" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:02.33" />
                    <SPLIT distance="125" swimtime="00:01:19.38" />
                    <SPLIT distance="150" swimtime="00:01:36.96" />
                    <SPLIT distance="175" swimtime="00:01:54.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="109444" heatid="110804" lane="7" entrytime="00:01:06.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="109445">
              <RESULTS>
                <RESULT eventid="98940" points="359" reactiontime="+75" swimtime="00:03:09.30" resultid="109446" heatid="110664" lane="8" entrytime="00:03:08.59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.23" />
                    <SPLIT distance="50" swimtime="00:00:43.81" />
                    <SPLIT distance="75" swimtime="00:01:07.63" />
                    <SPLIT distance="100" swimtime="00:01:31.79" />
                    <SPLIT distance="125" swimtime="00:01:55.87" />
                    <SPLIT distance="150" swimtime="00:02:20.51" />
                    <SPLIT distance="175" swimtime="00:02:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="371" reactiontime="+84" swimtime="00:01:26.75" resultid="109447" heatid="110724" lane="3" entrytime="00:01:27.16">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.06" />
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                    <SPLIT distance="75" swimtime="00:01:03.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="289" swimtime="00:02:47.48" resultid="109448" heatid="110767" lane="0" entrytime="00:02:45.81">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.72" />
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="75" swimtime="00:00:58.99" />
                    <SPLIT distance="100" swimtime="00:01:21.11" />
                    <SPLIT distance="125" swimtime="00:01:42.73" />
                    <SPLIT distance="150" swimtime="00:02:04.82" />
                    <SPLIT distance="175" swimtime="00:02:26.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="353" reactiontime="+80" swimtime="00:00:40.72" resultid="109449" heatid="110821" lane="5" entrytime="00:00:40.28">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="305" reactiontime="+77" swimtime="00:05:48.16" resultid="109450" heatid="110840" lane="8" entrytime="00:05:50.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.27" />
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                    <SPLIT distance="75" swimtime="00:01:01.56" />
                    <SPLIT distance="100" swimtime="00:01:24.47" />
                    <SPLIT distance="125" swimtime="00:01:47.06" />
                    <SPLIT distance="150" swimtime="00:02:09.74" />
                    <SPLIT distance="175" swimtime="00:02:32.16" />
                    <SPLIT distance="200" swimtime="00:02:55.05" />
                    <SPLIT distance="225" swimtime="00:03:16.50" />
                    <SPLIT distance="250" swimtime="00:03:38.13" />
                    <SPLIT distance="275" swimtime="00:03:59.69" />
                    <SPLIT distance="300" swimtime="00:04:21.88" />
                    <SPLIT distance="325" swimtime="00:04:43.79" />
                    <SPLIT distance="350" swimtime="00:05:06.16" />
                    <SPLIT distance="375" swimtime="00:05:27.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-28" firstname="Paweł" gender="M" lastname="Rogosz" nation="POL" athleteid="109336">
              <RESULTS>
                <RESULT eventid="98830" points="370" reactiontime="+92" swimtime="00:02:32.62" resultid="109337" heatid="110625" lane="4" entrytime="00:02:35.79">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.27" />
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="75" swimtime="00:00:54.87" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="125" swimtime="00:01:36.23" />
                    <SPLIT distance="150" swimtime="00:01:57.83" />
                    <SPLIT distance="175" swimtime="00:02:15.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="328" reactiontime="+104" swimtime="00:10:42.77" resultid="109338" heatid="110635" lane="0" entrytime="00:10:41.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.54" />
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="75" swimtime="00:00:54.42" />
                    <SPLIT distance="100" swimtime="00:01:14.48" />
                    <SPLIT distance="125" swimtime="00:01:34.79" />
                    <SPLIT distance="150" swimtime="00:01:55.08" />
                    <SPLIT distance="175" swimtime="00:02:15.50" />
                    <SPLIT distance="200" swimtime="00:02:35.79" />
                    <SPLIT distance="225" swimtime="00:02:56.62" />
                    <SPLIT distance="250" swimtime="00:03:17.25" />
                    <SPLIT distance="275" swimtime="00:03:38.12" />
                    <SPLIT distance="300" swimtime="00:03:58.71" />
                    <SPLIT distance="325" swimtime="00:04:19.17" />
                    <SPLIT distance="350" swimtime="00:04:39.59" />
                    <SPLIT distance="375" swimtime="00:05:00.16" />
                    <SPLIT distance="400" swimtime="00:05:20.67" />
                    <SPLIT distance="425" swimtime="00:05:41.06" />
                    <SPLIT distance="450" swimtime="00:06:01.34" />
                    <SPLIT distance="475" swimtime="00:06:21.63" />
                    <SPLIT distance="500" swimtime="00:06:41.91" />
                    <SPLIT distance="525" swimtime="00:07:02.31" />
                    <SPLIT distance="550" swimtime="00:07:22.80" />
                    <SPLIT distance="575" swimtime="00:07:43.12" />
                    <SPLIT distance="600" swimtime="00:08:03.77" />
                    <SPLIT distance="625" swimtime="00:08:23.80" />
                    <SPLIT distance="650" swimtime="00:08:44.12" />
                    <SPLIT distance="675" swimtime="00:09:04.57" />
                    <SPLIT distance="700" swimtime="00:09:24.82" />
                    <SPLIT distance="725" swimtime="00:09:44.75" />
                    <SPLIT distance="750" swimtime="00:10:04.44" />
                    <SPLIT distance="775" swimtime="00:10:24.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="381" reactiontime="+97" swimtime="00:02:46.18" resultid="109339" heatid="110669" lane="6" entrytime="00:02:55.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.30" />
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="75" swimtime="00:00:58.88" />
                    <SPLIT distance="100" swimtime="00:01:20.34" />
                    <SPLIT distance="125" swimtime="00:01:41.66" />
                    <SPLIT distance="150" swimtime="00:02:03.12" />
                    <SPLIT distance="175" swimtime="00:02:24.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="315" reactiontime="+97" swimtime="00:02:39.54" resultid="109340" heatid="110712" lane="4" entrytime="00:02:45.79">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.20" />
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="75" swimtime="00:00:56.30" />
                    <SPLIT distance="100" swimtime="00:01:17.21" />
                    <SPLIT distance="125" swimtime="00:01:37.51" />
                    <SPLIT distance="150" swimtime="00:01:58.26" />
                    <SPLIT distance="175" swimtime="00:02:18.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="109341" heatid="110791" lane="3" entrytime="00:05:39.32" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="109342" heatid="110813" lane="2" entrytime="00:02:55.79" />
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="109343" heatid="110846" lane="2" entrytime="00:05:14.79" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="109412">
              <RESULTS>
                <RESULT eventid="98798" points="148" reactiontime="+75" swimtime="00:00:38.28" resultid="109413" heatid="110598" lane="5" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="104" swimtime="00:15:41.35" resultid="109414" heatid="110638" lane="1" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.31" />
                    <SPLIT distance="50" swimtime="00:00:50.59" />
                    <SPLIT distance="75" swimtime="00:01:18.97" />
                    <SPLIT distance="100" swimtime="00:01:47.81" />
                    <SPLIT distance="125" swimtime="00:02:16.36" />
                    <SPLIT distance="150" swimtime="00:02:46.49" />
                    <SPLIT distance="175" swimtime="00:03:15.72" />
                    <SPLIT distance="200" swimtime="00:03:46.38" />
                    <SPLIT distance="225" swimtime="00:04:16.85" />
                    <SPLIT distance="250" swimtime="00:04:47.81" />
                    <SPLIT distance="275" swimtime="00:05:17.88" />
                    <SPLIT distance="300" swimtime="00:05:49.06" />
                    <SPLIT distance="325" swimtime="00:06:20.06" />
                    <SPLIT distance="350" swimtime="00:06:51.67" />
                    <SPLIT distance="375" swimtime="00:07:21.79" />
                    <SPLIT distance="400" swimtime="00:07:52.56" />
                    <SPLIT distance="425" swimtime="00:08:23.26" />
                    <SPLIT distance="450" swimtime="00:08:53.56" />
                    <SPLIT distance="475" swimtime="00:09:24.01" />
                    <SPLIT distance="500" swimtime="00:09:53.84" />
                    <SPLIT distance="525" swimtime="00:10:23.24" />
                    <SPLIT distance="550" swimtime="00:10:52.89" />
                    <SPLIT distance="575" swimtime="00:11:23.24" />
                    <SPLIT distance="600" swimtime="00:11:52.83" />
                    <SPLIT distance="625" swimtime="00:12:23.01" />
                    <SPLIT distance="650" swimtime="00:12:53.38" />
                    <SPLIT distance="675" swimtime="00:13:23.15" />
                    <SPLIT distance="700" swimtime="00:13:52.63" />
                    <SPLIT distance="725" swimtime="00:14:21.48" />
                    <SPLIT distance="750" swimtime="00:14:50.60" />
                    <SPLIT distance="775" swimtime="00:15:17.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="85" reactiontime="+81" swimtime="00:00:50.46" resultid="109415" heatid="110652" lane="4" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="138" reactiontime="+72" swimtime="00:01:26.96" resultid="109416" heatid="110680" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.66" />
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="75" swimtime="00:01:03.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="80" reactiontime="+91" swimtime="00:01:53.23" resultid="109417" heatid="110758" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.57" />
                    <SPLIT distance="50" swimtime="00:00:55.46" />
                    <SPLIT distance="75" swimtime="00:01:24.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="115" swimtime="00:03:24.17" resultid="109418" heatid="110770" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="75" swimtime="00:01:04.66" />
                    <SPLIT distance="100" swimtime="00:01:31.46" />
                    <SPLIT distance="125" swimtime="00:02:00.43" />
                    <SPLIT distance="150" swimtime="00:02:29.34" />
                    <SPLIT distance="175" swimtime="00:02:57.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="75" reactiontime="+98" swimtime="00:04:09.39" resultid="109419" heatid="110811" lane="1" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.20" />
                    <SPLIT distance="50" swimtime="00:00:57.23" />
                    <SPLIT distance="75" swimtime="00:01:28.99" />
                    <SPLIT distance="100" swimtime="00:02:01.13" />
                    <SPLIT distance="125" swimtime="00:02:32.95" />
                    <SPLIT distance="150" swimtime="00:03:05.94" />
                    <SPLIT distance="175" swimtime="00:03:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="97" reactiontime="+77" swimtime="00:07:41.31" resultid="109420" heatid="110851" lane="3" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.36" />
                    <SPLIT distance="50" swimtime="00:00:46.23" />
                    <SPLIT distance="75" swimtime="00:01:13.34" />
                    <SPLIT distance="100" swimtime="00:01:40.80" />
                    <SPLIT distance="125" swimtime="00:02:09.69" />
                    <SPLIT distance="150" swimtime="00:02:39.07" />
                    <SPLIT distance="175" swimtime="00:03:08.29" />
                    <SPLIT distance="200" swimtime="00:03:37.12" />
                    <SPLIT distance="225" swimtime="00:04:08.31" />
                    <SPLIT distance="250" swimtime="00:04:38.27" />
                    <SPLIT distance="275" swimtime="00:05:10.22" />
                    <SPLIT distance="300" swimtime="00:05:41.51" />
                    <SPLIT distance="325" swimtime="00:06:13.50" />
                    <SPLIT distance="350" swimtime="00:06:44.38" />
                    <SPLIT distance="375" swimtime="00:07:17.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="109428">
              <RESULTS>
                <RESULT eventid="98777" points="101" swimtime="00:00:49.89" resultid="109429" heatid="110586" lane="5" entrytime="00:00:48.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="116" swimtime="00:16:21.50" resultid="109430" heatid="110634" lane="1" entrytime="00:16:12.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.03" />
                    <SPLIT distance="50" swimtime="00:00:53.32" />
                    <SPLIT distance="75" swimtime="00:01:23.44" />
                    <SPLIT distance="100" swimtime="00:01:54.74" />
                    <SPLIT distance="125" swimtime="00:02:26.45" />
                    <SPLIT distance="150" swimtime="00:02:58.22" />
                    <SPLIT distance="175" swimtime="00:03:30.10" />
                    <SPLIT distance="200" swimtime="00:04:01.59" />
                    <SPLIT distance="225" swimtime="00:04:33.66" />
                    <SPLIT distance="250" swimtime="00:05:05.22" />
                    <SPLIT distance="275" swimtime="00:05:37.20" />
                    <SPLIT distance="300" swimtime="00:06:08.36" />
                    <SPLIT distance="325" swimtime="00:06:39.20" />
                    <SPLIT distance="350" swimtime="00:07:11.23" />
                    <SPLIT distance="375" swimtime="00:07:41.87" />
                    <SPLIT distance="400" swimtime="00:08:12.69" />
                    <SPLIT distance="425" swimtime="00:08:44.17" />
                    <SPLIT distance="450" swimtime="00:09:15.26" />
                    <SPLIT distance="475" swimtime="00:09:46.07" />
                    <SPLIT distance="500" swimtime="00:10:17.42" />
                    <SPLIT distance="525" swimtime="00:10:47.77" />
                    <SPLIT distance="550" swimtime="00:11:18.81" />
                    <SPLIT distance="575" swimtime="00:11:49.13" />
                    <SPLIT distance="600" swimtime="00:12:19.04" />
                    <SPLIT distance="625" swimtime="00:12:51.22" />
                    <SPLIT distance="650" swimtime="00:13:21.00" />
                    <SPLIT distance="675" swimtime="00:13:52.00" />
                    <SPLIT distance="700" swimtime="00:14:22.42" />
                    <SPLIT distance="725" swimtime="00:14:52.82" />
                    <SPLIT distance="750" swimtime="00:15:23.78" />
                    <SPLIT distance="775" swimtime="00:15:53.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="87" swimtime="00:01:54.70" resultid="109431" heatid="110672" lane="1" entrytime="00:01:53.92">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.89" />
                    <SPLIT distance="50" swimtime="00:00:53.39" />
                    <SPLIT distance="75" swimtime="00:01:24.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="103" swimtime="00:08:18.93" resultid="109432" heatid="110842" lane="1" entrytime="00:08:13.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.42" />
                    <SPLIT distance="50" swimtime="00:00:55.83" />
                    <SPLIT distance="75" swimtime="00:01:26.23" />
                    <SPLIT distance="100" swimtime="00:01:58.42" />
                    <SPLIT distance="125" swimtime="00:02:29.96" />
                    <SPLIT distance="150" swimtime="00:03:03.28" />
                    <SPLIT distance="175" swimtime="00:03:35.67" />
                    <SPLIT distance="200" swimtime="00:04:07.85" />
                    <SPLIT distance="225" swimtime="00:04:40.16" />
                    <SPLIT distance="250" swimtime="00:05:12.48" />
                    <SPLIT distance="275" swimtime="00:05:44.58" />
                    <SPLIT distance="300" swimtime="00:06:16.37" />
                    <SPLIT distance="325" swimtime="00:06:47.39" />
                    <SPLIT distance="350" swimtime="00:07:18.48" />
                    <SPLIT distance="375" swimtime="00:07:49.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-29" firstname="Jan" gender="M" lastname="Boboli" nation="POL" athleteid="109467">
              <RESULTS>
                <RESULT eventid="98798" points="148" reactiontime="+99" swimtime="00:00:38.28" resultid="109468" heatid="110598" lane="2" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="54" reactiontime="+84" swimtime="00:00:58.68" resultid="109469" heatid="110652" lane="6" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="114" reactiontime="+90" swimtime="00:01:32.50" resultid="109470" heatid="110679" lane="6" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.57" />
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                    <SPLIT distance="75" swimtime="00:01:07.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="162" reactiontime="+87" swimtime="00:00:39.96" resultid="109471" heatid="110743" lane="8" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-13" firstname="Marcin" gender="M" lastname="Giejsztowt" nation="POL" athleteid="109384">
              <RESULTS>
                <RESULT eventid="106277" points="387" reactiontime="+73" swimtime="00:01:01.65" resultid="109385" heatid="110684" lane="7" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.18" />
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="75" swimtime="00:00:46.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="109386" heatid="110745" lane="8" entrytime="00:00:33.25" />
                <RESULT eventid="99218" points="390" reactiontime="+80" swimtime="00:02:15.93" resultid="109387" heatid="110775" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.00" />
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="75" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="125" swimtime="00:01:23.02" />
                    <SPLIT distance="150" swimtime="00:01:40.97" />
                    <SPLIT distance="175" swimtime="00:01:58.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="389" swimtime="00:04:50.60" resultid="109388" heatid="110845" lane="0" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="75" swimtime="00:00:49.59" />
                    <SPLIT distance="100" swimtime="00:01:07.18" />
                    <SPLIT distance="125" swimtime="00:01:25.02" />
                    <SPLIT distance="150" swimtime="00:01:43.28" />
                    <SPLIT distance="175" swimtime="00:02:01.87" />
                    <SPLIT distance="200" swimtime="00:02:21.09" />
                    <SPLIT distance="225" swimtime="00:02:39.69" />
                    <SPLIT distance="250" swimtime="00:02:58.88" />
                    <SPLIT distance="275" swimtime="00:03:17.91" />
                    <SPLIT distance="300" swimtime="00:03:37.58" />
                    <SPLIT distance="325" swimtime="00:03:55.93" />
                    <SPLIT distance="350" swimtime="00:04:14.73" />
                    <SPLIT distance="375" swimtime="00:04:33.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="109457">
              <RESULTS>
                <RESULT eventid="98798" status="WDR" swimtime="00:00:00.00" resultid="109458" heatid="110611" lane="1" entrytime="00:00:25.80" />
                <RESULT eventid="106277" status="WDR" swimtime="00:00:00.00" resultid="109459" heatid="110688" lane="6" entrytime="00:00:56.86" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="109461" heatid="110844" lane="7" entrytime="00:04:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="109472">
              <RESULTS>
                <RESULT eventid="98798" points="505" reactiontime="+67" swimtime="00:00:25.43" resultid="109473" heatid="110611" lane="6" entrytime="00:00:25.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="450" reactiontime="+77" swimtime="00:02:23.00" resultid="109474" heatid="110628" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                    <SPLIT distance="75" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:04.49" />
                    <SPLIT distance="125" swimtime="00:01:25.94" />
                    <SPLIT distance="150" swimtime="00:01:48.50" />
                    <SPLIT distance="175" swimtime="00:02:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="537" reactiontime="+66" swimtime="00:00:55.26" resultid="109475" heatid="110689" lane="8" entrytime="00:00:55.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.59" />
                    <SPLIT distance="50" swimtime="00:00:26.58" />
                    <SPLIT distance="75" swimtime="00:00:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="109476" heatid="110706" lane="1" entrytime="00:01:03.00" />
                <RESULT eventid="99170" points="551" reactiontime="+80" swimtime="00:00:26.59" resultid="109477" heatid="110751" lane="1" entrytime="00:00:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="WDR" swimtime="00:00:00.00" resultid="109478" heatid="110792" lane="2" entrytime="00:05:10.00" />
                <RESULT eventid="99361" points="524" reactiontime="+69" swimtime="00:01:00.05" resultid="109479" heatid="110805" lane="8" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="75" swimtime="00:00:42.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="203" reactiontime="+74" swimtime="00:02:48.92" resultid="110861" heatid="110777" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.16" />
                    <SPLIT distance="50" swimtime="00:00:25.90" />
                    <SPLIT distance="75" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:00:54.49" />
                    <SPLIT distance="125" swimtime="00:02:22.15" />
                    <SPLIT distance="150" swimtime="00:02:44.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="109462">
              <RESULTS>
                <RESULT eventid="98891" points="366" reactiontime="+72" swimtime="00:10:19.40" resultid="109463" heatid="110636" lane="4" entrytime="00:10:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.80" />
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="75" swimtime="00:00:52.19" />
                    <SPLIT distance="100" swimtime="00:01:10.83" />
                    <SPLIT distance="125" swimtime="00:01:29.68" />
                    <SPLIT distance="150" swimtime="00:01:48.81" />
                    <SPLIT distance="175" swimtime="00:02:07.72" />
                    <SPLIT distance="200" swimtime="00:02:26.98" />
                    <SPLIT distance="225" swimtime="00:02:46.37" />
                    <SPLIT distance="250" swimtime="00:03:05.52" />
                    <SPLIT distance="275" swimtime="00:03:24.86" />
                    <SPLIT distance="300" swimtime="00:03:44.41" />
                    <SPLIT distance="325" swimtime="00:04:04.09" />
                    <SPLIT distance="350" swimtime="00:04:23.79" />
                    <SPLIT distance="375" swimtime="00:04:43.46" />
                    <SPLIT distance="400" swimtime="00:05:03.28" />
                    <SPLIT distance="425" swimtime="00:05:22.61" />
                    <SPLIT distance="450" swimtime="00:05:42.52" />
                    <SPLIT distance="475" swimtime="00:06:02.21" />
                    <SPLIT distance="500" swimtime="00:06:21.95" />
                    <SPLIT distance="525" swimtime="00:06:41.60" />
                    <SPLIT distance="550" swimtime="00:07:01.57" />
                    <SPLIT distance="575" swimtime="00:07:21.34" />
                    <SPLIT distance="600" swimtime="00:07:41.30" />
                    <SPLIT distance="625" swimtime="00:08:01.50" />
                    <SPLIT distance="650" swimtime="00:08:21.94" />
                    <SPLIT distance="675" swimtime="00:08:42.25" />
                    <SPLIT distance="700" swimtime="00:09:02.41" />
                    <SPLIT distance="725" swimtime="00:09:22.28" />
                    <SPLIT distance="750" swimtime="00:09:42.33" />
                    <SPLIT distance="775" swimtime="00:10:01.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="368" reactiontime="+77" swimtime="00:01:02.68" resultid="109464" heatid="110685" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                    <SPLIT distance="75" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="405" reactiontime="+79" swimtime="00:02:14.26" resultid="109465" heatid="110775" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.15" />
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="75" swimtime="00:00:48.69" />
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                    <SPLIT distance="125" swimtime="00:01:22.92" />
                    <SPLIT distance="150" swimtime="00:01:40.44" />
                    <SPLIT distance="175" swimtime="00:01:57.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="373" swimtime="00:04:54.71" resultid="109466" heatid="110845" lane="9" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.68" />
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="75" swimtime="00:00:51.71" />
                    <SPLIT distance="100" swimtime="00:01:10.26" />
                    <SPLIT distance="125" swimtime="00:01:28.84" />
                    <SPLIT distance="150" swimtime="00:01:47.33" />
                    <SPLIT distance="175" swimtime="00:02:06.02" />
                    <SPLIT distance="200" swimtime="00:02:24.96" />
                    <SPLIT distance="225" swimtime="00:02:43.81" />
                    <SPLIT distance="250" swimtime="00:03:02.50" />
                    <SPLIT distance="275" swimtime="00:03:21.52" />
                    <SPLIT distance="300" swimtime="00:03:40.45" />
                    <SPLIT distance="325" swimtime="00:03:59.33" />
                    <SPLIT distance="350" swimtime="00:04:18.26" />
                    <SPLIT distance="375" swimtime="00:04:36.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="109406">
              <RESULTS>
                <RESULT eventid="98798" points="354" reactiontime="+88" swimtime="00:00:28.63" resultid="109407" heatid="110605" lane="3" entrytime="00:00:28.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="362" reactiontime="+93" swimtime="00:01:03.01" resultid="109408" heatid="110684" lane="1" entrytime="00:01:04.65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.58" />
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                    <SPLIT distance="75" swimtime="00:00:46.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="316" reactiontime="+93" swimtime="00:01:14.35" resultid="109409" heatid="110700" lane="3" entrytime="00:01:15.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.43" />
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="75" swimtime="00:00:57.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="290" reactiontime="+74" swimtime="00:01:13.86" resultid="109410" heatid="110761" lane="8" entrytime="00:01:15.84">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.29" />
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="75" swimtime="00:00:55.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="300" reactiontime="+81" swimtime="00:02:37.72" resultid="109411" heatid="110814" lane="2" entrytime="00:02:43.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.39" />
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="75" swimtime="00:00:56.98" />
                    <SPLIT distance="100" swimtime="00:01:17.23" />
                    <SPLIT distance="125" swimtime="00:01:36.82" />
                    <SPLIT distance="150" swimtime="00:01:57.20" />
                    <SPLIT distance="175" swimtime="00:02:17.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-17" firstname="Waldemar" gender="M" lastname="de Makay" nation="POL" athleteid="109376">
              <RESULTS>
                <RESULT eventid="98798" points="250" reactiontime="+85" swimtime="00:00:32.12" resultid="109377" heatid="110601" lane="4" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="277" reactiontime="+104" swimtime="00:21:40.38" resultid="109378" heatid="110642" lane="6" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.08" />
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="75" swimtime="00:00:58.96" />
                    <SPLIT distance="100" swimtime="00:01:20.01" />
                    <SPLIT distance="125" swimtime="00:01:40.98" />
                    <SPLIT distance="150" swimtime="00:02:02.41" />
                    <SPLIT distance="175" swimtime="00:02:23.98" />
                    <SPLIT distance="200" swimtime="00:02:45.74" />
                    <SPLIT distance="225" swimtime="00:03:07.21" />
                    <SPLIT distance="250" swimtime="00:03:28.81" />
                    <SPLIT distance="275" swimtime="00:03:50.59" />
                    <SPLIT distance="300" swimtime="00:04:12.35" />
                    <SPLIT distance="325" swimtime="00:04:34.21" />
                    <SPLIT distance="350" swimtime="00:04:55.85" />
                    <SPLIT distance="375" swimtime="00:05:17.30" />
                    <SPLIT distance="400" swimtime="00:05:39.22" />
                    <SPLIT distance="425" swimtime="00:06:00.79" />
                    <SPLIT distance="450" swimtime="00:06:22.73" />
                    <SPLIT distance="475" swimtime="00:06:44.15" />
                    <SPLIT distance="500" swimtime="00:07:06.11" />
                    <SPLIT distance="525" swimtime="00:07:28.07" />
                    <SPLIT distance="550" swimtime="00:07:49.74" />
                    <SPLIT distance="575" swimtime="00:08:11.29" />
                    <SPLIT distance="600" swimtime="00:08:33.03" />
                    <SPLIT distance="625" swimtime="00:08:54.56" />
                    <SPLIT distance="650" swimtime="00:09:16.47" />
                    <SPLIT distance="675" swimtime="00:09:38.48" />
                    <SPLIT distance="700" swimtime="00:10:00.38" />
                    <SPLIT distance="725" swimtime="00:10:21.95" />
                    <SPLIT distance="750" swimtime="00:10:43.54" />
                    <SPLIT distance="775" swimtime="00:11:05.40" />
                    <SPLIT distance="800" swimtime="00:11:27.24" />
                    <SPLIT distance="825" swimtime="00:11:49.22" />
                    <SPLIT distance="850" swimtime="00:12:11.22" />
                    <SPLIT distance="875" swimtime="00:12:33.06" />
                    <SPLIT distance="900" swimtime="00:12:54.86" />
                    <SPLIT distance="925" swimtime="00:13:16.31" />
                    <SPLIT distance="950" swimtime="00:13:38.23" />
                    <SPLIT distance="975" swimtime="00:14:00.44" />
                    <SPLIT distance="1000" swimtime="00:14:22.64" />
                    <SPLIT distance="1025" swimtime="00:14:44.66" />
                    <SPLIT distance="1050" swimtime="00:15:06.58" />
                    <SPLIT distance="1075" swimtime="00:15:28.63" />
                    <SPLIT distance="1100" swimtime="00:15:50.39" />
                    <SPLIT distance="1125" swimtime="00:16:12.55" />
                    <SPLIT distance="1150" swimtime="00:16:34.42" />
                    <SPLIT distance="1175" swimtime="00:16:56.72" />
                    <SPLIT distance="1200" swimtime="00:17:18.62" />
                    <SPLIT distance="1225" swimtime="00:17:40.60" />
                    <SPLIT distance="1250" swimtime="00:18:02.51" />
                    <SPLIT distance="1275" swimtime="00:18:24.41" />
                    <SPLIT distance="1300" swimtime="00:18:46.23" />
                    <SPLIT distance="1325" swimtime="00:19:07.79" />
                    <SPLIT distance="1350" swimtime="00:19:29.91" />
                    <SPLIT distance="1375" swimtime="00:19:52.01" />
                    <SPLIT distance="1400" swimtime="00:20:14.07" />
                    <SPLIT distance="1425" swimtime="00:20:36.19" />
                    <SPLIT distance="1450" swimtime="00:20:58.17" />
                    <SPLIT distance="1475" swimtime="00:21:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="162" reactiontime="+92" swimtime="00:00:40.70" resultid="109379" heatid="110654" lane="2" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="237" swimtime="00:01:12.59" resultid="109380" heatid="110682" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="75" swimtime="00:00:53.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="163" reactiontime="+84" swimtime="00:01:29.43" resultid="109381" heatid="110759" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.72" />
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                    <SPLIT distance="75" swimtime="00:01:06.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="255" reactiontime="+103" swimtime="00:02:36.58" resultid="109382" heatid="110773" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.72" />
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="75" swimtime="00:00:56.07" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="125" swimtime="00:01:35.75" />
                    <SPLIT distance="150" swimtime="00:01:56.39" />
                    <SPLIT distance="175" swimtime="00:02:17.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="273" reactiontime="+106" swimtime="00:05:27.13" resultid="109383" heatid="110847" lane="8" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.86" />
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                    <SPLIT distance="75" swimtime="00:00:56.76" />
                    <SPLIT distance="100" swimtime="00:01:17.10" />
                    <SPLIT distance="125" swimtime="00:01:37.76" />
                    <SPLIT distance="150" swimtime="00:01:58.71" />
                    <SPLIT distance="175" swimtime="00:02:19.46" />
                    <SPLIT distance="200" swimtime="00:02:40.34" />
                    <SPLIT distance="225" swimtime="00:03:00.93" />
                    <SPLIT distance="250" swimtime="00:03:22.11" />
                    <SPLIT distance="275" swimtime="00:03:43.21" />
                    <SPLIT distance="300" swimtime="00:04:04.31" />
                    <SPLIT distance="325" swimtime="00:04:25.65" />
                    <SPLIT distance="350" swimtime="00:04:46.81" />
                    <SPLIT distance="375" swimtime="00:05:07.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="330" reactiontime="+113" swimtime="00:01:59.51" resultid="109480" heatid="110783" lane="1" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.07" />
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                    <SPLIT distance="75" swimtime="00:00:46.35" />
                    <SPLIT distance="100" swimtime="00:01:02.80" />
                    <SPLIT distance="125" swimtime="00:01:16.88" />
                    <SPLIT distance="150" swimtime="00:01:32.36" />
                    <SPLIT distance="175" swimtime="00:01:45.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109370" number="1" reactiontime="+113" />
                    <RELAYPOSITION athleteid="109376" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="109406" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="109397" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="253" reactiontime="+88" swimtime="00:02:22.99" resultid="109481" heatid="110717" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.77" />
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="75" swimtime="00:00:55.04" />
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="125" swimtime="00:01:33.08" />
                    <SPLIT distance="150" swimtime="00:01:51.23" />
                    <SPLIT distance="175" swimtime="00:02:06.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109370" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="109433" number="2" />
                    <RELAYPOSITION athleteid="109406" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="109376" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="99059" points="390" reactiontime="+84" swimtime="00:02:03.83" resultid="109482" heatid="110719" lane="9" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.88" />
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="75" swimtime="00:00:47.57" />
                    <SPLIT distance="100" swimtime="00:01:05.50" />
                    <SPLIT distance="125" swimtime="00:01:19.29" />
                    <SPLIT distance="150" swimtime="00:01:36.46" />
                    <SPLIT distance="175" swimtime="00:01:49.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109397" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="109462" number="2" />
                    <RELAYPOSITION athleteid="109439" number="3" />
                    <RELAYPOSITION athleteid="109457" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="99250" points="413" reactiontime="+79" swimtime="00:01:50.86" resultid="109483" heatid="110784" lane="8" entrytime="00:01:47.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.22" />
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="75" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:00:56.29" />
                    <SPLIT distance="125" swimtime="00:01:09.76" />
                    <SPLIT distance="150" swimtime="00:01:24.77" />
                    <SPLIT distance="175" swimtime="00:01:37.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109352" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="109462" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="109439" number="3" reactiontime="+2" />
                    <RELAYPOSITION athleteid="109457" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="106680" name="Weteran Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" phone="604 522 654" street="ŚW.JANA  4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="502611100009" athleteid="106708">
              <RESULTS>
                <RESULT eventid="98863" points="471" reactiontime="+82" swimtime="00:10:15.75" resultid="106709" heatid="110633" lane="4" entrytime="00:10:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.56" />
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="75" swimtime="00:00:53.07" />
                    <SPLIT distance="100" swimtime="00:01:11.64" />
                    <SPLIT distance="125" swimtime="00:01:30.40" />
                    <SPLIT distance="150" swimtime="00:01:49.23" />
                    <SPLIT distance="175" swimtime="00:02:08.29" />
                    <SPLIT distance="200" swimtime="00:02:27.37" />
                    <SPLIT distance="225" swimtime="00:02:46.56" />
                    <SPLIT distance="250" swimtime="00:03:05.59" />
                    <SPLIT distance="275" swimtime="00:03:24.97" />
                    <SPLIT distance="300" swimtime="00:03:44.16" />
                    <SPLIT distance="325" swimtime="00:04:03.65" />
                    <SPLIT distance="350" swimtime="00:04:23.05" />
                    <SPLIT distance="375" swimtime="00:04:42.61" />
                    <SPLIT distance="400" swimtime="00:05:02.07" />
                    <SPLIT distance="425" swimtime="00:05:21.80" />
                    <SPLIT distance="450" swimtime="00:05:41.21" />
                    <SPLIT distance="475" swimtime="00:06:01.06" />
                    <SPLIT distance="500" swimtime="00:06:20.59" />
                    <SPLIT distance="525" swimtime="00:06:40.59" />
                    <SPLIT distance="550" swimtime="00:07:00.28" />
                    <SPLIT distance="575" swimtime="00:07:20.10" />
                    <SPLIT distance="600" swimtime="00:07:39.67" />
                    <SPLIT distance="625" swimtime="00:07:59.66" />
                    <SPLIT distance="650" swimtime="00:08:19.35" />
                    <SPLIT distance="675" swimtime="00:08:38.96" />
                    <SPLIT distance="700" swimtime="00:08:58.59" />
                    <SPLIT distance="725" swimtime="00:09:18.65" />
                    <SPLIT distance="750" swimtime="00:09:38.30" />
                    <SPLIT distance="775" swimtime="00:09:57.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="437" reactiontime="+74" swimtime="00:02:57.30" resultid="106710" heatid="110664" lane="2" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.50" />
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                    <SPLIT distance="75" swimtime="00:01:01.61" />
                    <SPLIT distance="100" swimtime="00:01:23.91" />
                    <SPLIT distance="125" swimtime="00:01:46.80" />
                    <SPLIT distance="150" swimtime="00:02:10.24" />
                    <SPLIT distance="175" swimtime="00:02:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="450" reactiontime="+88" swimtime="00:01:21.37" resultid="106711" heatid="110725" lane="1" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.01" />
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="75" swimtime="00:00:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="451" swimtime="00:02:24.41" resultid="106712" heatid="110768" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.16" />
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="75" swimtime="00:00:51.50" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="125" swimtime="00:01:28.54" />
                    <SPLIT distance="150" swimtime="00:01:47.48" />
                    <SPLIT distance="175" swimtime="00:02:06.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="418" swimtime="00:00:38.49" resultid="106713" heatid="110822" lane="5" entrytime="00:00:38.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="469" swimtime="00:05:01.83" resultid="106714" heatid="110839" lane="6" entrytime="00:05:01.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.31" />
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="75" swimtime="00:00:52.50" />
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="125" swimtime="00:01:29.59" />
                    <SPLIT distance="150" swimtime="00:01:48.56" />
                    <SPLIT distance="175" swimtime="00:02:07.78" />
                    <SPLIT distance="200" swimtime="00:02:27.00" />
                    <SPLIT distance="225" swimtime="00:02:46.20" />
                    <SPLIT distance="250" swimtime="00:03:05.72" />
                    <SPLIT distance="275" swimtime="00:03:25.11" />
                    <SPLIT distance="300" swimtime="00:03:44.65" />
                    <SPLIT distance="325" swimtime="00:04:04.10" />
                    <SPLIT distance="350" swimtime="00:04:23.87" />
                    <SPLIT distance="375" swimtime="00:04:43.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-07-16" firstname="Ewald" gender="M" lastname="Bastek" nation="POL" license="502611200001" athleteid="106686">
              <RESULTS>
                <RESULT eventid="98798" points="158" reactiontime="+103" swimtime="00:00:37.43" resultid="106687" heatid="110598" lane="0" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="146" reactiontime="+112" swimtime="00:01:25.25" resultid="106688" heatid="110680" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.33" />
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                    <SPLIT distance="75" swimtime="00:01:02.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="137" reactiontime="+96" swimtime="00:03:12.42" resultid="106689" heatid="110770" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.17" />
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                    <SPLIT distance="75" swimtime="00:01:09.59" />
                    <SPLIT distance="100" swimtime="00:01:34.83" />
                    <SPLIT distance="125" swimtime="00:02:00.16" />
                    <SPLIT distance="150" swimtime="00:02:24.68" />
                    <SPLIT distance="175" swimtime="00:02:49.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="74" swimtime="00:01:54.99" resultid="106690" heatid="110798" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.15" />
                    <SPLIT distance="50" swimtime="00:00:55.83" />
                    <SPLIT distance="75" swimtime="00:01:25.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-05" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" license="502611100005" athleteid="106719">
              <RESULTS>
                <RESULT eventid="98777" points="181" reactiontime="+97" swimtime="00:00:41.06" resultid="106720" heatid="110587" lane="7" entrytime="00:00:42.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" license="502611200004" athleteid="106721">
              <RESULTS>
                <RESULT eventid="98924" points="142" reactiontime="+59" swimtime="00:00:42.54" resultid="106722" heatid="110653" lane="3" entrytime="00:00:42.59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="125" reactiontime="+76" swimtime="00:01:37.75" resultid="106723" heatid="110758" lane="4" entrytime="00:01:37.37">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.70" />
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                    <SPLIT distance="75" swimtime="00:01:12.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="107" reactiontime="+72" swimtime="00:03:42.20" resultid="106724" heatid="110812" lane="9" entrytime="00:03:36.72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.21" />
                    <SPLIT distance="50" swimtime="00:00:49.68" />
                    <SPLIT distance="75" swimtime="00:01:19.20" />
                    <SPLIT distance="100" swimtime="00:01:46.27" />
                    <SPLIT distance="125" swimtime="00:02:14.99" />
                    <SPLIT distance="150" swimtime="00:02:43.94" />
                    <SPLIT distance="175" swimtime="00:03:13.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="502611200005" athleteid="106715">
              <RESULTS>
                <RESULT eventid="98798" points="134" reactiontime="+107" swimtime="00:00:39.54" resultid="106716" heatid="110598" lane="1" entrytime="00:00:38.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="74" reactiontime="+95" swimtime="00:00:52.70" resultid="106717" heatid="110652" lane="3" entrytime="00:00:51.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="86" swimtime="00:00:49.23" resultid="106718" heatid="110742" lane="5" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-28" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="502611200007" athleteid="106704">
              <RESULTS>
                <RESULT eventid="98798" points="251" reactiontime="+84" swimtime="00:00:32.10" resultid="106705" heatid="110601" lane="5" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="165" reactiontime="+86" swimtime="00:01:32.33" resultid="106706" heatid="110697" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.48" />
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="75" swimtime="00:01:12.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="228" reactiontime="+94" swimtime="00:00:35.64" resultid="106707" heatid="110743" lane="5" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-14" firstname="Maciej" gender="M" lastname="Kunicki" nation="POL" license="502611200011" athleteid="106699">
              <RESULTS>
                <RESULT eventid="98830" points="276" reactiontime="+87" swimtime="00:02:48.18" resultid="106700" heatid="110623" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.10" />
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="75" swimtime="00:00:56.38" />
                    <SPLIT distance="100" swimtime="00:01:18.56" />
                    <SPLIT distance="125" swimtime="00:01:45.02" />
                    <SPLIT distance="150" swimtime="00:02:10.70" />
                    <SPLIT distance="175" swimtime="00:02:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="239" reactiontime="+87" swimtime="00:02:54.80" resultid="106701" heatid="110712" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.07" />
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                    <SPLIT distance="75" swimtime="00:01:00.44" />
                    <SPLIT distance="100" swimtime="00:01:23.20" />
                    <SPLIT distance="125" swimtime="00:01:45.97" />
                    <SPLIT distance="150" swimtime="00:02:09.73" />
                    <SPLIT distance="175" swimtime="00:02:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="316" swimtime="00:00:31.98" resultid="106702" heatid="110746" lane="9" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="262" reactiontime="+91" swimtime="00:01:15.67" resultid="106703" heatid="110801" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.07" />
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="75" swimtime="00:00:56.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="502611100001" athleteid="106691">
              <RESULTS>
                <RESULT eventid="98777" points="237" reactiontime="+85" swimtime="00:00:37.54" resultid="106692" heatid="110588" lane="6" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106294" points="159" reactiontime="+71" swimtime="00:00:47.34" resultid="106693" heatid="110648" lane="9" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="200" swimtime="00:01:27.05" resultid="106694" heatid="110673" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.77" />
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                    <SPLIT distance="75" swimtime="00:01:05.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="116" reactiontime="+81" swimtime="00:00:49.95" resultid="106695" heatid="110736" lane="5" entrytime="00:00:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-22" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" license="502611100004" athleteid="106696">
              <RESULTS>
                <RESULT eventid="106294" points="95" reactiontime="+96" swimtime="00:00:56.25" resultid="106697" heatid="110646" lane="1" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="160" swimtime="00:00:53.03" resultid="106698" heatid="110818" lane="6" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="146" reactiontime="+82" swimtime="00:02:51.64" resultid="106726" heatid="110717" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.69" />
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                    <SPLIT distance="75" swimtime="00:01:08.59" />
                    <SPLIT distance="100" swimtime="00:01:35.01" />
                    <SPLIT distance="125" swimtime="00:01:51.85" />
                    <SPLIT distance="150" swimtime="00:02:12.70" />
                    <SPLIT distance="175" swimtime="00:02:31.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106721" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="106686" number="2" />
                    <RELAYPOSITION athleteid="106704" number="3" />
                    <RELAYPOSITION athleteid="106715" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="99250" points="162" swimtime="00:02:31.23" resultid="106727" heatid="110782" lane="9" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.90" />
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                    <SPLIT distance="75" swimtime="00:00:55.94" />
                    <SPLIT distance="100" swimtime="00:01:16.76" />
                    <SPLIT distance="125" swimtime="00:01:35.18" />
                    <SPLIT distance="150" swimtime="00:01:55.90" />
                    <SPLIT distance="175" swimtime="00:02:12.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106686" number="1" />
                    <RELAYPOSITION athleteid="106721" number="2" />
                    <RELAYPOSITION athleteid="106715" number="3" />
                    <RELAYPOSITION athleteid="106704" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="99036" points="215" reactiontime="+73" swimtime="00:02:53.65" resultid="106729" heatid="110715" lane="0" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.37" />
                    <SPLIT distance="50" swimtime="00:00:45.16" />
                    <SPLIT distance="75" swimtime="00:01:09.39" />
                    <SPLIT distance="100" swimtime="00:01:38.67" />
                    <SPLIT distance="125" swimtime="00:01:54.43" />
                    <SPLIT distance="150" swimtime="00:02:12.99" />
                    <SPLIT distance="175" swimtime="00:02:31.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106691" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="106696" number="2" />
                    <RELAYPOSITION athleteid="106708" number="3" />
                    <RELAYPOSITION athleteid="106719" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="99441" points="143" reactiontime="+74" swimtime="00:02:52.92" resultid="106728" heatid="110836" lane="8" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.46" />
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                    <SPLIT distance="75" swimtime="00:01:10.03" />
                    <SPLIT distance="100" swimtime="00:01:39.29" />
                    <SPLIT distance="125" swimtime="00:01:55.57" />
                    <SPLIT distance="150" swimtime="00:02:15.35" />
                    <SPLIT distance="175" swimtime="00:02:33.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106691" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="106696" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="106704" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="106686" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="98846" points="162" reactiontime="+79" swimtime="00:02:31.44" resultid="106725" heatid="110629" lane="4" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.17" />
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="75" swimtime="00:00:56.75" />
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="125" swimtime="00:01:35.52" />
                    <SPLIT distance="150" swimtime="00:01:56.83" />
                    <SPLIT distance="175" swimtime="00:02:13.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106691" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="106686" number="2" reactiontime="+71" />
                    <RELAYPOSITION athleteid="106719" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="106704" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WKS" nation="POL" region="DOL" clubid="107733" name="WKS Śląsk Wrocław">
          <CONTACT email="marrot68@wp.pl" name="Rother Marek" />
          <ATHLETES>
            <ATHLETE birthdate="1968-05-21" firstname="Marek" gender="M" lastname="Rother" nation="POL" athleteid="107734">
              <RESULTS>
                <RESULT eventid="98830" points="406" reactiontime="+87" swimtime="00:02:28.00" resultid="107735" heatid="110626" lane="0" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.24" />
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="75" swimtime="00:00:50.61" />
                    <SPLIT distance="100" swimtime="00:01:08.65" />
                    <SPLIT distance="125" swimtime="00:01:30.39" />
                    <SPLIT distance="150" swimtime="00:01:53.05" />
                    <SPLIT distance="175" swimtime="00:02:11.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="423" reactiontime="+60" swimtime="00:00:29.58" resultid="107736" heatid="110660" lane="9" entrytime="00:00:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="425" reactiontime="+73" swimtime="00:01:07.38" resultid="107737" heatid="110704" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="75" swimtime="00:00:50.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="441" reactiontime="+73" swimtime="00:01:04.24" resultid="107738" heatid="110763" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.22" />
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="75" swimtime="00:00:47.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="408" reactiontime="+64" swimtime="00:02:22.39" resultid="107739" heatid="110816" lane="8" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.63" />
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="75" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:08.47" />
                    <SPLIT distance="125" swimtime="00:01:26.74" />
                    <SPLIT distance="150" swimtime="00:01:45.08" />
                    <SPLIT distance="175" swimtime="00:02:03.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="108942" name="Wyższa Szkoła Biznesu w Dąbrowie Górniczej" shortname="WS Biznesu w Dąbrowie Gr.">
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" swrid="4086800" athleteid="108943">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="108945" heatid="110610" lane="2" entrytime="00:00:26.00" entrycourse="SCM" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="108946" heatid="110623" lane="9" entrytime="00:03:00.00" entrycourse="SCM" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="108947" heatid="110658" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="98956" points="302" swimtime="00:02:59.41" resultid="108948" heatid="110668" lane="6" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.28" />
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="75" swimtime="00:00:58.66" />
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                    <SPLIT distance="125" swimtime="00:01:44.22" />
                    <SPLIT distance="150" swimtime="00:02:08.23" />
                    <SPLIT distance="175" swimtime="00:02:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="368" reactiontime="+77" swimtime="00:01:17.60" resultid="108949" heatid="110734" lane="1" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.54" />
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="75" swimtime="00:00:55.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="262" reactiontime="+70" swimtime="00:01:16.43" resultid="108951" heatid="110760" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.36" />
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="75" swimtime="00:00:56.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="218" reactiontime="+65" swimtime="00:02:55.30" resultid="108952" heatid="110813" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.63" />
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="75" swimtime="00:01:02.56" />
                    <SPLIT distance="100" swimtime="00:01:25.24" />
                    <SPLIT distance="125" swimtime="00:01:47.90" />
                    <SPLIT distance="150" swimtime="00:02:10.79" />
                    <SPLIT distance="175" swimtime="00:02:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="432" reactiontime="+58" swimtime="00:00:33.38" resultid="108953" heatid="110833" lane="5" entrytime="00:00:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="108941" name="Wyższa Szkoła Humanitas w Sosnowcu" shortname="WS Humanitas w Sosnowcu">
          <ATHLETES>
            <ATHLETE birthdate="1996-03-24" firstname="KINGA" gender="F" lastname="PLUTA" nation="POL" athleteid="108944">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="108954" heatid="110591" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="108955" heatid="110616" lane="6" entrytime="00:03:10.00" />
                <RESULT eventid="98940" points="391" reactiontime="+88" swimtime="00:03:03.97" resultid="108956" heatid="110664" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.09" />
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="75" swimtime="00:01:03.41" />
                    <SPLIT distance="100" swimtime="00:01:26.27" />
                    <SPLIT distance="125" swimtime="00:01:50.14" />
                    <SPLIT distance="150" swimtime="00:02:14.65" />
                    <SPLIT distance="175" swimtime="00:02:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="108957" heatid="110694" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="99089" points="432" reactiontime="+83" swimtime="00:01:22.48" resultid="108958" heatid="110724" lane="4" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.09" />
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="75" swimtime="00:01:00.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="388" swimtime="00:02:31.78" resultid="108959" heatid="110767" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.77" />
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="75" swimtime="00:00:52.27" />
                    <SPLIT distance="100" swimtime="00:01:11.41" />
                    <SPLIT distance="125" swimtime="00:01:31.18" />
                    <SPLIT distance="150" swimtime="00:01:51.64" />
                    <SPLIT distance="175" swimtime="00:02:12.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="295" reactiontime="+83" swimtime="00:02:58.98" resultid="108960" heatid="110808" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.49" />
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                    <SPLIT distance="75" swimtime="00:01:05.54" />
                    <SPLIT distance="100" swimtime="00:01:28.31" />
                    <SPLIT distance="125" swimtime="00:01:51.55" />
                    <SPLIT distance="150" swimtime="00:02:14.69" />
                    <SPLIT distance="175" swimtime="00:02:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="468" reactiontime="+85" swimtime="00:00:37.09" resultid="108961" heatid="110823" lane="3" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="106326" name="Zawodnik Niezrzeszony">
          <CONTACT city="KRAKÓW" email="piotr_urbanczyk@onet.pl" name="URBAŃCZYK" phone="608172201" />
          <ATHLETES>
            <ATHLETE birthdate="1986-08-06" firstname="Oleksandr" gender="M" lastname="Broshevan" nation="POL" athleteid="110418">
              <RESULTS>
                <RESULT eventid="98798" points="385" reactiontime="+94" swimtime="00:00:27.84" resultid="110419" heatid="110595" lane="3" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="276" reactiontime="+104" swimtime="00:02:48.33" resultid="110420" heatid="110626" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.46" />
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="75" swimtime="00:00:56.21" />
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                    <SPLIT distance="125" swimtime="00:01:43.77" />
                    <SPLIT distance="150" swimtime="00:02:09.47" />
                    <SPLIT distance="175" swimtime="00:02:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="295" reactiontime="+101" swimtime="00:00:33.35" resultid="110421" heatid="110658" lane="0" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="328" reactiontime="+102" swimtime="00:01:05.10" resultid="110422" heatid="110687" lane="5" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.43" />
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                    <SPLIT distance="75" swimtime="00:00:47.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="231" reactiontime="+97" swimtime="00:02:51.92" resultid="110423" heatid="110811" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.30" />
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="75" swimtime="00:01:00.98" />
                    <SPLIT distance="100" swimtime="00:01:23.62" />
                    <SPLIT distance="125" swimtime="00:01:47.09" />
                    <SPLIT distance="150" swimtime="00:02:11.14" />
                    <SPLIT distance="175" swimtime="00:02:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="325" swimtime="00:00:36.72" resultid="110424" heatid="110830" lane="9" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="110858" heatid="110726" lane="6" late="yes" />
                <RESULT eventid="99186" points="255" reactiontime="+101" swimtime="00:01:17.05" resultid="110859" heatid="110757" lane="0" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.59" />
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="75" swimtime="00:00:57.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="385" reactiontime="+92" swimtime="00:00:29.96" resultid="110863" heatid="110741" lane="7" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-11-22" firstname="Marek" gender="M" lastname="Pałysa" nation="POL" athleteid="110495">
              <RESULTS>
                <RESULT eventid="98891" points="253" reactiontime="+94" swimtime="00:11:40.79" resultid="110496" heatid="110637" lane="5" entrytime="00:11:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.56" />
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                    <SPLIT distance="75" swimtime="00:00:58.28" />
                    <SPLIT distance="100" swimtime="00:01:19.14" />
                    <SPLIT distance="125" swimtime="00:01:40.61" />
                    <SPLIT distance="150" swimtime="00:02:02.72" />
                    <SPLIT distance="175" swimtime="00:02:25.46" />
                    <SPLIT distance="200" swimtime="00:02:47.70" />
                    <SPLIT distance="225" swimtime="00:03:10.14" />
                    <SPLIT distance="250" swimtime="00:03:32.68" />
                    <SPLIT distance="275" swimtime="00:03:54.77" />
                    <SPLIT distance="300" swimtime="00:04:17.13" />
                    <SPLIT distance="325" swimtime="00:04:39.03" />
                    <SPLIT distance="350" swimtime="00:05:01.30" />
                    <SPLIT distance="375" swimtime="00:05:23.29" />
                    <SPLIT distance="400" swimtime="00:05:45.68" />
                    <SPLIT distance="425" swimtime="00:06:07.91" />
                    <SPLIT distance="450" swimtime="00:06:30.64" />
                    <SPLIT distance="475" swimtime="00:06:52.63" />
                    <SPLIT distance="500" swimtime="00:07:15.58" />
                    <SPLIT distance="525" swimtime="00:07:38.10" />
                    <SPLIT distance="550" swimtime="00:08:00.73" />
                    <SPLIT distance="575" swimtime="00:08:22.98" />
                    <SPLIT distance="600" swimtime="00:08:45.73" />
                    <SPLIT distance="625" swimtime="00:09:08.03" />
                    <SPLIT distance="650" swimtime="00:09:30.49" />
                    <SPLIT distance="675" swimtime="00:09:52.68" />
                    <SPLIT distance="700" swimtime="00:10:15.05" />
                    <SPLIT distance="725" swimtime="00:10:37.15" />
                    <SPLIT distance="750" swimtime="00:10:59.53" />
                    <SPLIT distance="775" swimtime="00:11:21.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="257" reactiontime="+88" swimtime="00:05:33.45" resultid="110497" heatid="110847" lane="4" entrytime="00:05:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.91" />
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="75" swimtime="00:00:52.51" />
                    <SPLIT distance="100" swimtime="00:01:11.94" />
                    <SPLIT distance="125" swimtime="00:01:32.01" />
                    <SPLIT distance="150" swimtime="00:01:52.47" />
                    <SPLIT distance="175" swimtime="00:02:13.88" />
                    <SPLIT distance="200" swimtime="00:02:35.81" />
                    <SPLIT distance="225" swimtime="00:02:57.81" />
                    <SPLIT distance="250" swimtime="00:03:19.93" />
                    <SPLIT distance="275" swimtime="00:03:42.84" />
                    <SPLIT distance="300" swimtime="00:04:04.62" />
                    <SPLIT distance="325" swimtime="00:04:27.49" />
                    <SPLIT distance="350" swimtime="00:04:50.55" />
                    <SPLIT distance="375" swimtime="00:05:13.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Bartłomiej" gender="M" lastname="Kurek" nation="POL" swrid="4104735" athleteid="110414">
              <RESULTS>
                <RESULT eventid="98924" points="400" reactiontime="+74" swimtime="00:00:30.14" resultid="110415" heatid="110659" lane="5" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="402" reactiontime="+73" swimtime="00:01:08.59" resultid="110416" heatid="110705" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="75" swimtime="00:00:52.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="497" reactiontime="+69" swimtime="00:00:27.52" resultid="110417" heatid="110749" lane="4" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-07" firstname="Marcin" gender="M" lastname="Musialik" nation="POL" swrid="4509577" athleteid="110430">
              <RESULTS>
                <RESULT eventid="98830" points="421" reactiontime="+89" swimtime="00:02:26.17" resultid="110431" heatid="110626" lane="5" entrytime="00:02:30.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="75" swimtime="00:00:50.26" />
                    <SPLIT distance="100" swimtime="00:01:08.51" />
                    <SPLIT distance="125" swimtime="00:01:30.37" />
                    <SPLIT distance="150" swimtime="00:01:52.38" />
                    <SPLIT distance="175" swimtime="00:02:09.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="472" reactiontime="+87" swimtime="00:18:08.63" resultid="110432" heatid="110641" lane="6" entrytime="00:19:00.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.43" />
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="75" swimtime="00:00:50.24" />
                    <SPLIT distance="100" swimtime="00:01:08.13" />
                    <SPLIT distance="125" swimtime="00:01:25.86" />
                    <SPLIT distance="150" swimtime="00:01:44.16" />
                    <SPLIT distance="175" swimtime="00:02:02.01" />
                    <SPLIT distance="200" swimtime="00:02:20.51" />
                    <SPLIT distance="225" swimtime="00:02:38.81" />
                    <SPLIT distance="250" swimtime="00:02:57.43" />
                    <SPLIT distance="275" swimtime="00:03:15.90" />
                    <SPLIT distance="300" swimtime="00:03:34.59" />
                    <SPLIT distance="325" swimtime="00:03:52.96" />
                    <SPLIT distance="350" swimtime="00:04:11.56" />
                    <SPLIT distance="375" swimtime="00:04:29.80" />
                    <SPLIT distance="400" swimtime="00:04:48.56" />
                    <SPLIT distance="425" swimtime="00:05:06.80" />
                    <SPLIT distance="450" swimtime="00:05:25.53" />
                    <SPLIT distance="475" swimtime="00:05:43.80" />
                    <SPLIT distance="500" swimtime="00:06:02.08" />
                    <SPLIT distance="525" swimtime="00:06:20.35" />
                    <SPLIT distance="550" swimtime="00:06:38.61" />
                    <SPLIT distance="575" swimtime="00:06:56.71" />
                    <SPLIT distance="600" swimtime="00:07:15.10" />
                    <SPLIT distance="625" swimtime="00:07:33.29" />
                    <SPLIT distance="650" swimtime="00:07:51.81" />
                    <SPLIT distance="675" swimtime="00:08:09.93" />
                    <SPLIT distance="700" swimtime="00:08:28.30" />
                    <SPLIT distance="725" swimtime="00:08:46.30" />
                    <SPLIT distance="750" swimtime="00:09:04.71" />
                    <SPLIT distance="775" swimtime="00:09:23.08" />
                    <SPLIT distance="800" swimtime="00:09:41.58" />
                    <SPLIT distance="825" swimtime="00:09:59.83" />
                    <SPLIT distance="850" swimtime="00:10:18.40" />
                    <SPLIT distance="875" swimtime="00:10:36.64" />
                    <SPLIT distance="900" swimtime="00:10:55.23" />
                    <SPLIT distance="925" swimtime="00:11:13.55" />
                    <SPLIT distance="950" swimtime="00:11:32.12" />
                    <SPLIT distance="975" swimtime="00:11:50.36" />
                    <SPLIT distance="1000" swimtime="00:12:08.99" />
                    <SPLIT distance="1025" swimtime="00:12:27.26" />
                    <SPLIT distance="1050" swimtime="00:12:45.91" />
                    <SPLIT distance="1075" swimtime="00:13:04.25" />
                    <SPLIT distance="1100" swimtime="00:13:23.19" />
                    <SPLIT distance="1125" swimtime="00:13:41.28" />
                    <SPLIT distance="1150" swimtime="00:13:59.59" />
                    <SPLIT distance="1175" swimtime="00:14:17.11" />
                    <SPLIT distance="1200" swimtime="00:14:35.33" />
                    <SPLIT distance="1225" swimtime="00:14:53.41" />
                    <SPLIT distance="1250" swimtime="00:15:11.97" />
                    <SPLIT distance="1275" swimtime="00:15:30.24" />
                    <SPLIT distance="1300" swimtime="00:15:48.47" />
                    <SPLIT distance="1325" swimtime="00:16:05.59" />
                    <SPLIT distance="1350" swimtime="00:16:23.16" />
                    <SPLIT distance="1375" swimtime="00:16:40.41" />
                    <SPLIT distance="1400" swimtime="00:16:58.26" />
                    <SPLIT distance="1425" swimtime="00:17:15.61" />
                    <SPLIT distance="1450" swimtime="00:17:33.44" />
                    <SPLIT distance="1475" swimtime="00:17:51.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="304" reactiontime="+66" swimtime="00:00:33.04" resultid="110433" heatid="110656" lane="5" entrytime="00:00:34.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="357" reactiontime="+87" swimtime="00:02:32.94" resultid="110434" heatid="110713" lane="1" entrytime="00:02:35.84">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.31" />
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="75" swimtime="00:00:54.14" />
                    <SPLIT distance="100" swimtime="00:01:14.08" />
                    <SPLIT distance="125" swimtime="00:01:33.89" />
                    <SPLIT distance="150" swimtime="00:01:53.84" />
                    <SPLIT distance="175" swimtime="00:02:13.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="349" reactiontime="+66" swimtime="00:01:09.43" resultid="110435" heatid="110762" lane="9" entrytime="00:01:12.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.59" />
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="75" swimtime="00:00:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="432" reactiontime="+98" swimtime="00:05:11.49" resultid="110436" heatid="110792" lane="1" entrytime="00:05:23.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.63" />
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="75" swimtime="00:00:51.48" />
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                    <SPLIT distance="125" swimtime="00:01:30.83" />
                    <SPLIT distance="150" swimtime="00:01:50.35" />
                    <SPLIT distance="175" swimtime="00:02:09.86" />
                    <SPLIT distance="200" swimtime="00:02:29.53" />
                    <SPLIT distance="225" swimtime="00:02:52.10" />
                    <SPLIT distance="250" swimtime="00:03:14.34" />
                    <SPLIT distance="275" swimtime="00:03:37.09" />
                    <SPLIT distance="300" swimtime="00:04:00.38" />
                    <SPLIT distance="325" swimtime="00:04:18.50" />
                    <SPLIT distance="350" swimtime="00:04:36.19" />
                    <SPLIT distance="375" swimtime="00:04:54.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="374" reactiontime="+71" swimtime="00:02:26.48" resultid="110437" heatid="110815" lane="4" entrytime="00:02:28.43">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="75" swimtime="00:00:53.78" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="125" swimtime="00:01:31.31" />
                    <SPLIT distance="150" swimtime="00:01:49.79" />
                    <SPLIT distance="175" swimtime="00:02:08.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="473" reactiontime="+85" swimtime="00:04:32.41" resultid="110438" heatid="110843" lane="8" entrytime="00:04:38.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.45" />
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="75" swimtime="00:00:47.73" />
                    <SPLIT distance="100" swimtime="00:01:04.69" />
                    <SPLIT distance="125" swimtime="00:01:21.55" />
                    <SPLIT distance="150" swimtime="00:01:38.65" />
                    <SPLIT distance="175" swimtime="00:01:55.95" />
                    <SPLIT distance="200" swimtime="00:02:13.47" />
                    <SPLIT distance="225" swimtime="00:02:30.95" />
                    <SPLIT distance="250" swimtime="00:02:48.29" />
                    <SPLIT distance="275" swimtime="00:03:05.76" />
                    <SPLIT distance="300" swimtime="00:03:23.12" />
                    <SPLIT distance="325" swimtime="00:03:40.60" />
                    <SPLIT distance="350" swimtime="00:03:58.20" />
                    <SPLIT distance="375" swimtime="00:04:15.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Mateusz" gender="M" lastname="Jaskier" nation="POL" swrid="4363436" athleteid="110529">
              <RESULTS>
                <RESULT eventid="98798" points="517" reactiontime="+73" swimtime="00:00:25.24" resultid="110530" heatid="110611" lane="7" entrytime="00:00:25.68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="433" reactiontime="+84" swimtime="00:02:24.80" resultid="110531" heatid="110627" lane="4" entrytime="00:02:25.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="75" swimtime="00:00:50.26" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="125" swimtime="00:01:29.74" />
                    <SPLIT distance="150" swimtime="00:01:50.26" />
                    <SPLIT distance="175" swimtime="00:02:08.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="480" reactiontime="+77" swimtime="00:02:33.82" resultid="110532" heatid="110670" lane="3" entrytime="00:02:31.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.97" />
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="75" swimtime="00:00:51.38" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="125" swimtime="00:01:31.05" />
                    <SPLIT distance="150" swimtime="00:01:51.67" />
                    <SPLIT distance="175" swimtime="00:02:12.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="535" swimtime="00:01:02.38" resultid="110533" heatid="110705" lane="6" entrytime="00:01:05.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.63" />
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                    <SPLIT distance="75" swimtime="00:00:47.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="569" swimtime="00:01:07.07" resultid="110534" heatid="110734" lane="6" entrytime="00:01:07.19">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.33" />
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="75" swimtime="00:00:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="524" reactiontime="+64" swimtime="00:00:27.04" resultid="110535" heatid="110750" lane="7" entrytime="00:00:27.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="473" reactiontime="+78" swimtime="00:01:02.16" resultid="110536" heatid="110804" lane="1" entrytime="00:01:06.64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.86" />
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                    <SPLIT distance="75" swimtime="00:00:45.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="570" swimtime="00:00:30.45" resultid="110537" heatid="110834" lane="6" entrytime="00:00:30.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-11-19" firstname="Judyta" gender="F" lastname="Sołtyk" nation="POL" athleteid="110465">
              <RESULTS>
                <RESULT eventid="99457" points="461" reactiontime="+93" swimtime="00:05:03.46" resultid="110466" heatid="110839" lane="2" entrytime="00:05:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.33" />
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="75" swimtime="00:00:51.97" />
                    <SPLIT distance="100" swimtime="00:01:10.65" />
                    <SPLIT distance="125" swimtime="00:01:29.50" />
                    <SPLIT distance="150" swimtime="00:01:48.80" />
                    <SPLIT distance="175" swimtime="00:02:08.19" />
                    <SPLIT distance="200" swimtime="00:02:27.57" />
                    <SPLIT distance="225" swimtime="00:02:46.86" />
                    <SPLIT distance="250" swimtime="00:03:06.52" />
                    <SPLIT distance="275" swimtime="00:03:26.04" />
                    <SPLIT distance="300" swimtime="00:03:45.94" />
                    <SPLIT distance="325" swimtime="00:04:05.65" />
                    <SPLIT distance="350" swimtime="00:04:25.35" />
                    <SPLIT distance="375" swimtime="00:04:44.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Piotr" gender="M" lastname="Kister" nation="POL" athleteid="110385">
              <RESULTS>
                <RESULT eventid="98956" points="298" reactiontime="+82" swimtime="00:03:00.35" resultid="110386" heatid="110669" lane="1" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.35" />
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="75" swimtime="00:01:04.22" />
                    <SPLIT distance="100" swimtime="00:01:27.28" />
                    <SPLIT distance="125" swimtime="00:01:50.93" />
                    <SPLIT distance="150" swimtime="00:02:14.58" />
                    <SPLIT distance="175" swimtime="00:02:37.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="286" reactiontime="+77" swimtime="00:02:44.65" resultid="110387" heatid="110712" lane="5" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.28" />
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="75" swimtime="00:00:55.63" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="125" swimtime="00:01:38.07" />
                    <SPLIT distance="150" swimtime="00:02:00.15" />
                    <SPLIT distance="175" swimtime="00:02:22.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="332" swimtime="00:01:20.25" resultid="110388" heatid="110733" lane="9" entrytime="00:01:19.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.93" />
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="75" swimtime="00:00:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="354" reactiontime="+86" swimtime="00:00:30.80" resultid="110389" heatid="110747" lane="1" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="316" reactiontime="+68" swimtime="00:01:11.10" resultid="110390" heatid="110802" lane="4" entrytime="00:01:10.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.56" />
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="75" swimtime="00:00:51.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="339" reactiontime="+86" swimtime="00:00:36.21" resultid="110391" heatid="110831" lane="1" entrytime="00:00:35.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="110565">
              <RESULTS>
                <RESULT eventid="98940" status="DNS" swimtime="00:00:00.00" resultid="110566" heatid="110663" lane="9" entrytime="00:03:30.00" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="110567" heatid="110693" lane="0" entrytime="00:01:27.00" />
                <RESULT eventid="99089" points="263" reactiontime="+96" swimtime="00:01:37.22" resultid="110568" heatid="110723" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.01" />
                    <SPLIT distance="50" swimtime="00:00:45.67" />
                    <SPLIT distance="75" swimtime="00:01:11.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="274" swimtime="00:06:39.45" resultid="110569" heatid="110787" lane="9" entrytime="00:06:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.96" />
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="75" swimtime="00:01:08.23" />
                    <SPLIT distance="100" swimtime="00:01:36.89" />
                    <SPLIT distance="125" swimtime="00:02:03.33" />
                    <SPLIT distance="150" swimtime="00:02:27.02" />
                    <SPLIT distance="175" swimtime="00:02:50.72" />
                    <SPLIT distance="200" swimtime="00:03:13.76" />
                    <SPLIT distance="225" swimtime="00:03:41.14" />
                    <SPLIT distance="250" swimtime="00:04:08.52" />
                    <SPLIT distance="275" swimtime="00:04:35.98" />
                    <SPLIT distance="300" swimtime="00:05:03.79" />
                    <SPLIT distance="325" swimtime="00:05:28.69" />
                    <SPLIT distance="350" swimtime="00:05:52.78" />
                    <SPLIT distance="375" swimtime="00:06:16.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" status="DNS" swimtime="00:00:00.00" resultid="110570" heatid="110808" lane="0" entrytime="00:03:15.00" />
                <RESULT eventid="99457" status="DNS" swimtime="00:00:00.00" resultid="110571" heatid="110841" lane="6" entrytime="00:06:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Mateusz" gender="M" lastname="Burzawa" nation="POL" athleteid="110550">
              <RESULTS>
                <RESULT eventid="98798" points="502" reactiontime="+71" swimtime="00:00:25.49" resultid="110551" heatid="110610" lane="6" entrytime="00:00:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="507" reactiontime="+71" swimtime="00:02:17.41" resultid="110552" heatid="110628" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.23" />
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="75" swimtime="00:00:47.59" />
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                    <SPLIT distance="125" swimtime="00:01:25.62" />
                    <SPLIT distance="150" swimtime="00:01:45.69" />
                    <SPLIT distance="175" swimtime="00:02:02.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="404" reactiontime="+90" swimtime="00:00:30.05" resultid="110553" heatid="110659" lane="1" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="467" reactiontime="+77" swimtime="00:02:35.19" resultid="110554" heatid="110669" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="75" swimtime="00:00:54.58" />
                    <SPLIT distance="100" swimtime="00:01:14.62" />
                    <SPLIT distance="125" swimtime="00:01:34.83" />
                    <SPLIT distance="150" swimtime="00:01:55.09" />
                    <SPLIT distance="175" swimtime="00:02:15.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="474" reactiontime="+75" swimtime="00:01:11.28" resultid="110555" heatid="110733" lane="4" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.50" />
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="75" swimtime="00:00:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="572" swimtime="00:01:59.70" resultid="110556" heatid="110778" lane="0" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.03" />
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                    <SPLIT distance="75" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:00:58.32" />
                    <SPLIT distance="125" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:29.16" />
                    <SPLIT distance="175" swimtime="00:01:44.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Bogusław" gender="M" lastname="Ogrodnik" nation="POL" athleteid="110406">
              <RESULTS>
                <RESULT eventid="98798" points="214" reactiontime="+110" swimtime="00:00:33.85" resultid="110407" heatid="110600" lane="2" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="176" reactiontime="+110" swimtime="00:25:12.84" resultid="110408" heatid="110643" lane="5" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.85" />
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                    <SPLIT distance="75" swimtime="00:01:06.17" />
                    <SPLIT distance="100" swimtime="00:01:30.62" />
                    <SPLIT distance="125" swimtime="00:01:55.34" />
                    <SPLIT distance="150" swimtime="00:02:19.98" />
                    <SPLIT distance="175" swimtime="00:02:44.89" />
                    <SPLIT distance="200" swimtime="00:03:09.84" />
                    <SPLIT distance="225" swimtime="00:03:35.33" />
                    <SPLIT distance="250" swimtime="00:04:00.15" />
                    <SPLIT distance="275" swimtime="00:04:25.36" />
                    <SPLIT distance="300" swimtime="00:04:50.07" />
                    <SPLIT distance="325" swimtime="00:05:15.92" />
                    <SPLIT distance="350" swimtime="00:05:41.47" />
                    <SPLIT distance="375" swimtime="00:06:06.70" />
                    <SPLIT distance="400" swimtime="00:06:32.35" />
                    <SPLIT distance="425" swimtime="00:06:57.04" />
                    <SPLIT distance="450" swimtime="00:07:22.70" />
                    <SPLIT distance="475" swimtime="00:07:48.43" />
                    <SPLIT distance="500" swimtime="00:08:14.00" />
                    <SPLIT distance="525" swimtime="00:08:39.20" />
                    <SPLIT distance="550" swimtime="00:09:04.76" />
                    <SPLIT distance="575" swimtime="00:09:29.99" />
                    <SPLIT distance="600" swimtime="00:09:54.82" />
                    <SPLIT distance="625" swimtime="00:10:20.36" />
                    <SPLIT distance="650" swimtime="00:10:45.81" />
                    <SPLIT distance="675" swimtime="00:11:10.90" />
                    <SPLIT distance="700" swimtime="00:11:36.38" />
                    <SPLIT distance="725" swimtime="00:12:02.40" />
                    <SPLIT distance="750" swimtime="00:12:28.06" />
                    <SPLIT distance="775" swimtime="00:12:53.80" />
                    <SPLIT distance="800" swimtime="00:13:18.49" />
                    <SPLIT distance="825" swimtime="00:13:44.60" />
                    <SPLIT distance="850" swimtime="00:14:10.06" />
                    <SPLIT distance="875" swimtime="00:14:35.89" />
                    <SPLIT distance="900" swimtime="00:15:00.41" />
                    <SPLIT distance="925" swimtime="00:15:26.31" />
                    <SPLIT distance="950" swimtime="00:15:51.19" />
                    <SPLIT distance="975" swimtime="00:16:17.07" />
                    <SPLIT distance="1000" swimtime="00:16:41.69" />
                    <SPLIT distance="1025" swimtime="00:17:07.28" />
                    <SPLIT distance="1050" swimtime="00:17:32.09" />
                    <SPLIT distance="1075" swimtime="00:17:57.77" />
                    <SPLIT distance="1100" swimtime="00:18:22.45" />
                    <SPLIT distance="1125" swimtime="00:18:48.02" />
                    <SPLIT distance="1150" swimtime="00:19:13.48" />
                    <SPLIT distance="1175" swimtime="00:19:39.66" />
                    <SPLIT distance="1200" swimtime="00:20:05.90" />
                    <SPLIT distance="1225" swimtime="00:20:31.86" />
                    <SPLIT distance="1250" swimtime="00:20:57.70" />
                    <SPLIT distance="1275" swimtime="00:21:23.37" />
                    <SPLIT distance="1300" swimtime="00:21:48.92" />
                    <SPLIT distance="1325" swimtime="00:22:14.95" />
                    <SPLIT distance="1350" swimtime="00:22:40.87" />
                    <SPLIT distance="1375" swimtime="00:23:07.70" />
                    <SPLIT distance="1400" swimtime="00:23:33.87" />
                    <SPLIT distance="1425" swimtime="00:24:00.14" />
                    <SPLIT distance="1450" swimtime="00:24:26.22" />
                    <SPLIT distance="1475" swimtime="00:24:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="193" swimtime="00:01:17.67" resultid="110409" heatid="110681" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.92" />
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="75" swimtime="00:00:56.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="165" reactiontime="+101" swimtime="00:01:41.27" resultid="110410" heatid="110730" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.52" />
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="75" swimtime="00:01:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="158" swimtime="00:03:03.60" resultid="110411" heatid="110771" lane="6" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.75" />
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="75" swimtime="00:00:59.26" />
                    <SPLIT distance="100" swimtime="00:01:22.52" />
                    <SPLIT distance="125" swimtime="00:01:47.51" />
                    <SPLIT distance="150" swimtime="00:02:13.01" />
                    <SPLIT distance="175" swimtime="00:02:39.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="215" reactiontime="+99" swimtime="00:00:42.12" resultid="110412" heatid="110826" lane="3" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="143" swimtime="00:06:45.33" resultid="110413" heatid="110849" lane="9" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.38" />
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="75" swimtime="00:01:06.54" />
                    <SPLIT distance="100" swimtime="00:01:31.86" />
                    <SPLIT distance="125" swimtime="00:01:58.84" />
                    <SPLIT distance="150" swimtime="00:02:25.09" />
                    <SPLIT distance="175" swimtime="00:02:51.52" />
                    <SPLIT distance="200" swimtime="00:03:17.66" />
                    <SPLIT distance="225" swimtime="00:03:43.41" />
                    <SPLIT distance="250" swimtime="00:04:09.47" />
                    <SPLIT distance="275" swimtime="00:04:36.18" />
                    <SPLIT distance="300" swimtime="00:05:02.39" />
                    <SPLIT distance="325" swimtime="00:05:29.74" />
                    <SPLIT distance="350" swimtime="00:05:57.02" />
                    <SPLIT distance="375" swimtime="00:06:23.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="PAWEŁ" gender="M" lastname="CIESIELSKI" nation="POL" athleteid="110577">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="110578" heatid="110605" lane="0" entrytime="00:00:29.15" />
                <RESULT eventid="106277" points="288" reactiontime="+72" swimtime="00:01:08.00" resultid="110579" heatid="110682" lane="6" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                    <SPLIT distance="75" swimtime="00:00:48.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="278" reactiontime="+73" swimtime="00:01:17.55" resultid="110580" heatid="110701" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.10" />
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="75" swimtime="00:00:57.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="336" reactiontime="+66" swimtime="00:00:31.35" resultid="110581" heatid="110745" lane="4" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="110582" heatid="110829" lane="8" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Włodzimierz" gender="M" lastname="Zieliński" nation="POL" athleteid="110498">
              <RESULTS>
                <RESULT eventid="98798" status="WDR" swimtime="00:00:00.00" resultid="110499" heatid="110600" lane="3" entrytime="00:00:33.50" />
                <RESULT eventid="106256" status="WDR" swimtime="00:00:00.00" resultid="110500" heatid="110644" lane="2" entrytime="00:27:20.00" />
                <RESULT eventid="98924" status="WDR" swimtime="00:00:00.00" resultid="110501" heatid="110653" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="106277" status="WDR" swimtime="00:00:00.00" resultid="110502" heatid="110680" lane="4" entrytime="00:01:18.00" />
                <RESULT eventid="99218" status="WDR" swimtime="00:00:00.00" resultid="110503" heatid="110771" lane="0" entrytime="00:03:03.00" />
                <RESULT eventid="99393" status="WDR" swimtime="00:00:00.00" resultid="110504" heatid="110812" lane="0" entrytime="00:03:35.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="110505" heatid="110850" lane="6" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Marek" gender="M" lastname="Baranowski" nation="POL" swrid="4072629" athleteid="110380">
              <RESULTS>
                <RESULT eventid="98798" points="480" swimtime="00:00:25.87" resultid="110381" heatid="110611" lane="9" entrytime="00:00:25.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="478" swimtime="00:00:57.46" resultid="110382" heatid="110689" lane="0" entrytime="00:00:55.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.95" />
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                    <SPLIT distance="75" swimtime="00:00:42.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="500" reactiontime="+61" swimtime="00:02:05.14" resultid="110383" heatid="110776" lane="5" entrytime="00:02:14.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="75" swimtime="00:00:42.57" />
                    <SPLIT distance="100" swimtime="00:00:58.41" />
                    <SPLIT distance="125" swimtime="00:01:14.43" />
                    <SPLIT distance="150" swimtime="00:01:31.03" />
                    <SPLIT distance="175" swimtime="00:01:48.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="452" reactiontime="+75" swimtime="00:04:36.47" resultid="110384" heatid="110844" lane="3" entrytime="00:04:40.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.94" />
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="75" swimtime="00:00:46.45" />
                    <SPLIT distance="100" swimtime="00:01:03.40" />
                    <SPLIT distance="125" swimtime="00:01:20.81" />
                    <SPLIT distance="150" swimtime="00:01:38.47" />
                    <SPLIT distance="175" swimtime="00:01:56.11" />
                    <SPLIT distance="200" swimtime="00:02:14.01" />
                    <SPLIT distance="225" swimtime="00:02:31.64" />
                    <SPLIT distance="250" swimtime="00:02:49.38" />
                    <SPLIT distance="275" swimtime="00:03:07.10" />
                    <SPLIT distance="300" swimtime="00:03:24.92" />
                    <SPLIT distance="325" swimtime="00:03:42.84" />
                    <SPLIT distance="350" swimtime="00:04:01.10" />
                    <SPLIT distance="375" swimtime="00:04:18.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" swrid="4992696" athleteid="110447">
              <RESULTS>
                <RESULT eventid="98798" points="231" reactiontime="+88" swimtime="00:00:33.00" resultid="110448" heatid="110601" lane="8" entrytime="00:00:32.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="132" swimtime="00:14:30.29" resultid="110449" heatid="110637" lane="9" entrytime="00:13:12.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.08" />
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                    <SPLIT distance="75" swimtime="00:01:05.34" />
                    <SPLIT distance="100" swimtime="00:01:28.97" />
                    <SPLIT distance="125" swimtime="00:01:53.92" />
                    <SPLIT distance="150" swimtime="00:02:19.77" />
                    <SPLIT distance="175" swimtime="00:02:45.12" />
                    <SPLIT distance="200" swimtime="00:03:10.80" />
                    <SPLIT distance="225" swimtime="00:03:37.22" />
                    <SPLIT distance="250" swimtime="00:04:03.69" />
                    <SPLIT distance="275" swimtime="00:04:31.07" />
                    <SPLIT distance="300" swimtime="00:04:58.54" />
                    <SPLIT distance="325" swimtime="00:05:26.94" />
                    <SPLIT distance="350" swimtime="00:05:55.15" />
                    <SPLIT distance="375" swimtime="00:06:23.18" />
                    <SPLIT distance="400" swimtime="00:06:51.65" />
                    <SPLIT distance="425" swimtime="00:07:20.63" />
                    <SPLIT distance="450" swimtime="00:07:49.83" />
                    <SPLIT distance="475" swimtime="00:08:19.45" />
                    <SPLIT distance="500" swimtime="00:08:47.81" />
                    <SPLIT distance="525" swimtime="00:09:16.98" />
                    <SPLIT distance="550" swimtime="00:09:46.59" />
                    <SPLIT distance="575" swimtime="00:10:15.30" />
                    <SPLIT distance="600" swimtime="00:10:44.94" />
                    <SPLIT distance="625" swimtime="00:11:14.14" />
                    <SPLIT distance="650" swimtime="00:11:43.19" />
                    <SPLIT distance="675" swimtime="00:12:12.31" />
                    <SPLIT distance="700" swimtime="00:12:40.33" />
                    <SPLIT distance="725" swimtime="00:13:07.72" />
                    <SPLIT distance="750" swimtime="00:13:35.85" />
                    <SPLIT distance="775" swimtime="00:14:04.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="173" reactiontime="+80" swimtime="00:00:39.85" resultid="110450" heatid="110654" lane="4" entrytime="00:00:39.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="161" swimtime="00:01:33.03" resultid="110451" heatid="110698" lane="0" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.50" />
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                    <SPLIT distance="75" swimtime="00:01:09.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="157" swimtime="00:01:30.51" resultid="110452" heatid="110759" lane="3" entrytime="00:01:27.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.32" />
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                    <SPLIT distance="75" swimtime="00:01:07.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="134" swimtime="00:07:39.14" resultid="110453" heatid="110788" lane="4" entrytime="00:07:12.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.63" />
                    <SPLIT distance="50" swimtime="00:00:54.50" />
                    <SPLIT distance="75" swimtime="00:01:26.41" />
                    <SPLIT distance="100" swimtime="00:01:58.54" />
                    <SPLIT distance="125" swimtime="00:02:29.26" />
                    <SPLIT distance="150" swimtime="00:02:57.04" />
                    <SPLIT distance="175" swimtime="00:03:25.23" />
                    <SPLIT distance="200" swimtime="00:03:53.35" />
                    <SPLIT distance="225" swimtime="00:04:28.15" />
                    <SPLIT distance="250" swimtime="00:05:00.55" />
                    <SPLIT distance="275" swimtime="00:05:32.30" />
                    <SPLIT distance="300" swimtime="00:06:05.49" />
                    <SPLIT distance="325" swimtime="00:06:29.95" />
                    <SPLIT distance="350" swimtime="00:06:54.44" />
                    <SPLIT distance="375" swimtime="00:07:18.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="130" reactiontime="+91" swimtime="00:03:28.21" resultid="110454" heatid="110812" lane="2" entrytime="00:03:19.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.16" />
                    <SPLIT distance="75" swimtime="00:01:13.55" />
                    <SPLIT distance="100" swimtime="00:01:40.38" />
                    <SPLIT distance="125" swimtime="00:02:07.49" />
                    <SPLIT distance="150" swimtime="00:02:34.96" />
                    <SPLIT distance="175" swimtime="00:03:02.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="146" reactiontime="+90" swimtime="00:06:42.41" resultid="110455" heatid="110849" lane="8" entrytime="00:06:15.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.07" />
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                    <SPLIT distance="75" swimtime="00:01:06.26" />
                    <SPLIT distance="100" swimtime="00:01:30.59" />
                    <SPLIT distance="125" swimtime="00:01:56.16" />
                    <SPLIT distance="150" swimtime="00:02:22.49" />
                    <SPLIT distance="175" swimtime="00:02:48.83" />
                    <SPLIT distance="200" swimtime="00:03:14.30" />
                    <SPLIT distance="225" swimtime="00:03:40.92" />
                    <SPLIT distance="250" swimtime="00:04:07.35" />
                    <SPLIT distance="275" swimtime="00:04:34.52" />
                    <SPLIT distance="300" swimtime="00:05:01.19" />
                    <SPLIT distance="325" swimtime="00:05:28.82" />
                    <SPLIT distance="350" swimtime="00:05:54.65" />
                    <SPLIT distance="375" swimtime="00:06:19.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" swrid="4967127" athleteid="110524">
              <RESULTS>
                <RESULT eventid="98891" points="129" reactiontime="+106" swimtime="00:14:37.55" resultid="110525" heatid="110638" lane="5" entrytime="00:14:13.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.55" />
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                    <SPLIT distance="75" swimtime="00:01:10.89" />
                    <SPLIT distance="100" swimtime="00:01:37.55" />
                    <SPLIT distance="125" swimtime="00:02:04.26" />
                    <SPLIT distance="150" swimtime="00:02:32.12" />
                    <SPLIT distance="175" swimtime="00:02:59.65" />
                    <SPLIT distance="200" swimtime="00:03:26.91" />
                    <SPLIT distance="225" swimtime="00:03:54.19" />
                    <SPLIT distance="250" swimtime="00:04:21.83" />
                    <SPLIT distance="275" swimtime="00:04:49.80" />
                    <SPLIT distance="300" swimtime="00:05:17.50" />
                    <SPLIT distance="325" swimtime="00:05:44.99" />
                    <SPLIT distance="350" swimtime="00:06:13.05" />
                    <SPLIT distance="375" swimtime="00:06:41.18" />
                    <SPLIT distance="400" swimtime="00:07:09.42" />
                    <SPLIT distance="425" swimtime="00:07:38.08" />
                    <SPLIT distance="450" swimtime="00:08:06.13" />
                    <SPLIT distance="475" swimtime="00:08:34.50" />
                    <SPLIT distance="500" swimtime="00:09:03.12" />
                    <SPLIT distance="525" swimtime="00:09:31.20" />
                    <SPLIT distance="550" swimtime="00:09:59.35" />
                    <SPLIT distance="575" swimtime="00:10:27.92" />
                    <SPLIT distance="600" swimtime="00:10:56.46" />
                    <SPLIT distance="625" swimtime="00:11:25.01" />
                    <SPLIT distance="650" swimtime="00:11:53.48" />
                    <SPLIT distance="675" swimtime="00:12:21.64" />
                    <SPLIT distance="700" swimtime="00:12:49.81" />
                    <SPLIT distance="725" swimtime="00:13:18.40" />
                    <SPLIT distance="750" swimtime="00:13:45.99" />
                    <SPLIT distance="775" swimtime="00:14:13.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="130" reactiontime="+102" swimtime="00:01:28.68" resultid="110526" heatid="110679" lane="4" entrytime="00:01:29.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.16" />
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                    <SPLIT distance="75" swimtime="00:01:06.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="121" reactiontime="+94" swimtime="00:03:20.79" resultid="110527" heatid="110770" lane="2" entrytime="00:03:22.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.10" />
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                    <SPLIT distance="75" swimtime="00:01:10.13" />
                    <SPLIT distance="100" swimtime="00:01:35.50" />
                    <SPLIT distance="125" swimtime="00:02:02.36" />
                    <SPLIT distance="150" swimtime="00:02:29.94" />
                    <SPLIT distance="175" swimtime="00:02:57.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="119" reactiontime="+115" swimtime="00:07:11.19" resultid="110528" heatid="110851" lane="4" entrytime="00:07:11.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.33" />
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                    <SPLIT distance="75" swimtime="00:01:11.44" />
                    <SPLIT distance="100" swimtime="00:01:38.40" />
                    <SPLIT distance="125" swimtime="00:02:06.69" />
                    <SPLIT distance="150" swimtime="00:02:34.11" />
                    <SPLIT distance="175" swimtime="00:03:03.02" />
                    <SPLIT distance="200" swimtime="00:03:30.62" />
                    <SPLIT distance="225" swimtime="00:03:59.14" />
                    <SPLIT distance="250" swimtime="00:04:27.25" />
                    <SPLIT distance="275" swimtime="00:04:55.74" />
                    <SPLIT distance="300" swimtime="00:05:23.92" />
                    <SPLIT distance="325" swimtime="00:05:52.68" />
                    <SPLIT distance="350" swimtime="00:06:21.34" />
                    <SPLIT distance="375" swimtime="00:06:48.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="Edward" gender="M" lastname="Dziekoński" nation="POL" swrid="4992707" athleteid="110515">
              <RESULTS>
                <RESULT eventid="98798" points="130" reactiontime="+97" swimtime="00:00:39.95" resultid="110516" heatid="110596" lane="4" entrytime="00:00:40.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="117" reactiontime="+142" swimtime="00:15:05.63" resultid="110517" heatid="110638" lane="3" entrytime="00:15:09.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.12" />
                    <SPLIT distance="50" swimtime="00:00:49.42" />
                    <SPLIT distance="75" swimtime="00:01:17.03" />
                    <SPLIT distance="100" swimtime="00:01:45.14" />
                    <SPLIT distance="125" swimtime="00:02:13.87" />
                    <SPLIT distance="150" swimtime="00:02:42.31" />
                    <SPLIT distance="175" swimtime="00:03:11.17" />
                    <SPLIT distance="200" swimtime="00:03:40.01" />
                    <SPLIT distance="225" swimtime="00:04:09.01" />
                    <SPLIT distance="250" swimtime="00:04:37.16" />
                    <SPLIT distance="275" swimtime="00:05:05.35" />
                    <SPLIT distance="300" swimtime="00:05:33.83" />
                    <SPLIT distance="325" swimtime="00:06:02.72" />
                    <SPLIT distance="350" swimtime="00:06:31.66" />
                    <SPLIT distance="375" swimtime="00:07:00.44" />
                    <SPLIT distance="400" swimtime="00:07:29.15" />
                    <SPLIT distance="425" swimtime="00:07:57.85" />
                    <SPLIT distance="450" swimtime="00:08:26.92" />
                    <SPLIT distance="475" swimtime="00:08:56.21" />
                    <SPLIT distance="500" swimtime="00:09:25.02" />
                    <SPLIT distance="525" swimtime="00:09:53.95" />
                    <SPLIT distance="550" swimtime="00:10:22.85" />
                    <SPLIT distance="575" swimtime="00:10:51.65" />
                    <SPLIT distance="600" swimtime="00:11:20.59" />
                    <SPLIT distance="625" swimtime="00:11:49.15" />
                    <SPLIT distance="650" swimtime="00:12:17.18" />
                    <SPLIT distance="675" swimtime="00:12:45.76" />
                    <SPLIT distance="700" swimtime="00:13:14.53" />
                    <SPLIT distance="725" swimtime="00:13:43.05" />
                    <SPLIT distance="750" swimtime="00:14:11.26" />
                    <SPLIT distance="775" swimtime="00:14:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="81" reactiontime="+104" swimtime="00:00:51.33" resultid="110518" heatid="110652" lane="5" entrytime="00:00:50.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="94" reactiontime="+106" swimtime="00:01:51.07" resultid="110519" heatid="110696" lane="4" entrytime="00:01:55.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.69" />
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                    <SPLIT distance="75" swimtime="00:01:25.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="120" swimtime="00:00:44.08" resultid="110520" heatid="110743" lane="9" entrytime="00:00:43.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="113" reactiontime="+107" swimtime="00:03:24.96" resultid="110521" heatid="110770" lane="8" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.59" />
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="75" swimtime="00:01:11.64" />
                    <SPLIT distance="100" swimtime="00:01:38.13" />
                    <SPLIT distance="125" swimtime="00:02:05.44" />
                    <SPLIT distance="150" swimtime="00:02:32.70" />
                    <SPLIT distance="175" swimtime="00:02:59.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="70" swimtime="00:01:57.16" resultid="110522" heatid="110799" lane="9" entrytime="00:01:57.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.63" />
                    <SPLIT distance="50" swimtime="00:00:54.32" />
                    <SPLIT distance="75" swimtime="00:01:25.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="114" swimtime="00:07:17.51" resultid="110523" heatid="110851" lane="2" entrytime="00:07:31.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.20" />
                    <SPLIT distance="50" swimtime="00:00:47.89" />
                    <SPLIT distance="75" swimtime="00:01:14.57" />
                    <SPLIT distance="100" swimtime="00:01:41.54" />
                    <SPLIT distance="125" swimtime="00:02:09.24" />
                    <SPLIT distance="150" swimtime="00:02:37.52" />
                    <SPLIT distance="175" swimtime="00:03:05.62" />
                    <SPLIT distance="200" swimtime="00:03:34.60" />
                    <SPLIT distance="225" swimtime="00:04:03.20" />
                    <SPLIT distance="250" swimtime="00:04:31.09" />
                    <SPLIT distance="275" swimtime="00:04:59.09" />
                    <SPLIT distance="300" swimtime="00:05:26.68" />
                    <SPLIT distance="325" swimtime="00:05:54.74" />
                    <SPLIT distance="350" swimtime="00:06:22.90" />
                    <SPLIT distance="375" swimtime="00:06:51.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-18" firstname="Kazimierz" gender="M" lastname="Sinicki" nation="POL" athleteid="110538">
              <RESULTS>
                <RESULT eventid="98798" points="309" reactiontime="+74" swimtime="00:00:29.94" resultid="110539" heatid="110603" lane="8" entrytime="00:00:30.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="287" reactiontime="+99" swimtime="00:01:08.08" resultid="110540" heatid="110683" lane="1" entrytime="00:01:07.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.48" />
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="75" swimtime="00:00:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="243" reactiontime="+84" swimtime="00:00:34.90" resultid="110541" heatid="110743" lane="4" entrytime="00:00:35.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Andrzej" gender="M" lastname="Fajdasz" nation="POL" athleteid="110392">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="110393" heatid="110603" lane="2" entrytime="00:00:30.35" />
                <RESULT eventid="98830" points="224" reactiontime="+86" swimtime="00:03:00.38" resultid="110394" heatid="110622" lane="7" entrytime="00:03:05.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="75" swimtime="00:01:01.98" />
                    <SPLIT distance="100" swimtime="00:01:25.71" />
                    <SPLIT distance="125" swimtime="00:01:51.96" />
                    <SPLIT distance="150" swimtime="00:02:18.56" />
                    <SPLIT distance="175" swimtime="00:02:40.25" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4" eventid="106277" status="DSQ" swimtime="00:00:00.00" resultid="110395" heatid="110686" lane="2" entrytime="00:01:01.20" />
                <RESULT eventid="98988" points="269" swimtime="00:01:18.42" resultid="110396" heatid="110700" lane="0" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.60" />
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="75" swimtime="00:01:01.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="224" reactiontime="+92" swimtime="00:01:20.50" resultid="110397" heatid="110760" lane="7" entrytime="00:01:20.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.83" />
                    <SPLIT distance="50" swimtime="00:01:20.49" />
                    <SPLIT distance="75" swimtime="00:01:00.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="289" reactiontime="+89" swimtime="00:02:30.17" resultid="110398" heatid="110772" lane="5" entrytime="00:02:40.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.22" />
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="75" swimtime="00:00:52.99" />
                    <SPLIT distance="100" swimtime="00:01:12.31" />
                    <SPLIT distance="125" swimtime="00:01:31.64" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                    <SPLIT distance="175" swimtime="00:02:11.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="216" reactiontime="+87" swimtime="00:02:56.03" resultid="110399" heatid="110813" lane="7" entrytime="00:02:58.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.97" />
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="75" swimtime="00:01:02.53" />
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                    <SPLIT distance="125" swimtime="00:01:47.98" />
                    <SPLIT distance="150" swimtime="00:02:11.35" />
                    <SPLIT distance="175" swimtime="00:02:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="258" swimtime="00:05:33.13" resultid="110400" heatid="110848" lane="6" entrytime="00:05:48.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.74" />
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="75" swimtime="00:00:54.90" />
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="125" swimtime="00:01:35.40" />
                    <SPLIT distance="150" swimtime="00:01:56.37" />
                    <SPLIT distance="175" swimtime="00:02:17.28" />
                    <SPLIT distance="200" swimtime="00:02:38.39" />
                    <SPLIT distance="225" swimtime="00:02:59.54" />
                    <SPLIT distance="250" swimtime="00:03:20.97" />
                    <SPLIT distance="275" swimtime="00:03:42.65" />
                    <SPLIT distance="300" swimtime="00:04:04.89" />
                    <SPLIT distance="325" swimtime="00:04:26.90" />
                    <SPLIT distance="350" swimtime="00:04:49.34" />
                    <SPLIT distance="375" swimtime="00:05:11.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-06-30" firstname="Alan" gender="M" lastname="Bistron" nation="POL" athleteid="110369">
              <RESULTS>
                <RESULT eventid="98798" points="247" reactiontime="+66" swimtime="00:00:32.28" resultid="110370" heatid="110598" lane="4" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" swrid="4186249" athleteid="110478">
              <RESULTS>
                <RESULT eventid="98798" points="392" swimtime="00:00:27.68" resultid="110479" heatid="110607" lane="9" entrytime="00:00:28.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="359" reactiontime="+95" swimtime="00:02:34.19" resultid="110480" heatid="110625" lane="2" entrytime="00:02:38.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.65" />
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="75" swimtime="00:00:52.53" />
                    <SPLIT distance="100" swimtime="00:01:12.08" />
                    <SPLIT distance="125" swimtime="00:01:34.67" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                    <SPLIT distance="175" swimtime="00:02:16.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="400" reactiontime="+77" swimtime="00:00:29.57" resultid="110481" heatid="110748" lane="8" entrytime="00:00:30.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="110482" heatid="110775" lane="2" entrytime="00:02:20.25" />
                <RESULT eventid="106277" points="395" reactiontime="+83" swimtime="00:01:01.21" resultid="110483" heatid="110685" lane="7" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.24" />
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="75" swimtime="00:00:45.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z2/G3" eventid="98988" status="DSQ" swimtime="00:00:00.00" resultid="110484" heatid="110703" lane="9" entrytime="00:01:11.25" />
                <RESULT eventid="99361" points="354" reactiontime="+95" swimtime="00:01:08.43" resultid="110485" heatid="110803" lane="1" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.69" />
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="75" swimtime="00:00:50.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="333" swimtime="00:00:36.41" resultid="110486" heatid="110829" lane="4" entrytime="00:00:37.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-06-06" firstname="Jolanta" gender="F" lastname="Lipińska" nation="POL" athleteid="110471">
              <RESULTS>
                <RESULT eventid="98814" points="25" reactiontime="+129" swimtime="00:06:53.13" resultid="110472" heatid="110614" lane="1" entrytime="00:06:42.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:48.12" />
                    <SPLIT distance="50" swimtime="00:01:45.87" />
                    <SPLIT distance="75" swimtime="00:02:35.39" />
                    <SPLIT distance="100" swimtime="00:03:25.12" />
                    <SPLIT distance="125" swimtime="00:04:22.67" />
                    <SPLIT distance="150" swimtime="00:05:19.14" />
                    <SPLIT distance="175" swimtime="00:06:07.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="47" reactiontime="+126" swimtime="00:06:11.32" resultid="110473" heatid="110661" lane="7" entrytime="00:05:49.73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:42.48" />
                    <SPLIT distance="50" swimtime="00:01:27.78" />
                    <SPLIT distance="75" swimtime="00:02:16.05" />
                    <SPLIT distance="100" swimtime="00:03:03.73" />
                    <SPLIT distance="125" swimtime="00:03:52.78" />
                    <SPLIT distance="150" swimtime="00:04:40.86" />
                    <SPLIT distance="175" swimtime="00:05:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="43" reactiontime="+144" swimtime="00:02:57.71" resultid="110474" heatid="110721" lane="1" entrytime="00:02:50.78">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:37.82" />
                    <SPLIT distance="50" swimtime="00:01:23.09" />
                    <SPLIT distance="75" swimtime="00:02:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="31" reactiontime="+52" swimtime="00:02:53.62" resultid="110475" heatid="110753" lane="2" entrytime="00:02:56.78">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:38.96" />
                    <SPLIT distance="50" swimtime="00:01:22.88" />
                    <SPLIT distance="75" swimtime="00:02:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="33" reactiontime="+69" swimtime="00:06:11.27" resultid="110476" heatid="110806" lane="2" entrytime="00:06:05.74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:42.26" />
                    <SPLIT distance="50" swimtime="00:01:26.02" />
                    <SPLIT distance="75" swimtime="00:02:13.94" />
                    <SPLIT distance="100" swimtime="00:03:00.84" />
                    <SPLIT distance="125" swimtime="00:03:49.26" />
                    <SPLIT distance="150" swimtime="00:04:36.46" />
                    <SPLIT distance="175" swimtime="00:05:26.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="58" reactiontime="+128" swimtime="00:01:14.23" resultid="110477" heatid="110817" lane="3" entrytime="00:01:16.16">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="31" reactiontime="+78" swimtime="00:03:00.23" resultid="110583" heatid="110690" lane="6" entrytime="00:02:58.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:46.80" />
                    <SPLIT distance="50" swimtime="00:01:29.80" />
                    <SPLIT distance="75" swimtime="00:02:16.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-02" firstname="Janusz" gender="M" lastname="Płonka" nation="POL" athleteid="110361">
              <RESULTS>
                <RESULT eventid="98830" points="56" reactiontime="+114" swimtime="00:04:44.99" resultid="110362" heatid="110619" lane="3" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.67" />
                    <SPLIT distance="50" swimtime="00:01:01.69" />
                    <SPLIT distance="75" swimtime="00:01:40.52" />
                    <SPLIT distance="100" swimtime="00:02:20.69" />
                    <SPLIT distance="125" swimtime="00:03:02.39" />
                    <SPLIT distance="150" swimtime="00:03:43.43" />
                    <SPLIT distance="175" swimtime="00:04:16.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="62" reactiontime="+103" swimtime="00:05:04.25" resultid="110363" heatid="110665" lane="3" entrytime="00:05:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.40" />
                    <SPLIT distance="50" swimtime="00:01:11.50" />
                    <SPLIT distance="75" swimtime="00:01:52.91" />
                    <SPLIT distance="100" swimtime="00:02:32.90" />
                    <SPLIT distance="125" swimtime="00:03:12.81" />
                    <SPLIT distance="150" swimtime="00:03:53.16" />
                    <SPLIT distance="175" swimtime="00:04:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="36" reactiontime="+107" swimtime="00:05:25.87" resultid="110364" heatid="110709" lane="4" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.60" />
                    <SPLIT distance="50" swimtime="00:01:08.71" />
                    <SPLIT distance="75" swimtime="00:01:51.27" />
                    <SPLIT distance="100" swimtime="00:02:34.02" />
                    <SPLIT distance="125" swimtime="00:03:15.76" />
                    <SPLIT distance="175" swimtime="00:04:43.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="76" reactiontime="+99" swimtime="00:00:51.38" resultid="110365" heatid="110742" lane="8" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="52" reactiontime="+84" swimtime="00:02:10.70" resultid="110366" heatid="110758" lane="8" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.10" />
                    <SPLIT distance="50" swimtime="00:01:06.31" />
                    <SPLIT distance="75" swimtime="00:01:38.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="40" reactiontime="+117" swimtime="00:02:20.76" resultid="110367" heatid="110798" lane="7" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.40" />
                    <SPLIT distance="50" swimtime="00:01:05.86" />
                    <SPLIT distance="75" swimtime="00:01:44.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="83" reactiontime="+117" swimtime="00:00:57.87" resultid="110368" heatid="110824" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="110487">
              <RESULTS>
                <RESULT eventid="98798" points="264" reactiontime="+89" swimtime="00:00:31.57" resultid="110488" heatid="110601" lane="6" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106256" points="192" swimtime="00:24:29.86" resultid="110489" heatid="110643" lane="6" entrytime="00:25:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.45" />
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="75" swimtime="00:01:05.86" />
                    <SPLIT distance="100" swimtime="00:01:30.25" />
                    <SPLIT distance="125" swimtime="00:01:54.61" />
                    <SPLIT distance="150" swimtime="00:02:18.85" />
                    <SPLIT distance="175" swimtime="00:02:44.28" />
                    <SPLIT distance="200" swimtime="00:03:07.95" />
                    <SPLIT distance="225" swimtime="00:03:32.87" />
                    <SPLIT distance="250" swimtime="00:03:57.89" />
                    <SPLIT distance="275" swimtime="00:04:22.87" />
                    <SPLIT distance="300" swimtime="00:04:47.87" />
                    <SPLIT distance="325" swimtime="00:05:12.60" />
                    <SPLIT distance="350" swimtime="00:05:37.15" />
                    <SPLIT distance="375" swimtime="00:06:01.37" />
                    <SPLIT distance="400" swimtime="00:06:27.35" />
                    <SPLIT distance="425" swimtime="00:06:52.79" />
                    <SPLIT distance="450" swimtime="00:07:17.27" />
                    <SPLIT distance="475" swimtime="00:07:41.87" />
                    <SPLIT distance="500" swimtime="00:08:06.06" />
                    <SPLIT distance="525" swimtime="00:08:32.16" />
                    <SPLIT distance="550" swimtime="00:08:57.20" />
                    <SPLIT distance="575" swimtime="00:09:22.22" />
                    <SPLIT distance="600" swimtime="00:09:47.84" />
                    <SPLIT distance="625" swimtime="00:10:12.20" />
                    <SPLIT distance="650" swimtime="00:11:27.90" />
                    <SPLIT distance="675" swimtime="00:11:02.82" />
                    <SPLIT distance="700" swimtime="00:12:17.77" />
                    <SPLIT distance="725" swimtime="00:11:52.96" />
                    <SPLIT distance="750" swimtime="00:13:07.07" />
                    <SPLIT distance="775" swimtime="00:12:42.38" />
                    <SPLIT distance="800" swimtime="00:13:56.32" />
                    <SPLIT distance="825" swimtime="00:13:31.73" />
                    <SPLIT distance="850" swimtime="00:14:44.75" />
                    <SPLIT distance="875" swimtime="00:14:20.71" />
                    <SPLIT distance="900" swimtime="00:15:34.69" />
                    <SPLIT distance="925" swimtime="00:15:09.13" />
                    <SPLIT distance="950" swimtime="00:16:24.52" />
                    <SPLIT distance="975" swimtime="00:15:59.73" />
                    <SPLIT distance="1000" swimtime="00:17:14.06" />
                    <SPLIT distance="1025" swimtime="00:16:49.25" />
                    <SPLIT distance="1075" swimtime="00:17:38.61" />
                    <SPLIT distance="1125" swimtime="00:18:29.50" />
                    <SPLIT distance="1150" swimtime="00:18:54.03" />
                    <SPLIT distance="1175" swimtime="00:19:18.62" />
                    <SPLIT distance="1200" swimtime="00:19:43.62" />
                    <SPLIT distance="1225" swimtime="00:20:08.59" />
                    <SPLIT distance="1250" swimtime="00:20:32.96" />
                    <SPLIT distance="1275" swimtime="00:20:56.76" />
                    <SPLIT distance="1300" swimtime="00:21:20.01" />
                    <SPLIT distance="1325" swimtime="00:21:44.14" />
                    <SPLIT distance="1375" swimtime="00:22:33.28" />
                    <SPLIT distance="1400" swimtime="00:22:57.88" />
                    <SPLIT distance="1425" swimtime="00:23:21.45" />
                    <SPLIT distance="1450" swimtime="00:23:46.33" />
                    <SPLIT distance="1475" swimtime="00:24:09.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="110490" heatid="110654" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="106277" points="247" reactiontime="+89" swimtime="00:01:11.57" resultid="110491" heatid="110681" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.52" />
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="75" swimtime="00:00:52.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="176" reactiontime="+109" swimtime="00:00:38.89" resultid="110492" heatid="110743" lane="2" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="207" reactiontime="+103" swimtime="00:02:47.77" resultid="110493" heatid="110772" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.98" />
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="75" swimtime="00:00:59.04" />
                    <SPLIT distance="100" swimtime="00:01:20.49" />
                    <SPLIT distance="125" swimtime="00:01:42.22" />
                    <SPLIT distance="150" swimtime="00:02:04.83" />
                    <SPLIT distance="175" swimtime="00:02:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="110494" heatid="110849" lane="5" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-03-13" firstname="Konrad" gender="M" lastname="Szydło" nation="POL" athleteid="110456">
              <RESULTS>
                <RESULT eventid="98798" points="314" reactiontime="+90" swimtime="00:00:29.80" resultid="110457" heatid="110604" lane="2" entrytime="00:00:29.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="239" swimtime="00:02:56.60" resultid="110458" heatid="110622" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.20" />
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="75" swimtime="00:01:01.28" />
                    <SPLIT distance="100" swimtime="00:01:23.21" />
                    <SPLIT distance="125" swimtime="00:01:50.11" />
                    <SPLIT distance="150" swimtime="00:02:17.07" />
                    <SPLIT distance="175" swimtime="00:02:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="226" reactiontime="+78" swimtime="00:00:36.43" resultid="110459" heatid="110655" lane="7" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" points="314" reactiontime="+96" swimtime="00:01:06.06" resultid="110460" heatid="110683" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.05" />
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="75" swimtime="00:00:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="228" reactiontime="+85" swimtime="00:01:19.97" resultid="110461" heatid="110759" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.35" />
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="75" swimtime="00:00:59.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="306" reactiontime="+88" swimtime="00:02:27.45" resultid="110462" heatid="110772" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.78" />
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="75" swimtime="00:00:52.28" />
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                    <SPLIT distance="125" swimtime="00:01:30.67" />
                    <SPLIT distance="150" swimtime="00:01:50.74" />
                    <SPLIT distance="175" swimtime="00:02:09.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="220" reactiontime="+73" swimtime="00:02:54.78" resultid="110463" heatid="110812" lane="6" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.14" />
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="75" swimtime="00:01:03.69" />
                    <SPLIT distance="100" swimtime="00:01:26.13" />
                    <SPLIT distance="125" swimtime="00:01:48.59" />
                    <SPLIT distance="150" swimtime="00:02:10.94" />
                    <SPLIT distance="175" swimtime="00:02:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="291" reactiontime="+90" swimtime="00:05:20.03" resultid="110464" heatid="110848" lane="5" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="75" swimtime="00:00:54.36" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="125" swimtime="00:01:34.46" />
                    <SPLIT distance="150" swimtime="00:01:54.61" />
                    <SPLIT distance="175" swimtime="00:02:15.19" />
                    <SPLIT distance="200" swimtime="00:02:35.86" />
                    <SPLIT distance="225" swimtime="00:02:56.56" />
                    <SPLIT distance="250" swimtime="00:03:17.34" />
                    <SPLIT distance="275" swimtime="00:03:38.38" />
                    <SPLIT distance="300" swimtime="00:03:59.50" />
                    <SPLIT distance="325" swimtime="00:04:20.55" />
                    <SPLIT distance="350" swimtime="00:04:41.54" />
                    <SPLIT distance="375" swimtime="00:05:01.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Bernard" gender="M" lastname="Wierzbik" nation="POL" athleteid="110572">
              <RESULTS>
                <RESULT eventid="99020" points="167" swimtime="00:03:16.84" resultid="110573" heatid="110711" lane="0" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.90" />
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="75" swimtime="00:01:02.44" />
                    <SPLIT distance="100" swimtime="00:01:28.02" />
                    <SPLIT distance="125" swimtime="00:01:54.75" />
                    <SPLIT distance="150" swimtime="00:02:22.56" />
                    <SPLIT distance="175" swimtime="00:02:50.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="263" reactiontime="+97" swimtime="00:00:33.99" resultid="110574" heatid="110744" lane="3" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="220" swimtime="00:06:30.09" resultid="110575" heatid="110789" lane="0" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.00" />
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="75" swimtime="00:01:01.18" />
                    <SPLIT distance="100" swimtime="00:01:25.79" />
                    <SPLIT distance="150" swimtime="00:02:17.70" />
                    <SPLIT distance="200" swimtime="00:03:08.13" />
                    <SPLIT distance="225" swimtime="00:03:35.06" />
                    <SPLIT distance="250" swimtime="00:04:01.95" />
                    <SPLIT distance="275" swimtime="00:04:29.49" />
                    <SPLIT distance="300" swimtime="00:04:58.33" />
                    <SPLIT distance="325" swimtime="00:05:21.98" />
                    <SPLIT distance="350" swimtime="00:05:45.54" />
                    <SPLIT distance="375" swimtime="00:06:09.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="219" reactiontime="+92" swimtime="00:01:20.26" resultid="110576" heatid="110800" lane="5" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.38" />
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="75" swimtime="00:00:57.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Paweł" gender="M" lastname="Marudziński" nation="POL" athleteid="110557">
              <RESULTS>
                <RESULT eventid="98830" points="278" reactiontime="+88" swimtime="00:02:47.78" resultid="110558" heatid="110623" lane="8" entrytime="00:02:57.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.48" />
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="75" swimtime="00:00:54.85" />
                    <SPLIT distance="100" swimtime="00:01:16.73" />
                    <SPLIT distance="125" swimtime="00:01:40.62" />
                    <SPLIT distance="150" swimtime="00:02:04.90" />
                    <SPLIT distance="175" swimtime="00:02:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="272" reactiontime="+95" swimtime="00:03:05.90" resultid="110559" heatid="110667" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.16" />
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="75" swimtime="00:01:03.73" />
                    <SPLIT distance="100" swimtime="00:01:27.85" />
                    <SPLIT distance="125" swimtime="00:01:52.73" />
                    <SPLIT distance="150" swimtime="00:02:17.73" />
                    <SPLIT distance="175" swimtime="00:02:42.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="311" reactiontime="+88" swimtime="00:01:14.71" resultid="110560" heatid="110701" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.11" />
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="75" swimtime="00:00:56.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="289" reactiontime="+68" swimtime="00:01:24.05" resultid="110561" heatid="110732" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.75" />
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="75" swimtime="00:01:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="351" reactiontime="+89" swimtime="00:00:30.90" resultid="110562" heatid="110744" lane="4" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="110563" heatid="110803" lane="9" entrytime="00:01:10.00" />
                <RESULT eventid="99425" points="297" reactiontime="+101" swimtime="00:00:37.84" resultid="110564" heatid="110826" lane="2" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Adriana" gender="F" lastname="Hofman" nation="POL" swrid="4236095" athleteid="110401">
              <RESULTS>
                <RESULT eventid="98777" points="470" reactiontime="+82" swimtime="00:00:29.88" resultid="110402" heatid="110591" lane="1" entrytime="00:00:32.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="469" reactiontime="+76" swimtime="00:01:20.25" resultid="110403" heatid="110725" lane="8" entrytime="00:01:22.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.24" />
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                    <SPLIT distance="75" swimtime="00:00:59.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="436" swimtime="00:01:14.71" resultid="110404" heatid="110693" lane="4" entrytime="00:01:20.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.70" />
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="75" swimtime="00:00:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="550" reactiontime="+75" swimtime="00:00:35.14" resultid="110405" heatid="110823" lane="7" entrytime="00:00:36.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Patryk" gender="M" lastname="Suchodolski" nation="POL" athleteid="110506">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="110507" heatid="110610" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="110508" heatid="110624" lane="7" entrytime="00:02:45.00" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="110509" heatid="110660" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="110510" heatid="110670" lane="7" entrytime="00:02:40.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="110511" heatid="110734" lane="7" entrytime="00:01:10.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="110512" heatid="110750" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="110513" heatid="110804" lane="2" entrytime="00:01:05.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="110514" heatid="110834" lane="3" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Weronika" gender="F" lastname="Kabut" nation="POL" athleteid="110371">
              <RESULTS>
                <RESULT eventid="98777" points="473" reactiontime="+78" swimtime="00:00:29.82" resultid="110372" heatid="110592" lane="0" entrytime="00:00:30.14">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98814" points="356" reactiontime="+87" swimtime="00:02:51.81" resultid="110373" heatid="110617" lane="3" entrytime="00:02:53.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.37" />
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="75" swimtime="00:00:58.63" />
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="125" swimtime="00:01:45.55" />
                    <SPLIT distance="150" swimtime="00:02:10.55" />
                    <SPLIT distance="175" swimtime="00:02:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="465" reactiontime="+69" swimtime="00:01:05.71" resultid="110374" heatid="110675" lane="5" entrytime="00:01:07.39">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.93" />
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="75" swimtime="00:00:48.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="382" reactiontime="+61" swimtime="00:01:18.08" resultid="110375" heatid="110694" lane="6" entrytime="00:01:18.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.05" />
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="75" swimtime="00:01:00.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="380" reactiontime="+89" swimtime="00:00:33.65" resultid="110376" heatid="110739" lane="2" entrytime="00:00:34.85">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="413" swimtime="00:02:28.71" resultid="110377" heatid="110767" lane="6" entrytime="00:02:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.32" />
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="75" swimtime="00:00:51.30" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="125" swimtime="00:01:29.74" />
                    <SPLIT distance="150" swimtime="00:01:49.72" />
                    <SPLIT distance="175" swimtime="00:02:09.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="352" reactiontime="+87" swimtime="00:00:40.78" resultid="110378" heatid="110821" lane="7" entrytime="00:00:40.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="350" swimtime="00:05:32.54" resultid="110379" heatid="110839" lane="9" entrytime="00:05:37.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.87" />
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="75" swimtime="00:00:53.54" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="125" swimtime="00:01:34.51" />
                    <SPLIT distance="150" swimtime="00:01:55.90" />
                    <SPLIT distance="175" swimtime="00:02:16.90" />
                    <SPLIT distance="200" swimtime="00:02:38.99" />
                    <SPLIT distance="225" swimtime="00:03:00.66" />
                    <SPLIT distance="250" swimtime="00:03:22.65" />
                    <SPLIT distance="275" swimtime="00:03:44.50" />
                    <SPLIT distance="300" swimtime="00:04:07.11" />
                    <SPLIT distance="325" swimtime="00:04:28.64" />
                    <SPLIT distance="350" swimtime="00:04:50.88" />
                    <SPLIT distance="375" swimtime="00:05:12.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Piotr" gender="M" lastname="Urbańczyk" nation="POL" swrid="4186188" athleteid="110467">
              <RESULTS>
                <RESULT eventid="98924" points="456" reactiontime="+79" swimtime="00:00:28.85" resultid="110468" heatid="110660" lane="2" entrytime="00:00:28.47">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="480" reactiontime="+69" swimtime="00:01:02.46" resultid="110469" heatid="110763" lane="6" entrytime="00:01:00.94">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.08" />
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="75" swimtime="00:00:47.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="419" reactiontime="+71" swimtime="00:02:21.12" resultid="110470" heatid="110816" lane="6" entrytime="00:02:15.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.94" />
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="75" swimtime="00:00:50.10" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="125" swimtime="00:01:26.81" />
                    <SPLIT distance="150" swimtime="00:01:45.40" />
                    <SPLIT distance="175" swimtime="00:02:03.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-11" firstname="Paweł" gender="M" lastname="Adamowicz" nation="POL" athleteid="110425">
              <RESULTS>
                <RESULT eventid="98798" points="71" reactiontime="+82" swimtime="00:00:48.84" resultid="110426" heatid="110596" lane="5" entrytime="00:00:41.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106277" status="DNS" swimtime="00:00:00.00" resultid="110427" heatid="110677" lane="3" />
                <RESULT eventid="99091" points="162" reactiontime="+79" swimtime="00:01:41.91" resultid="110428" heatid="110728" lane="5" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.45" />
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="75" swimtime="00:01:15.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="180" reactiontime="+87" swimtime="00:00:44.70" resultid="110429" heatid="110826" lane="1" entrytime="00:00:45.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Aleksandra" gender="F" lastname="Mazurkiewicz" nation="POL" swrid="4170963" athleteid="110439">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="110440" heatid="110592" lane="6" entrytime="00:00:29.50" />
                <RESULT eventid="106294" status="DNS" swimtime="00:00:00.00" resultid="110441" heatid="110650" lane="0" entrytime="00:00:33.15" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="110442" heatid="110675" lane="6" entrytime="00:01:09.50" />
                <RESULT eventid="99089" status="DNS" swimtime="00:00:00.00" resultid="110443" heatid="110725" lane="7" entrytime="00:01:22.00" />
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="110444" heatid="110756" lane="2" entrytime="00:01:13.44" />
                <RESULT eventid="99377" status="DNS" swimtime="00:00:00.00" resultid="110445" heatid="110809" lane="3" entrytime="00:02:38.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="110446" heatid="110822" lane="6" entrytime="00:00:38.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="1077" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:22.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:43.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1103" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:11:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:21:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.25">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:57.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:07.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:22.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:42.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1075" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:13:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:52.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:22.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1101" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:11:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:22:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:22.50">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:05.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:25.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:52.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1073" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:47.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1099" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:12:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:22:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:12.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:12.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:52.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1071" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:15:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:50.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:50.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:07.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1097" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:12:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:37.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1069" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:15:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:50.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:52.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1095" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1067" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:16:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1093" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:13:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:52.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1065" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:16:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:57.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1091" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1063" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:17:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:52.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1089" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:15:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1059" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:20:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:21.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1085" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:17:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:02.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1057" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:21:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1083" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:18:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1615" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:19:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:57.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1617" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:23:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1619" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="89" agemin="85" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:20:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1621" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="89" agemin="85" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:24:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1623" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="94" agemin="90" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:23:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1625" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="94" agemin="90" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:26:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1627" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="95" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:27:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1629" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="95" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:29:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1061" course="LCM" gender="F" type="DEFAULT">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:15:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:12.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1087" course="LCM" gender="M" type="DEFAULT">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:16:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="KS Warszawianka" version="11.76727">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Warszawa" name="LETNIE OTWARTE MISTRZOSTWA POLSKI W PŁYWANIU W KATEGORIACH MASTERS" course="LCM" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2023-06-02" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Warszawa" nation="POL" />
      <POINTTABLE pointtableid="3123" name="FINA Master Point Scoring" version="2023" />
      <SESSIONS>
        <SESSION date="2023-06-02" daytime="14:00" endtime="18:39" name="I BLOK" number="1" warmupfrom="13:00" warmupuntil="13:55">
          <EVENTS>
            <EVENT eventid="1059" daytime="14:00" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4008" />
                    <RANKING order="2" place="2" resultid="2644" />
                    <RANKING order="3" place="3" resultid="3641" />
                    <RANKING order="4" place="4" resultid="3097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3423" />
                    <RANKING order="2" place="2" resultid="3956" />
                    <RANKING order="3" place="3" resultid="3739" />
                    <RANKING order="4" place="4" resultid="3378" />
                    <RANKING order="5" place="5" resultid="2743" />
                    <RANKING order="6" place="6" resultid="1822" />
                    <RANKING order="7" place="7" resultid="3771" />
                    <RANKING order="8" place="8" resultid="3947" />
                    <RANKING order="9" place="9" resultid="3068" />
                    <RANKING order="10" place="-1" resultid="3254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3583" />
                    <RANKING order="2" place="2" resultid="2165" />
                    <RANKING order="3" place="3" resultid="3175" />
                    <RANKING order="4" place="4" resultid="2767" />
                    <RANKING order="5" place="5" resultid="3232" />
                    <RANKING order="6" place="6" resultid="3180" />
                    <RANKING order="7" place="7" resultid="3459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3466" />
                    <RANKING order="2" place="2" resultid="2630" />
                    <RANKING order="3" place="3" resultid="3414" />
                    <RANKING order="4" place="4" resultid="2914" />
                    <RANKING order="5" place="5" resultid="3406" />
                    <RANKING order="6" place="6" resultid="2978" />
                    <RANKING order="7" place="7" resultid="3322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2303" />
                    <RANKING order="2" place="2" resultid="2884" />
                    <RANKING order="3" place="3" resultid="2114" />
                    <RANKING order="4" place="4" resultid="2957" />
                    <RANKING order="5" place="5" resultid="3238" />
                    <RANKING order="6" place="6" resultid="3650" />
                    <RANKING order="7" place="7" resultid="2406" />
                    <RANKING order="8" place="-1" resultid="2397" />
                    <RANKING order="9" place="-1" resultid="2931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3091" />
                    <RANKING order="2" place="2" resultid="2963" />
                    <RANKING order="3" place="3" resultid="2463" />
                    <RANKING order="4" place="4" resultid="2498" />
                    <RANKING order="5" place="5" resultid="2261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2422" />
                    <RANKING order="2" place="2" resultid="3494" />
                    <RANKING order="3" place="3" resultid="3781" />
                    <RANKING order="4" place="-1" resultid="1891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2107" />
                    <RANKING order="2" place="2" resultid="2429" />
                    <RANKING order="3" place="3" resultid="2875" />
                    <RANKING order="4" place="4" resultid="3011" />
                    <RANKING order="5" place="5" resultid="3455" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2413" />
                    <RANKING order="2" place="2" resultid="3103" />
                    <RANKING order="3" place="3" resultid="1797" />
                    <RANKING order="4" place="4" resultid="3119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3712" />
                    <RANKING order="2" place="2" resultid="3904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2199" />
                    <RANKING order="2" place="2" resultid="3912" />
                    <RANKING order="3" place="3" resultid="3786" />
                    <RANKING order="4" place="4" resultid="3210" />
                    <RANKING order="5" place="5" resultid="1898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1072" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1073" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1074" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1075" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4596" daytime="14:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4597" daytime="14:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4598" daytime="14:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4599" daytime="14:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4600" daytime="14:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4601" daytime="14:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4602" daytime="14:10" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1090" daytime="14:10" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1091" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2938" />
                    <RANKING order="2" place="2" resultid="2657" />
                    <RANKING order="3" place="3" resultid="3746" />
                    <RANKING order="4" place="4" resultid="2681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3799" />
                    <RANKING order="2" place="2" resultid="3365" />
                    <RANKING order="3" place="3" resultid="2675" />
                    <RANKING order="4" place="4" resultid="3963" />
                    <RANKING order="5" place="5" resultid="2626" />
                    <RANKING order="6" place="6" resultid="3981" />
                    <RANKING order="7" place="7" resultid="2781" />
                    <RANKING order="8" place="8" resultid="2825" />
                    <RANKING order="9" place="9" resultid="3161" />
                    <RANKING order="10" place="10" resultid="3046" />
                    <RANKING order="11" place="11" resultid="2872" />
                    <RANKING order="12" place="12" resultid="3972" />
                    <RANKING order="13" place="13" resultid="2638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2709" />
                    <RANKING order="2" place="2" resultid="3766" />
                    <RANKING order="3" place="3" resultid="3065" />
                    <RANKING order="4" place="4" resultid="3816" />
                    <RANKING order="5" place="5" resultid="3354" />
                    <RANKING order="6" place="6" resultid="3042" />
                    <RANKING order="7" place="7" resultid="2807" />
                    <RANKING order="8" place="8" resultid="3430" />
                    <RANKING order="9" place="9" resultid="2688" />
                    <RANKING order="10" place="10" resultid="1989" />
                    <RANKING order="11" place="11" resultid="3291" />
                    <RANKING order="12" place="12" resultid="2549" />
                    <RANKING order="13" place="13" resultid="2345" />
                    <RANKING order="14" place="14" resultid="2755" />
                    <RANKING order="15" place="15" resultid="3601" />
                    <RANKING order="16" place="-1" resultid="2354" />
                    <RANKING order="17" place="-1" resultid="2838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2727" />
                    <RANKING order="2" place="2" resultid="2722" />
                    <RANKING order="3" place="3" resultid="2974" />
                    <RANKING order="4" place="4" resultid="3894" />
                    <RANKING order="5" place="5" resultid="3388" />
                    <RANKING order="6" place="6" resultid="2787" />
                    <RANKING order="7" place="7" resultid="1812" />
                    <RANKING order="8" place="8" resultid="3005" />
                    <RANKING order="9" place="9" resultid="2929" />
                    <RANKING order="10" place="10" resultid="2671" />
                    <RANKING order="11" place="11" resultid="2217" />
                    <RANKING order="12" place="12" resultid="2701" />
                    <RANKING order="13" place="13" resultid="2981" />
                    <RANKING order="14" place="14" resultid="2520" />
                    <RANKING order="15" place="15" resultid="2666" />
                    <RANKING order="16" place="-1" resultid="2955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3485" />
                    <RANKING order="2" place="2" resultid="2917" />
                    <RANKING order="3" place="3" resultid="3803" />
                    <RANKING order="4" place="4" resultid="3146" />
                    <RANKING order="5" place="5" resultid="3809" />
                    <RANKING order="6" place="6" resultid="4020" />
                    <RANKING order="7" place="7" resultid="1852" />
                    <RANKING order="8" place="8" resultid="2545" />
                    <RANKING order="9" place="9" resultid="2758" />
                    <RANKING order="10" place="10" resultid="2922" />
                    <RANKING order="11" place="11" resultid="4003" />
                    <RANKING order="12" place="12" resultid="2694" />
                    <RANKING order="13" place="13" resultid="2765" />
                    <RANKING order="14" place="-1" resultid="3837" />
                    <RANKING order="15" place="-1" resultid="3166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3350" />
                    <RANKING order="2" place="2" resultid="3656" />
                    <RANKING order="3" place="3" resultid="3247" />
                    <RANKING order="4" place="4" resultid="1845" />
                    <RANKING order="5" place="5" resultid="2770" />
                    <RANKING order="6" place="6" resultid="2300" />
                    <RANKING order="7" place="7" resultid="1873" />
                    <RANKING order="8" place="8" resultid="3664" />
                    <RANKING order="9" place="9" resultid="3019" />
                    <RANKING order="10" place="10" resultid="3194" />
                    <RANKING order="11" place="11" resultid="2965" />
                    <RANKING order="12" place="12" resultid="2011" />
                    <RANKING order="13" place="13" resultid="2846" />
                    <RANKING order="14" place="14" resultid="3478" />
                    <RANKING order="15" place="15" resultid="2472" />
                    <RANKING order="16" place="16" resultid="2738" />
                    <RANKING order="17" place="17" resultid="2925" />
                    <RANKING order="18" place="18" resultid="2763" />
                    <RANKING order="19" place="19" resultid="2761" />
                    <RANKING order="20" place="20" resultid="2248" />
                    <RANKING order="21" place="21" resultid="3678" />
                    <RANKING order="22" place="-1" resultid="3673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3760" />
                    <RANKING order="2" place="2" resultid="2794" />
                    <RANKING order="3" place="3" resultid="2851" />
                    <RANKING order="4" place="4" resultid="3751" />
                    <RANKING order="5" place="5" resultid="3917" />
                    <RANKING order="6" place="6" resultid="2242" />
                    <RANKING order="7" place="7" resultid="3054" />
                    <RANKING order="8" place="-1" resultid="1816" />
                    <RANKING order="9" place="-1" resultid="3469" />
                    <RANKING order="10" place="-1" resultid="3875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3185" />
                    <RANKING order="2" place="2" resultid="3447" />
                    <RANKING order="3" place="3" resultid="3792" />
                    <RANKING order="4" place="4" resultid="3622" />
                    <RANKING order="5" place="5" resultid="3050" />
                    <RANKING order="6" place="6" resultid="3438" />
                    <RANKING order="7" place="7" resultid="1937" />
                    <RANKING order="8" place="8" resultid="1966" />
                    <RANKING order="9" place="9" resultid="2997" />
                    <RANKING order="10" place="10" resultid="2968" />
                    <RANKING order="11" place="11" resultid="3498" />
                    <RANKING order="12" place="12" resultid="1945" />
                    <RANKING order="13" place="13" resultid="3201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3261" />
                    <RANKING order="2" place="2" resultid="1785" />
                    <RANKING order="3" place="3" resultid="2290" />
                    <RANKING order="4" place="4" resultid="1963" />
                    <RANKING order="5" place="5" resultid="3032" />
                    <RANKING order="6" place="6" resultid="2442" />
                    <RANKING order="7" place="7" resultid="2732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2210" />
                    <RANKING order="2" place="2" resultid="2363" />
                    <RANKING order="3" place="3" resultid="2801" />
                    <RANKING order="4" place="4" resultid="1802" />
                    <RANKING order="5" place="5" resultid="2489" />
                    <RANKING order="6" place="6" resultid="2155" />
                    <RANKING order="7" place="7" resultid="1882" />
                    <RANKING order="8" place="8" resultid="2609" />
                    <RANKING order="9" place="9" resultid="3926" />
                    <RANKING order="10" place="10" resultid="3452" />
                    <RANKING order="11" place="11" resultid="3219" />
                    <RANKING order="12" place="12" resultid="2123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3296" />
                    <RANKING order="2" place="2" resultid="2282" />
                    <RANKING order="3" place="3" resultid="3867" />
                    <RANKING order="4" place="4" resultid="2456" />
                    <RANKING order="5" place="5" resultid="2864" />
                    <RANKING order="6" place="6" resultid="3721" />
                    <RANKING order="7" place="7" resultid="2103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2016" />
                    <RANKING order="2" place="2" resultid="2205" />
                    <RANKING order="3" place="3" resultid="3853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2137" />
                    <RANKING order="2" place="2" resultid="2192" />
                    <RANKING order="3" place="3" resultid="3613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1105" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1106" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4603" daytime="14:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4604" daytime="14:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4605" daytime="14:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4606" daytime="14:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4607" daytime="14:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4608" daytime="14:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4609" daytime="14:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4610" daytime="14:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4611" daytime="14:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4612" daytime="14:25" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4613" daytime="14:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4614" daytime="14:30" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4615" daytime="14:30" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4616" daytime="14:35" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="4617" daytime="14:35" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="14:35" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2645" />
                    <RANKING order="2" place="2" resultid="3635" />
                    <RANKING order="3" place="3" resultid="3085" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3740" />
                    <RANKING order="2" place="2" resultid="3823" />
                    <RANKING order="3" place="3" resultid="3957" />
                    <RANKING order="4" place="4" resultid="3379" />
                    <RANKING order="5" place="5" resultid="1823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2166" />
                    <RANKING order="2" place="2" resultid="3590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3342" />
                    <RANKING order="2" place="2" resultid="3154" />
                    <RANKING order="3" place="3" resultid="3140" />
                    <RANKING order="4" place="4" resultid="3993" />
                    <RANKING order="5" place="-1" resultid="3323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2304" />
                    <RANKING order="2" place="2" resultid="2115" />
                    <RANKING order="3" place="3" resultid="2398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2330" />
                    <RANKING order="2" place="2" resultid="2529" />
                    <RANKING order="3" place="3" resultid="3934" />
                    <RANKING order="4" place="4" resultid="2480" />
                    <RANKING order="5" place="5" resultid="2464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2423" />
                    <RANKING order="2" place="2" resultid="3369" />
                    <RANKING order="3" place="3" resultid="2511" />
                    <RANKING order="4" place="4" resultid="2273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2108" />
                    <RANKING order="2" place="2" resultid="3012" />
                    <RANKING order="3" place="3" resultid="3077" />
                    <RANKING order="4" place="4" resultid="2746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2414" />
                    <RANKING order="2" place="2" resultid="2591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat" />
                <AGEGROUP agegroupid="1119" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1120" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1121" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1122" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1123" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4618" daytime="14:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4619" daytime="14:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4620" daytime="14:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4621" daytime="14:50" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="14:55" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2658" />
                    <RANKING order="2" place="2" resultid="3628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2812" />
                    <RANKING order="2" place="2" resultid="2826" />
                    <RANKING order="3" place="3" resultid="3646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3316" />
                    <RANKING order="2" place="2" resultid="2355" />
                    <RANKING order="3" place="3" resultid="2712" />
                    <RANKING order="4" place="4" resultid="3431" />
                    <RANKING order="5" place="5" resultid="1994" />
                    <RANKING order="6" place="6" resultid="2346" />
                    <RANKING order="7" place="7" resultid="3602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2728" />
                    <RANKING order="2" place="2" resultid="3895" />
                    <RANKING order="3" place="3" resultid="1933" />
                    <RANKING order="4" place="4" resultid="2236" />
                    <RANKING order="5" place="5" resultid="2982" />
                    <RANKING order="6" place="-1" resultid="2521" />
                    <RANKING order="7" place="-1" resultid="3687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3486" />
                    <RANKING order="2" place="2" resultid="2174" />
                    <RANKING order="3" place="3" resultid="3147" />
                    <RANKING order="4" place="-1" resultid="3167" />
                    <RANKING order="5" place="-1" resultid="3399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3195" />
                    <RANKING order="2" place="2" resultid="1874" />
                    <RANKING order="3" place="3" resultid="3335" />
                    <RANKING order="4" place="4" resultid="2299" />
                    <RANKING order="5" place="5" resultid="3393" />
                    <RANKING order="6" place="6" resultid="2473" />
                    <RANKING order="7" place="-1" resultid="2935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3025" />
                    <RANKING order="2" place="2" resultid="2852" />
                    <RANKING order="3" place="3" resultid="2264" />
                    <RANKING order="4" place="4" resultid="3876" />
                    <RANKING order="5" place="5" resultid="1927" />
                    <RANKING order="6" place="-1" resultid="2600" />
                    <RANKING order="7" place="-1" resultid="3470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1132" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3186" />
                    <RANKING order="2" place="2" resultid="3202" />
                    <RANKING order="3" place="3" resultid="1922" />
                    <RANKING order="4" place="4" resultid="1946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1133" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1786" />
                    <RANKING order="2" place="2" resultid="3033" />
                    <RANKING order="3" place="3" resultid="3357" />
                    <RANKING order="4" place="4" resultid="2733" />
                    <RANKING order="5" place="-1" resultid="2443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2211" />
                    <RANKING order="2" place="2" resultid="2156" />
                    <RANKING order="3" place="3" resultid="2490" />
                    <RANKING order="4" place="4" resultid="3998" />
                    <RANKING order="5" place="5" resultid="1978" />
                    <RANKING order="6" place="-1" resultid="2388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3297" />
                    <RANKING order="2" place="2" resultid="3281" />
                    <RANKING order="3" place="3" resultid="1859" />
                    <RANKING order="4" place="4" resultid="2457" />
                    <RANKING order="5" place="-1" resultid="2023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1912" />
                    <RANKING order="2" place="2" resultid="1981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1139" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1140" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4622" daytime="14:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4623" daytime="15:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4624" daytime="15:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4625" daytime="15:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4626" daytime="15:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4627" daytime="15:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4628" daytime="15:25" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1141" daytime="15:30" gender="X" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1142" agemax="-1" agemin="-1" name="&quot;0&quot; 0-99 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="119" agemin="100" name="&quot;A&quot; 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3505" />
                    <RANKING order="2" place="2" resultid="4037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="159" agemin="120" name="&quot;B&quot; 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4409" />
                    <RANKING order="2" place="2" resultid="3301" />
                    <RANKING order="3" place="3" resultid="3507" />
                    <RANKING order="4" place="4" resultid="3117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="199" agemin="160" name="&quot;C&quot; 160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3509" />
                    <RANKING order="2" place="2" resultid="3302" />
                    <RANKING order="3" place="3" resultid="2945" />
                    <RANKING order="4" place="4" resultid="3513" />
                    <RANKING order="5" place="5" resultid="2555" />
                    <RANKING order="6" place="-1" resultid="2990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="239" agemin="200" name="&quot;D&quot; 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3511" />
                    <RANKING order="2" place="2" resultid="2553" />
                    <RANKING order="3" place="3" resultid="3112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="279" agemin="240" name="&quot;E&quot; 240-279 lat " calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="-1" agemin="280" name="&quot;F&quot; 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4629" daytime="15:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4630" daytime="15:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1158" daytime="15:35" gender="F" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1166" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3086" />
                    <RANKING order="2" place="-1" resultid="3098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3948" />
                    <RANKING order="2" place="2" resultid="3824" />
                    <RANKING order="3" place="-1" resultid="3772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3695" />
                    <RANKING order="2" place="2" resultid="3233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3141" />
                    <RANKING order="2" place="2" resultid="3994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3239" />
                    <RANKING order="2" place="-1" resultid="2958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2331" />
                    <RANKING order="2" place="2" resultid="3092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1892" />
                    <RANKING order="2" place="2" resultid="2512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2592" />
                    <RANKING order="2" place="2" resultid="3104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat" />
                <AGEGROUP agegroupid="1176" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat" />
                <AGEGROUP agegroupid="1177" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1178" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1179" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1180" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1181" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4631" daytime="15:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4632" daytime="15:50" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1182" daytime="16:05" gender="M" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1183" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3964" />
                    <RANKING order="2" place="2" resultid="2823" />
                    <RANKING order="3" place="-1" resultid="3982" />
                    <RANKING order="4" place="-1" resultid="3973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2356" />
                    <RANKING order="2" place="2" resultid="2689" />
                    <RANKING order="3" place="3" resultid="1940" />
                    <RANKING order="4" place="4" resultid="1995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1813" />
                    <RANKING order="2" place="-1" resultid="3058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2175" />
                    <RANKING order="2" place="2" resultid="3810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3657" />
                    <RANKING order="2" place="2" resultid="1846" />
                    <RANKING order="3" place="3" resultid="2669" />
                    <RANKING order="4" place="4" resultid="2739" />
                    <RANKING order="5" place="5" resultid="2847" />
                    <RANKING order="6" place="-1" resultid="3679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3701" />
                    <RANKING order="2" place="2" resultid="2601" />
                    <RANKING order="3" place="3" resultid="3918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3623" />
                    <RANKING order="2" place="2" resultid="3439" />
                    <RANKING order="3" place="3" resultid="1967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3262" />
                    <RANKING order="2" place="2" resultid="3358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2389" />
                    <RANKING order="2" place="2" resultid="1883" />
                    <RANKING order="3" place="3" resultid="1803" />
                    <RANKING order="4" place="4" resultid="3999" />
                    <RANKING order="5" place="5" resultid="3220" />
                    <RANKING order="6" place="6" resultid="3453" />
                    <RANKING order="7" place="7" resultid="1979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3868" />
                    <RANKING order="2" place="2" resultid="2283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1913" />
                    <RANKING order="2" place="-1" resultid="3854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2138" />
                    <RANKING order="2" place="-1" resultid="3614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1197" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1198" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4633" daytime="16:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4634" daytime="16:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4635" daytime="16:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4636" daytime="16:55" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1199" daytime="17:10" gender="F" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1200" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat" />
                <AGEGROUP agegroupid="1201" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat" />
                <AGEGROUP agegroupid="1202" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat" />
                <AGEGROUP agegroupid="1203" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat" />
                <AGEGROUP agegroupid="1204" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat" />
                <AGEGROUP agegroupid="1210" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1212" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1213" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1214" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1215" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4637" daytime="17:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1216" daytime="17:45" gender="M" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1217" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat" />
                <AGEGROUP agegroupid="1218" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat" />
                <AGEGROUP agegroupid="1219" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat" />
                <AGEGROUP agegroupid="1221" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3665" />
                    <RANKING order="2" place="2" resultid="1835" />
                    <RANKING order="3" place="3" resultid="3226" />
                    <RANKING order="4" place="-1" resultid="2936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2795" />
                    <RANKING order="2" place="2" resultid="2265" />
                    <RANKING order="3" place="3" resultid="3752" />
                    <RANKING order="4" place="4" resultid="2434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1938" />
                    <RANKING order="2" place="-1" resultid="2184" />
                    <RANKING order="3" place="-1" resultid="1923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2451" />
                    <RANKING order="2" place="2" resultid="1839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3730" />
                    <RANKING order="2" place="2" resultid="2610" />
                    <RANKING order="3" place="-1" resultid="2383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2024" />
                    <RANKING order="2" place="2" resultid="3939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1229" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1230" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1231" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1232" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4638" daytime="17:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4639" daytime="18:15" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2023-06-03" daytime="09:00" endtime="11:35" name="II BLOK" number="2" officialmeeting="08:55" warmupfrom="08:15">
          <EVENTS>
            <EVENT eventid="1234" daytime="09:00" gender="F" number="10" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1236" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2908" />
                    <RANKING order="2" place="2" resultid="4009" />
                    <RANKING order="3" place="3" resultid="2646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3773" />
                    <RANKING order="2" place="2" resultid="3255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3591" />
                    <RANKING order="2" place="2" resultid="3181" />
                    <RANKING order="3" place="3" resultid="3460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3343" />
                    <RANKING order="2" place="2" resultid="2631" />
                    <RANKING order="3" place="3" resultid="3324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2920" />
                    <RANKING order="2" place="2" resultid="2305" />
                    <RANKING order="3" place="3" resultid="2116" />
                    <RANKING order="4" place="4" resultid="2368" />
                    <RANKING order="5" place="5" resultid="3651" />
                    <RANKING order="6" place="6" resultid="2620" />
                    <RANKING order="7" place="7" resultid="2985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2233" />
                    <RANKING order="2" place="2" resultid="2465" />
                    <RANKING order="3" place="3" resultid="2499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2424" />
                    <RANKING order="2" place="2" resultid="1905" />
                    <RANKING order="3" place="3" resultid="2513" />
                    <RANKING order="4" place="4" resultid="3495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2109" />
                    <RANKING order="2" place="2" resultid="2430" />
                    <RANKING order="3" place="3" resultid="2876" />
                    <RANKING order="4" place="4" resultid="3456" />
                    <RANKING order="5" place="5" resultid="2748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2415" />
                    <RANKING order="2" place="2" resultid="2593" />
                    <RANKING order="3" place="3" resultid="3105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3714" />
                    <RANKING order="2" place="2" resultid="3905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3913" />
                    <RANKING order="2" place="2" resultid="1899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1248" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1249" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1250" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1251" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4640" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4641" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4642" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4643" daytime="09:05" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1252" daytime="09:10" gender="M" number="11" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1253" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2659" />
                    <RANKING order="2" place="2" resultid="2682" />
                    <RANKING order="3" place="3" resultid="3630" />
                    <RANKING order="4" place="-1" resultid="1956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2676" />
                    <RANKING order="2" place="2" resultid="3384" />
                    <RANKING order="3" place="3" resultid="3366" />
                    <RANKING order="4" place="4" resultid="3848" />
                    <RANKING order="5" place="5" resultid="2782" />
                    <RANKING order="6" place="6" resultid="2775" />
                    <RANKING order="7" place="7" resultid="3983" />
                    <RANKING order="8" place="8" resultid="2639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3355" />
                    <RANKING order="2" place="2" resultid="3432" />
                    <RANKING order="3" place="3" resultid="2347" />
                    <RANKING order="4" place="4" resultid="1941" />
                    <RANKING order="5" place="-1" resultid="1996" />
                    <RANKING order="6" place="-1" resultid="2839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2723" />
                    <RANKING order="2" place="2" resultid="3269" />
                    <RANKING order="3" place="3" resultid="3006" />
                    <RANKING order="4" place="4" resultid="2522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3487" />
                    <RANKING order="2" place="2" resultid="3168" />
                    <RANKING order="3" place="2" resultid="3400" />
                    <RANKING order="4" place="4" resultid="3838" />
                    <RANKING order="5" place="-1" resultid="4013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3351" />
                    <RANKING order="2" place="2" resultid="3020" />
                    <RANKING order="3" place="3" resultid="3336" />
                    <RANKING order="4" place="4" resultid="2771" />
                    <RANKING order="5" place="5" resultid="3666" />
                    <RANKING order="6" place="6" resultid="2538" />
                    <RANKING order="7" place="7" resultid="2012" />
                    <RANKING order="8" place="8" resultid="2240" />
                    <RANKING order="9" place="9" resultid="2316" />
                    <RANKING order="10" place="10" resultid="2474" />
                    <RANKING order="11" place="-1" resultid="3680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3753" />
                    <RANKING order="2" place="2" resultid="2602" />
                    <RANKING order="3" place="3" resultid="3919" />
                    <RANKING order="4" place="4" resultid="3844" />
                    <RANKING order="5" place="-1" resultid="1817" />
                    <RANKING order="6" place="-1" resultid="3471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3793" />
                    <RANKING order="2" place="2" resultid="3187" />
                    <RANKING order="3" place="3" resultid="1968" />
                    <RANKING order="4" place="4" resultid="2185" />
                    <RANKING order="5" place="5" resultid="2969" />
                    <RANKING order="6" place="6" resultid="3203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat" />
                <AGEGROUP agegroupid="1262" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2212" />
                    <RANKING order="2" place="2" resultid="2802" />
                    <RANKING order="3" place="3" resultid="2491" />
                    <RANKING order="4" place="4" resultid="1884" />
                    <RANKING order="5" place="5" resultid="3927" />
                    <RANKING order="6" place="6" resultid="2124" />
                    <RANKING order="7" place="-1" resultid="1804" />
                    <RANKING order="8" place="-1" resultid="2390" />
                    <RANKING order="9" place="-1" resultid="3221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2025" />
                    <RANKING order="2" place="2" resultid="3869" />
                    <RANKING order="3" place="3" resultid="3940" />
                    <RANKING order="4" place="4" resultid="4805" />
                    <RANKING order="5" place="5" resultid="3722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2017" />
                    <RANKING order="2" place="2" resultid="1914" />
                    <RANKING order="3" place="3" resultid="3855" />
                    <RANKING order="4" place="4" resultid="2206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4016" />
                    <RANKING order="2" place="2" resultid="2193" />
                    <RANKING order="3" place="3" resultid="3615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1267" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1268" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4644" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4645" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4646" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4647" daytime="09:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4648" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4649" daytime="09:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4650" daytime="09:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4651" daytime="09:25" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1269" daytime="09:25" gender="F" number="12" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1270" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3087" />
                    <RANKING order="2" place="2" resultid="3636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3825" />
                    <RANKING order="2" place="2" resultid="3380" />
                    <RANKING order="3" place="3" resultid="1824" />
                    <RANKING order="4" place="-1" resultid="3774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2167" />
                    <RANKING order="2" place="2" resultid="3176" />
                    <RANKING order="3" place="3" resultid="3331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2613" />
                    <RANKING order="2" place="2" resultid="3407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2621" />
                    <RANKING order="2" place="2" resultid="2399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2332" />
                    <RANKING order="2" place="2" resultid="3935" />
                    <RANKING order="3" place="3" resultid="2466" />
                    <RANKING order="4" place="4" resultid="2482" />
                    <RANKING order="5" place="-1" resultid="2339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1893" />
                    <RANKING order="2" place="2" resultid="3371" />
                    <RANKING order="3" place="3" resultid="3782" />
                    <RANKING order="4" place="4" resultid="2274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3013" />
                    <RANKING order="2" place="2" resultid="3079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1282" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1283" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1284" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1285" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4652" daytime="09:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4653" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4654" daytime="09:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="09:40" gender="M" number="13" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1287" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3631" />
                    <RANKING order="2" place="2" resultid="1957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2813" />
                    <RANKING order="2" place="2" resultid="3974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3317" />
                    <RANKING order="2" place="2" resultid="2653" />
                    <RANKING order="3" place="3" resultid="2713" />
                    <RANKING order="4" place="4" resultid="3603" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3148" />
                    <RANKING order="2" place="2" resultid="2176" />
                    <RANKING order="3" place="3" resultid="2320" />
                    <RANKING order="4" place="-1" resultid="2004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3196" />
                    <RANKING order="2" place="2" resultid="2539" />
                    <RANKING order="3" place="3" resultid="3674" />
                    <RANKING order="4" place="-1" resultid="1830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3861" />
                    <RANKING order="2" place="2" resultid="2266" />
                    <RANKING order="3" place="3" resultid="2435" />
                    <RANKING order="4" place="-1" resultid="3472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3448" />
                    <RANKING order="2" place="2" resultid="3440" />
                    <RANKING order="3" place="3" resultid="2504" />
                    <RANKING order="4" place="4" resultid="3499" />
                    <RANKING order="5" place="5" resultid="1947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2359" />
                    <RANKING order="2" place="2" resultid="2130" />
                    <RANKING order="3" place="3" resultid="2444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2157" />
                    <RANKING order="2" place="2" resultid="2492" />
                    <RANKING order="3" place="3" resultid="3731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3282" />
                    <RANKING order="2" place="2" resultid="1860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1298" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2377" />
                    <RANKING order="2" place="2" resultid="1982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1299" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1300" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1301" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1302" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4655" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4656" daytime="09:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4657" daytime="09:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4658" daytime="10:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1303" daytime="10:05" gender="F" number="14" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1304" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4010" />
                    <RANKING order="2" place="2" resultid="2647" />
                    <RANKING order="3" place="3" resultid="3640" />
                    <RANKING order="4" place="4" resultid="3099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3424" />
                    <RANKING order="2" place="2" resultid="3958" />
                    <RANKING order="3" place="3" resultid="3741" />
                    <RANKING order="4" place="4" resultid="3256" />
                    <RANKING order="5" place="5" resultid="3949" />
                    <RANKING order="6" place="6" resultid="3826" />
                    <RANKING order="7" place="7" resultid="1825" />
                    <RANKING order="8" place="8" resultid="3069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2168" />
                    <RANKING order="2" place="2" resultid="3234" />
                    <RANKING order="3" place="3" resultid="3461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3344" />
                    <RANKING order="2" place="2" resultid="2632" />
                    <RANKING order="3" place="3" resultid="2614" />
                    <RANKING order="4" place="4" resultid="3415" />
                    <RANKING order="5" place="5" resultid="3408" />
                    <RANKING order="6" place="6" resultid="2979" />
                    <RANKING order="7" place="7" resultid="3325" />
                    <RANKING order="8" place="8" resultid="3610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2306" />
                    <RANKING order="2" place="2" resultid="2885" />
                    <RANKING order="3" place="3" resultid="2117" />
                    <RANKING order="4" place="4" resultid="3240" />
                    <RANKING order="5" place="5" resultid="2369" />
                    <RANKING order="6" place="6" resultid="2407" />
                    <RANKING order="7" place="-1" resultid="2400" />
                    <RANKING order="8" place="-1" resultid="2622" />
                    <RANKING order="9" place="-1" resultid="2959" />
                    <RANKING order="10" place="-1" resultid="3652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3093" />
                    <RANKING order="2" place="2" resultid="2500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3372" />
                    <RANKING order="2" place="2" resultid="2275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2110" />
                    <RANKING order="2" place="2" resultid="2431" />
                    <RANKING order="3" place="3" resultid="2877" />
                    <RANKING order="4" place="4" resultid="2749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2416" />
                    <RANKING order="2" place="2" resultid="1798" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3914" />
                    <RANKING order="2" place="2" resultid="3787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1316" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1317" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1318" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1319" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4659" daytime="10:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4660" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4661" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4662" daytime="10:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4663" daytime="10:15" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1320" daytime="10:15" gender="M" number="15" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1321" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2939" />
                    <RANKING order="2" place="2" resultid="3747" />
                    <RANKING order="3" place="3" resultid="2660" />
                    <RANKING order="4" place="4" resultid="2683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1322" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2677" />
                    <RANKING order="2" place="2" resultid="2827" />
                    <RANKING order="3" place="3" resultid="2776" />
                    <RANKING order="4" place="4" resultid="3965" />
                    <RANKING order="5" place="5" resultid="3984" />
                    <RANKING order="6" place="6" resultid="2873" />
                    <RANKING order="7" place="7" resultid="3162" />
                    <RANKING order="8" place="8" resultid="3975" />
                    <RANKING order="9" place="9" resultid="2640" />
                    <RANKING order="10" place="10" resultid="1954" />
                    <RANKING order="11" place="11" resultid="3647" />
                    <RANKING order="12" place="-1" resultid="2783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1323" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2719" />
                    <RANKING order="2" place="2" resultid="2808" />
                    <RANKING order="3" place="3" resultid="3817" />
                    <RANKING order="4" place="4" resultid="2690" />
                    <RANKING order="5" place="5" resultid="2756" />
                    <RANKING order="6" place="6" resultid="3604" />
                    <RANKING order="7" place="-1" resultid="2348" />
                    <RANKING order="8" place="-1" resultid="2840" />
                    <RANKING order="9" place="-1" resultid="3043" />
                    <RANKING order="10" place="-1" resultid="3433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1324" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2729" />
                    <RANKING order="2" place="2" resultid="2724" />
                    <RANKING order="3" place="3" resultid="3896" />
                    <RANKING order="4" place="4" resultid="3389" />
                    <RANKING order="5" place="5" resultid="2788" />
                    <RANKING order="6" place="6" resultid="1934" />
                    <RANKING order="7" place="7" resultid="3270" />
                    <RANKING order="8" place="8" resultid="2237" />
                    <RANKING order="9" place="9" resultid="2704" />
                    <RANKING order="10" place="10" resultid="2672" />
                    <RANKING order="11" place="11" resultid="3059" />
                    <RANKING order="12" place="12" resultid="2218" />
                    <RANKING order="13" place="13" resultid="2702" />
                    <RANKING order="14" place="14" resultid="2667" />
                    <RANKING order="15" place="15" resultid="2523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1325" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3488" />
                    <RANKING order="2" place="2" resultid="2918" />
                    <RANKING order="3" place="3" resultid="3804" />
                    <RANKING order="4" place="4" resultid="2313" />
                    <RANKING order="5" place="5" resultid="4022" />
                    <RANKING order="6" place="6" resultid="3839" />
                    <RANKING order="7" place="7" resultid="3169" />
                    <RANKING order="8" place="8" resultid="2923" />
                    <RANKING order="9" place="9" resultid="2759" />
                    <RANKING order="10" place="10" resultid="2546" />
                    <RANKING order="11" place="11" resultid="2695" />
                    <RANKING order="12" place="12" resultid="4004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1326" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1847" />
                    <RANKING order="2" place="2" resultid="3248" />
                    <RANKING order="3" place="3" resultid="3227" />
                    <RANKING order="4" place="4" resultid="2298" />
                    <RANKING order="5" place="5" resultid="1875" />
                    <RANKING order="6" place="6" resultid="3667" />
                    <RANKING order="7" place="7" resultid="3420" />
                    <RANKING order="8" place="8" resultid="2013" />
                    <RANKING order="9" place="9" resultid="3479" />
                    <RANKING order="10" place="10" resultid="2475" />
                    <RANKING order="11" place="11" resultid="2740" />
                    <RANKING order="12" place="12" resultid="2926" />
                    <RANKING order="13" place="13" resultid="2988" />
                    <RANKING order="14" place="14" resultid="3681" />
                    <RANKING order="15" place="15" resultid="2249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3761" />
                    <RANKING order="2" place="2" resultid="2853" />
                    <RANKING order="3" place="3" resultid="2796" />
                    <RANKING order="4" place="4" resultid="3920" />
                    <RANKING order="5" place="5" resultid="2603" />
                    <RANKING order="6" place="6" resultid="2243" />
                    <RANKING order="7" place="7" resultid="3055" />
                    <RANKING order="8" place="-1" resultid="1818" />
                    <RANKING order="9" place="-1" resultid="3877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1328" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3188" />
                    <RANKING order="2" place="2" resultid="3624" />
                    <RANKING order="3" place="3" resultid="3051" />
                    <RANKING order="4" place="4" resultid="1969" />
                    <RANKING order="5" place="5" resultid="2998" />
                    <RANKING order="6" place="6" resultid="4044" />
                    <RANKING order="7" place="7" resultid="2970" />
                    <RANKING order="8" place="8" resultid="3204" />
                    <RANKING order="9" place="-1" resultid="3500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1329" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3263" />
                    <RANKING order="2" place="2" resultid="1787" />
                    <RANKING order="3" place="3" resultid="2294" />
                    <RANKING order="4" place="4" resultid="1964" />
                    <RANKING order="5" place="5" resultid="2452" />
                    <RANKING order="6" place="6" resultid="3359" />
                    <RANKING order="7" place="7" resultid="2734" />
                    <RANKING order="8" place="8" resultid="1840" />
                    <RANKING order="9" place="-1" resultid="2445" />
                    <RANKING order="10" place="-1" resultid="3034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1330" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2213" />
                    <RANKING order="2" place="2" resultid="2364" />
                    <RANKING order="3" place="3" resultid="1805" />
                    <RANKING order="4" place="4" resultid="1885" />
                    <RANKING order="5" place="5" resultid="3732" />
                    <RANKING order="6" place="6" resultid="3928" />
                    <RANKING order="7" place="7" resultid="2125" />
                    <RANKING order="8" place="-1" resultid="3222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1331" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3298" />
                    <RANKING order="2" place="2" resultid="3870" />
                    <RANKING order="3" place="3" resultid="2284" />
                    <RANKING order="4" place="4" resultid="2458" />
                    <RANKING order="5" place="5" resultid="2865" />
                    <RANKING order="6" place="6" resultid="3723" />
                    <RANKING order="7" place="7" resultid="2104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1332" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2018" />
                    <RANKING order="2" place="2" resultid="3856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1333" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2139" />
                    <RANKING order="2" place="2" resultid="3616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1334" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1335" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1336" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4664" daytime="10:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4665" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4666" daytime="10:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4667" daytime="10:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4668" daytime="10:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4669" daytime="10:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4670" daytime="10:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4671" daytime="10:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4672" daytime="10:35" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4673" daytime="10:40" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4674" daytime="10:40" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4675" daytime="10:45" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1337" daytime="10:45" gender="F" number="16" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1338" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat" />
                <AGEGROUP agegroupid="1339" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3959" />
                    <RANKING order="2" place="2" resultid="3950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1340" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1341" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1342" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2333" />
                    <RANKING order="2" place="2" resultid="2530" />
                    <RANKING order="3" place="3" resultid="2483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1906" />
                    <RANKING order="2" place="2" resultid="2514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat" />
                <AGEGROUP agegroupid="1346" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat" />
                <AGEGROUP agegroupid="1348" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat" />
                <AGEGROUP agegroupid="1349" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1350" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1351" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1352" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1353" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4676" daytime="10:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4677" daytime="10:50" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1354" daytime="10:55" gender="M" number="17" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1355" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1356" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3800" />
                    <RANKING order="2" place="2" resultid="3966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1357" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1997" />
                    <RANKING order="2" place="2" resultid="4041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1358" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3897" />
                    <RANKING order="2" place="2" resultid="3689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1359" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2177" />
                    <RANKING order="2" place="2" resultid="3811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1360" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3658" />
                    <RANKING order="2" place="2" resultid="1836" />
                    <RANKING order="3" place="3" resultid="3021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1361" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3026" />
                    <RANKING order="2" place="2" resultid="3702" />
                    <RANKING order="3" place="3" resultid="2854" />
                    <RANKING order="4" place="4" resultid="2267" />
                    <RANKING order="5" place="5" resultid="3878" />
                    <RANKING order="6" place="6" resultid="1928" />
                    <RANKING order="7" place="-1" resultid="2436" />
                    <RANKING order="8" place="-1" resultid="3754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1362" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3441" />
                    <RANKING order="2" place="2" resultid="2505" />
                    <RANKING order="3" place="3" resultid="1948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1363" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2131" />
                    <RANKING order="2" place="-1" resultid="3035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1364" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2391" />
                    <RANKING order="2" place="2" resultid="2158" />
                    <RANKING order="3" place="-1" resultid="2384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1365" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1366" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1915" />
                    <RANKING order="2" place="2" resultid="1983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1367" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1368" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1369" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1370" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4678" daytime="10:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4679" daytime="11:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4680" daytime="11:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4681" daytime="11:15" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1371" daytime="11:15" gender="F" number="18" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1388" agemax="-1" agemin="-1" name="&quot;0&quot; 0-99 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="1389" agemax="119" agemin="100" name="&quot;A&quot; 100-119 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="1390" agemax="159" agemin="120" name="&quot;B&quot; 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3521" />
                    <RANKING order="2" place="2" resultid="3303" />
                    <RANKING order="3" place="3" resultid="3304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="199" agemin="160" name="&quot;C&quot; 160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3523" />
                    <RANKING order="2" place="2" resultid="2556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1392" agemax="239" agemin="200" name="&quot;D&quot; 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2552" />
                    <RANKING order="2" place="2" resultid="3113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1393" agemax="279" agemin="240" name="&quot;E&quot; 240-279 lat " calculate="TOTAL" />
                <AGEGROUP agegroupid="1394" agemax="-1" agemin="280" name="&quot;F&quot; 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4682" daytime="11:15" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1395" daytime="11:20" gender="M" number="19" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1396" agemax="-1" agemin="-1" name="&quot;0&quot; 0-99 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="119" agemin="100" name="&quot;A&quot; 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3515" />
                    <RANKING order="2" place="2" resultid="4038" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="159" agemin="120" name="&quot;B&quot; 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4410" />
                    <RANKING order="2" place="2" resultid="3305" />
                    <RANKING order="3" place="-1" resultid="2804" />
                    <RANKING order="4" place="-1" resultid="2887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1399" agemax="199" agemin="160" name="&quot;C&quot; 160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3516" />
                    <RANKING order="2" place="2" resultid="3833" />
                    <RANKING order="3" place="3" resultid="2326" />
                    <RANKING order="4" place="4" resultid="3118" />
                    <RANKING order="5" place="5" resultid="2993" />
                    <RANKING order="6" place="6" resultid="2944" />
                    <RANKING order="7" place="7" resultid="2253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1400" agemax="239" agemin="200" name="&quot;D&quot; 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3518" />
                    <RANKING order="2" place="2" resultid="3520" />
                    <RANKING order="3" place="3" resultid="2560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1401" agemax="279" agemin="240" name="&quot;E&quot; 240-279 lat " calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2558" />
                    <RANKING order="2" place="2" resultid="2221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1402" agemax="-1" agemin="280" name="&quot;F&quot; 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4683" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4684" daytime="11:25" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2023-06-03" daytime="14:35" endtime="18:08" name="III BLOK" number="3" warmupfrom="13:30" warmupuntil="13:55">
          <EVENTS>
            <EVENT eventid="1404" daytime="14:35" gender="F" number="20" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1406" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1407" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3827" />
                    <RANKING order="2" place="2" resultid="3381" />
                    <RANKING order="3" place="3" resultid="1826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1408" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2256" />
                    <RANKING order="2" place="2" resultid="3177" />
                    <RANKING order="3" place="3" resultid="3592" />
                    <RANKING order="4" place="4" resultid="3332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1409" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3278" />
                    <RANKING order="2" place="2" resultid="2615" />
                    <RANKING order="3" place="3" resultid="2779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2932" />
                    <RANKING order="2" place="2" resultid="2401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2340" />
                    <RANKING order="2" place="2" resultid="2334" />
                    <RANKING order="3" place="3" resultid="2531" />
                    <RANKING order="4" place="4" resultid="3936" />
                    <RANKING order="5" place="5" resultid="3275" />
                    <RANKING order="6" place="6" resultid="2467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1412" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1894" />
                    <RANKING order="2" place="2" resultid="3373" />
                    <RANKING order="3" place="3" resultid="3783" />
                    <RANKING order="4" place="4" resultid="2276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2111" />
                    <RANKING order="2" place="2" resultid="3080" />
                    <RANKING order="3" place="3" resultid="3014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3107" />
                    <RANKING order="2" place="2" resultid="3120" />
                    <RANKING order="3" place="3" resultid="2033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1415" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3788" />
                    <RANKING order="2" place="2" resultid="2200" />
                    <RANKING order="3" place="3" resultid="1900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1417" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1418" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1419" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1420" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1421" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4685" daytime="14:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4686" daytime="14:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4687" daytime="14:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4688" daytime="14:45" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1422" daytime="14:45" gender="M" number="21" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1423" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1424" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2814" />
                    <RANKING order="2" place="2" resultid="3047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2654" />
                    <RANKING order="2" place="2" resultid="3767" />
                    <RANKING order="3" place="3" resultid="2714" />
                    <RANKING order="4" place="4" resultid="3292" />
                    <RANKING order="5" place="5" resultid="1942" />
                    <RANKING order="6" place="6" resultid="3605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2975" />
                    <RANKING order="2" place="2" resultid="3690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3149" />
                    <RANKING order="2" place="2" resultid="2321" />
                    <RANKING order="3" place="3" resultid="2696" />
                    <RANKING order="4" place="4" resultid="2324" />
                    <RANKING order="5" place="5" resultid="2006" />
                    <RANKING order="6" place="-1" resultid="4025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3249" />
                    <RANKING order="2" place="2" resultid="1876" />
                    <RANKING order="3" place="3" resultid="2540" />
                    <RANKING order="4" place="4" resultid="3675" />
                    <RANKING order="5" place="5" resultid="2250" />
                    <RANKING order="6" place="6" resultid="1831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3862" />
                    <RANKING order="2" place="2" resultid="2437" />
                    <RANKING order="3" place="3" resultid="3056" />
                    <RANKING order="4" place="-1" resultid="3473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3449" />
                    <RANKING order="2" place="2" resultid="3501" />
                    <RANKING order="3" place="3" resultid="2999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1431" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3264" />
                    <RANKING order="2" place="2" resultid="2360" />
                    <RANKING order="3" place="3" resultid="2132" />
                    <RANKING order="4" place="4" resultid="2446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1432" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2159" />
                    <RANKING order="2" place="2" resultid="2126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3283" />
                    <RANKING order="2" place="2" resultid="1861" />
                    <RANKING order="3" place="3" resultid="2866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1435" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2195" />
                    <RANKING order="2" place="2" resultid="2140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1436" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1437" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1438" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4689" daytime="14:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4690" daytime="14:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4691" daytime="14:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4692" daytime="14:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4693" daytime="15:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1439" daytime="15:00" gender="F" number="22" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1440" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4011" />
                    <RANKING order="2" place="2" resultid="2648" />
                    <RANKING order="3" place="3" resultid="3638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1441" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3742" />
                    <RANKING order="2" place="2" resultid="3425" />
                    <RANKING order="3" place="3" resultid="2744" />
                    <RANKING order="4" place="4" resultid="3960" />
                    <RANKING order="5" place="5" resultid="3257" />
                    <RANKING order="6" place="6" resultid="3951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3587" />
                    <RANKING order="2" place="2" resultid="3584" />
                    <RANKING order="3" place="3" resultid="2257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3467" />
                    <RANKING order="2" place="2" resultid="2616" />
                    <RANKING order="3" place="3" resultid="3416" />
                    <RANKING order="4" place="4" resultid="3156" />
                    <RANKING order="5" place="5" resultid="3215" />
                    <RANKING order="6" place="6" resultid="3142" />
                    <RANKING order="7" place="7" resultid="3326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2307" />
                    <RANKING order="2" place="2" resultid="2886" />
                    <RANKING order="3" place="3" resultid="2118" />
                    <RANKING order="4" place="4" resultid="3242" />
                    <RANKING order="5" place="5" resultid="2960" />
                    <RANKING order="6" place="6" resultid="2408" />
                    <RANKING order="7" place="7" resultid="2402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2425" />
                    <RANKING order="2" place="2" resultid="2515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3015" />
                    <RANKING order="2" place="2" resultid="3081" />
                    <RANKING order="3" place="3" resultid="2750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1451" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1452" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1453" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1454" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1455" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4694" daytime="15:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4695" daytime="15:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4696" daytime="15:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4697" daytime="15:05" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1456" daytime="15:10" gender="M" number="23" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1457" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2661" />
                    <RANKING order="2" place="2" resultid="2940" />
                    <RANKING order="3" place="3" resultid="2684" />
                    <RANKING order="4" place="4" resultid="1959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1458" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2832" />
                    <RANKING order="2" place="2" resultid="3967" />
                    <RANKING order="3" place="3" resultid="2784" />
                    <RANKING order="4" place="4" resultid="2777" />
                    <RANKING order="5" place="5" resultid="3985" />
                    <RANKING order="6" place="6" resultid="3163" />
                    <RANKING order="7" place="7" resultid="3976" />
                    <RANKING order="8" place="8" resultid="3648" />
                    <RANKING order="9" place="-1" resultid="3367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2710" />
                    <RANKING order="2" place="2" resultid="2809" />
                    <RANKING order="3" place="3" resultid="3818" />
                    <RANKING order="4" place="4" resultid="3066" />
                    <RANKING order="5" place="5" resultid="3434" />
                    <RANKING order="6" place="6" resultid="2841" />
                    <RANKING order="7" place="7" resultid="3044" />
                    <RANKING order="8" place="8" resultid="1998" />
                    <RANKING order="9" place="9" resultid="2349" />
                    <RANKING order="10" place="10" resultid="3293" />
                    <RANKING order="11" place="-1" resultid="1990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1460" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2730" />
                    <RANKING order="2" place="2" resultid="3340" />
                    <RANKING order="3" place="3" resultid="3898" />
                    <RANKING order="4" place="4" resultid="2789" />
                    <RANKING order="5" place="5" resultid="1935" />
                    <RANKING order="6" place="6" resultid="3007" />
                    <RANKING order="7" place="7" resultid="2219" />
                    <RANKING order="8" place="8" resultid="2983" />
                    <RANKING order="9" place="9" resultid="3060" />
                    <RANKING order="10" place="10" resultid="2524" />
                    <RANKING order="11" place="-1" resultid="2238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1461" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3489" />
                    <RANKING order="2" place="2" resultid="3805" />
                    <RANKING order="3" place="3" resultid="2882" />
                    <RANKING order="4" place="4" resultid="3150" />
                    <RANKING order="5" place="5" resultid="3170" />
                    <RANKING order="6" place="6" resultid="3643" />
                    <RANKING order="7" place="7" resultid="2547" />
                    <RANKING order="8" place="8" resultid="1853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1462" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3352" />
                    <RANKING order="2" place="2" resultid="3659" />
                    <RANKING order="3" place="3" resultid="1848" />
                    <RANKING order="4" place="4" resultid="3250" />
                    <RANKING order="5" place="5" resultid="3228" />
                    <RANKING order="6" place="6" resultid="3832" />
                    <RANKING order="7" place="7" resultid="3480" />
                    <RANKING order="8" place="8" resultid="2476" />
                    <RANKING order="9" place="-1" resultid="2251" />
                    <RANKING order="10" place="-1" resultid="2966" />
                    <RANKING order="11" place="-1" resultid="3682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1463" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3027" />
                    <RANKING order="2" place="2" resultid="3762" />
                    <RANKING order="3" place="3" resultid="2855" />
                    <RANKING order="4" place="4" resultid="3755" />
                    <RANKING order="5" place="5" resultid="2797" />
                    <RANKING order="6" place="6" resultid="2244" />
                    <RANKING order="7" place="7" resultid="1929" />
                    <RANKING order="8" place="-1" resultid="2861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1464" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3189" />
                    <RANKING order="2" place="2" resultid="3052" />
                    <RANKING order="3" place="3" resultid="2506" />
                    <RANKING order="4" place="4" resultid="3205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1788" />
                    <RANKING order="2" place="2" resultid="2293" />
                    <RANKING order="3" place="3" resultid="2447" />
                    <RANKING order="4" place="4" resultid="2735" />
                    <RANKING order="5" place="5" resultid="3287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1466" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2214" />
                    <RANKING order="2" place="2" resultid="2365" />
                    <RANKING order="3" place="-1" resultid="2392" />
                    <RANKING order="4" place="-1" resultid="2493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2285" />
                    <RANKING order="2" place="2" resultid="1862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1468" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2019" />
                    <RANKING order="2" place="2" resultid="2207" />
                    <RANKING order="3" place="3" resultid="1984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1469" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1470" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1471" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1472" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4698" daytime="15:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4699" daytime="15:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4700" daytime="15:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4701" daytime="15:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4702" daytime="15:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4703" daytime="15:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4704" daytime="15:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4705" daytime="15:20" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1473" daytime="15:20" gender="F" number="24" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1474" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2909" />
                    <RANKING order="2" place="2" resultid="2649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1475" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3775" />
                    <RANKING order="2" place="2" resultid="3258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1476" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3593" />
                    <RANKING order="2" place="2" resultid="3182" />
                    <RANKING order="3" place="3" resultid="3462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1477" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2633" />
                    <RANKING order="2" place="2" resultid="3345" />
                    <RANKING order="3" place="3" resultid="3409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1478" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2119" />
                    <RANKING order="2" place="2" resultid="3653" />
                    <RANKING order="3" place="3" resultid="2623" />
                    <RANKING order="4" place="4" resultid="2986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1479" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2234" />
                    <RANKING order="2" place="2" resultid="2468" />
                    <RANKING order="3" place="3" resultid="2501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1480" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2426" />
                    <RANKING order="2" place="2" resultid="1907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2432" />
                    <RANKING order="2" place="2" resultid="2878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2418" />
                    <RANKING order="2" place="2" resultid="3108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3717" />
                    <RANKING order="2" place="2" resultid="3908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1484" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3915" />
                    <RANKING order="2" place="2" resultid="2201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1485" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1486" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1487" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1488" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1489" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4706" daytime="15:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4707" daytime="15:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4708" daytime="15:30" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1490" daytime="15:30" gender="M" number="25" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1491" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2662" />
                    <RANKING order="2" place="2" resultid="3632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1492" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3385" />
                    <RANKING order="2" place="2" resultid="2678" />
                    <RANKING order="3" place="3" resultid="2535" />
                    <RANKING order="4" place="4" resultid="3986" />
                    <RANKING order="5" place="5" resultid="2641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2350" />
                    <RANKING order="2" place="2" resultid="4042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2725" />
                    <RANKING order="2" place="-1" resultid="3271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1495" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3490" />
                    <RANKING order="2" place="2" resultid="3401" />
                    <RANKING order="3" place="3" resultid="3840" />
                    <RANKING order="4" place="4" resultid="4026" />
                    <RANKING order="5" place="-1" resultid="3171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1496" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3337" />
                    <RANKING order="2" place="2" resultid="3022" />
                    <RANKING order="3" place="3" resultid="2772" />
                    <RANKING order="4" place="4" resultid="3394" />
                    <RANKING order="5" place="5" resultid="2541" />
                    <RANKING order="6" place="6" resultid="2014" />
                    <RANKING order="7" place="7" resultid="2317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1497" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3756" />
                    <RANKING order="2" place="2" resultid="3921" />
                    <RANKING order="3" place="3" resultid="2604" />
                    <RANKING order="4" place="4" resultid="3845" />
                    <RANKING order="5" place="-1" resultid="1819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1498" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3794" />
                    <RANKING order="2" place="2" resultid="1970" />
                    <RANKING order="3" place="3" resultid="2186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1499" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3002" />
                    <RANKING order="2" place="2" resultid="1789" />
                    <RANKING order="3" place="3" resultid="3360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1500" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2494" />
                    <RANKING order="2" place="2" resultid="1886" />
                    <RANKING order="3" place="3" resultid="3929" />
                    <RANKING order="4" place="4" resultid="3733" />
                    <RANKING order="5" place="-1" resultid="1806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3299" />
                    <RANKING order="2" place="2" resultid="2027" />
                    <RANKING order="3" place="3" resultid="3941" />
                    <RANKING order="4" place="4" resultid="4806" />
                    <RANKING order="5" place="5" resultid="3724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1502" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2379" />
                    <RANKING order="2" place="2" resultid="2020" />
                    <RANKING order="3" place="3" resultid="1916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1503" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4017" />
                    <RANKING order="2" place="2" resultid="2196" />
                    <RANKING order="3" place="3" resultid="3617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1504" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1505" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1506" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4709" daytime="15:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4710" daytime="15:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4711" daytime="15:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4712" daytime="15:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4713" daytime="15:45" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1507" daytime="15:45" gender="F" number="26" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1508" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2910" />
                    <RANKING order="2" place="2" resultid="3088" />
                    <RANKING order="3" place="3" resultid="3100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1509" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3426" />
                    <RANKING order="2" place="2" resultid="3743" />
                    <RANKING order="3" place="3" resultid="3961" />
                    <RANKING order="4" place="4" resultid="3952" />
                    <RANKING order="5" place="5" resultid="3070" />
                    <RANKING order="6" place="-1" resultid="1827" />
                    <RANKING order="7" place="-1" resultid="3776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2169" />
                    <RANKING order="2" place="2" resultid="3235" />
                    <RANKING order="3" place="3" resultid="3463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1511" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2634" />
                    <RANKING order="2" place="2" resultid="3216" />
                    <RANKING order="3" place="3" resultid="3417" />
                    <RANKING order="4" place="4" resultid="3410" />
                    <RANKING order="5" place="5" resultid="3327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1512" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1794" />
                    <RANKING order="2" place="2" resultid="2370" />
                    <RANKING order="3" place="3" resultid="3243" />
                    <RANKING order="4" place="4" resultid="2961" />
                    <RANKING order="5" place="5" resultid="2409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1513" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3094" />
                    <RANKING order="2" place="2" resultid="2484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1514" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1895" />
                    <RANKING order="2" place="2" resultid="3374" />
                    <RANKING order="3" place="3" resultid="2277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2879" />
                    <RANKING order="2" place="2" resultid="2751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2595" />
                    <RANKING order="2" place="2" resultid="1799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat" />
                <AGEGROUP agegroupid="1518" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3212" />
                    <RANKING order="2" place="2" resultid="3789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1519" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1520" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1521" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1522" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1523" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4714" daytime="15:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4715" daytime="15:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4716" daytime="15:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4717" daytime="16:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1524" daytime="16:05" gender="M" number="27" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1525" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2941" />
                    <RANKING order="2" place="2" resultid="2820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1526" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2870" />
                    <RANKING order="2" place="2" resultid="2828" />
                    <RANKING order="3" place="3" resultid="3968" />
                    <RANKING order="4" place="4" resultid="3849" />
                    <RANKING order="5" place="5" resultid="3977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1527" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2720" />
                    <RANKING order="2" place="2" resultid="3819" />
                    <RANKING order="3" place="3" resultid="2691" />
                    <RANKING order="4" place="4" resultid="1991" />
                    <RANKING order="5" place="5" resultid="3606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1528" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3390" />
                    <RANKING order="2" place="2" resultid="3899" />
                    <RANKING order="3" place="3" resultid="2790" />
                    <RANKING order="4" place="4" resultid="2705" />
                    <RANKING order="5" place="5" resultid="3061" />
                    <RANKING order="6" place="6" resultid="2220" />
                    <RANKING order="7" place="7" resultid="2525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1529" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2178" />
                    <RANKING order="2" place="2" resultid="3990" />
                    <RANKING order="3" place="3" resultid="4023" />
                    <RANKING order="4" place="4" resultid="2314" />
                    <RANKING order="5" place="5" resultid="3812" />
                    <RANKING order="6" place="6" resultid="3841" />
                    <RANKING order="7" place="7" resultid="1854" />
                    <RANKING order="8" place="8" resultid="2697" />
                    <RANKING order="9" place="9" resultid="4005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1530" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2297" />
                    <RANKING order="2" place="2" resultid="1877" />
                    <RANKING order="3" place="3" resultid="3229" />
                    <RANKING order="4" place="4" resultid="3668" />
                    <RANKING order="5" place="5" resultid="1849" />
                    <RANKING order="6" place="6" resultid="3421" />
                    <RANKING order="7" place="7" resultid="3683" />
                    <RANKING order="8" place="8" resultid="2477" />
                    <RANKING order="9" place="9" resultid="2927" />
                    <RANKING order="10" place="-1" resultid="3481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1531" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3028" />
                    <RANKING order="2" place="2" resultid="2856" />
                    <RANKING order="3" place="3" resultid="2798" />
                    <RANKING order="4" place="4" resultid="3703" />
                    <RANKING order="5" place="5" resultid="3922" />
                    <RANKING order="6" place="6" resultid="2268" />
                    <RANKING order="7" place="7" resultid="2245" />
                    <RANKING order="8" place="-1" resultid="3474" />
                    <RANKING order="9" place="-1" resultid="3879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1532" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3190" />
                    <RANKING order="2" place="2" resultid="3625" />
                    <RANKING order="3" place="3" resultid="3795" />
                    <RANKING order="4" place="4" resultid="2971" />
                    <RANKING order="5" place="5" resultid="3502" />
                    <RANKING order="6" place="6" resultid="1949" />
                    <RANKING order="7" place="7" resultid="3206" />
                    <RANKING order="8" place="-1" resultid="2187" />
                    <RANKING order="9" place="-1" resultid="3442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1533" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3265" />
                    <RANKING order="2" place="2" resultid="2292" />
                    <RANKING order="3" place="3" resultid="2453" />
                    <RANKING order="4" place="4" resultid="3361" />
                    <RANKING order="5" place="5" resultid="2736" />
                    <RANKING order="6" place="6" resultid="3288" />
                    <RANKING order="7" place="-1" resultid="3036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1534" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2215" />
                    <RANKING order="2" place="2" resultid="1887" />
                    <RANKING order="3" place="3" resultid="1807" />
                    <RANKING order="4" place="4" resultid="3734" />
                    <RANKING order="5" place="5" resultid="3223" />
                    <RANKING order="6" place="6" resultid="3930" />
                    <RANKING order="7" place="-1" resultid="2385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1535" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2286" />
                    <RANKING order="2" place="2" resultid="3871" />
                    <RANKING order="3" place="3" resultid="2459" />
                    <RANKING order="4" place="4" resultid="3725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1536" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3857" />
                    <RANKING order="2" place="2" resultid="1985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1537" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2141" />
                    <RANKING order="2" place="2" resultid="3618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1538" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1539" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1540" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4718" daytime="16:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4719" daytime="16:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4720" daytime="16:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4721" daytime="16:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4722" daytime="16:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4723" daytime="16:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4724" daytime="16:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4725" daytime="16:35" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1541" daytime="16:40" gender="F" number="28" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1558" agemax="-1" agemin="-1" name="&quot;0&quot; 0-99 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="1559" agemax="119" agemin="100" name="&quot;A&quot; 100-119 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="1560" agemax="159" agemin="120" name="&quot;B&quot; 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3522" />
                    <RANKING order="2" place="2" resultid="3306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1561" agemax="199" agemin="160" name="&quot;C&quot; 160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3307" />
                    <RANKING order="2" place="2" resultid="3524" />
                    <RANKING order="3" place="3" resultid="2557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1562" agemax="239" agemin="200" name="&quot;D&quot; 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2551" />
                    <RANKING order="2" place="2" resultid="3114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1563" agemax="279" agemin="240" name="&quot;E&quot; 240-279 lat " calculate="TOTAL" />
                <AGEGROUP agegroupid="1564" agemax="-1" agemin="280" name="&quot;F&quot; 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4726" daytime="16:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1565" daytime="16:40" gender="M" number="29" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1566" agemax="-1" agemin="-1" name="&quot;0&quot; 0-99 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3525" />
                    <RANKING order="2" place="-1" resultid="3708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1567" agemax="119" agemin="100" name="&quot;A&quot; 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2836" />
                    <RANKING order="2" place="2" resultid="4039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1568" agemax="159" agemin="120" name="&quot;B&quot; 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4411" />
                    <RANKING order="2" place="2" resultid="3115" />
                    <RANKING order="3" place="3" resultid="4412" />
                    <RANKING order="4" place="-1" resultid="2994" />
                    <RANKING order="5" place="-1" resultid="2888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1569" agemax="199" agemin="160" name="&quot;C&quot; 160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3517" />
                    <RANKING order="2" place="2" resultid="3308" />
                    <RANKING order="3" place="3" resultid="3834" />
                    <RANKING order="4" place="4" resultid="2943" />
                    <RANKING order="5" place="5" resultid="2327" />
                    <RANKING order="6" place="6" resultid="3309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="239" agemin="200" name="&quot;D&quot; 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2803" />
                    <RANKING order="2" place="2" resultid="3519" />
                    <RANKING order="3" place="3" resultid="2564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1571" agemax="279" agemin="240" name="&quot;E&quot; 240-279 lat " calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2559" />
                    <RANKING order="2" place="2" resultid="2222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1572" agemax="-1" agemin="280" name="&quot;F&quot; 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4727" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4728" daytime="16:45" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1573" daytime="16:50" gender="F" number="30" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1581" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat" />
                <AGEGROUP agegroupid="1582" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2170" />
                    <RANKING order="2" place="2" resultid="3697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1584" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3157" />
                    <RANKING order="2" place="-1" resultid="3995" />
                    <RANKING order="3" place="-1" resultid="3346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1586" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2335" />
                    <RANKING order="2" place="2" resultid="2532" />
                    <RANKING order="3" place="3" resultid="2485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1587" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1908" />
                    <RANKING order="2" place="2" resultid="2516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1588" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat" />
                <AGEGROUP agegroupid="1589" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1590" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat" />
                <AGEGROUP agegroupid="1591" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat" />
                <AGEGROUP agegroupid="1592" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1593" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1594" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1595" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1596" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4785" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4786" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1597" daytime="17:05" gender="M" number="31" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1598" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3318" />
                    <RANKING order="2" place="2" resultid="2715" />
                    <RANKING order="3" place="3" resultid="1999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2179" />
                    <RANKING order="2" place="2" resultid="3402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3660" />
                    <RANKING order="2" place="2" resultid="3197" />
                    <RANKING order="3" place="3" resultid="3669" />
                    <RANKING order="4" place="4" resultid="3395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2269" />
                    <RANKING order="2" place="2" resultid="3880" />
                    <RANKING order="3" place="3" resultid="2438" />
                    <RANKING order="4" place="4" resultid="2605" />
                    <RANKING order="5" place="5" resultid="1930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3443" />
                    <RANKING order="2" place="2" resultid="2507" />
                    <RANKING order="3" place="3" resultid="1950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1606" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3037" />
                    <RANKING order="2" place="2" resultid="2133" />
                    <RANKING order="3" place="3" resultid="1841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1607" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2393" />
                    <RANKING order="2" place="2" resultid="2160" />
                    <RANKING order="3" place="3" resultid="4000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1608" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3284" />
                    <RANKING order="2" place="2" resultid="2028" />
                    <RANKING order="3" place="-1" resultid="2460" />
                    <RANKING order="4" place="-1" resultid="3872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1609" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1610" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1611" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1612" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1613" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4787" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4788" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4789" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4790" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2023-06-04" daytime="09:00" endtime="12:43" name="IV BLOK" number="4" warmupfrom="08:00" warmupuntil="08:55">
          <EVENTS>
            <EVENT eventid="1615" daytime="09:00" gender="F" number="32" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1617" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3744" />
                    <RANKING order="2" place="2" resultid="3953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3588" />
                    <RANKING order="2" place="2" resultid="3698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1620" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3158" />
                    <RANKING order="2" place="2" resultid="3996" />
                    <RANKING order="3" place="-1" resultid="3328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1621" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2309" />
                    <RANKING order="2" place="2" resultid="2624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1622" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat " />
                <AGEGROUP agegroupid="1623" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2427" />
                    <RANKING order="2" place="2" resultid="2517" />
                    <RANKING order="3" place="3" resultid="2278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1624" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3016" />
                    <RANKING order="2" place="2" resultid="3082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1625" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1626" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1627" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat" />
                <AGEGROUP agegroupid="1628" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1629" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1630" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1631" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1632" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4735" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4736" daytime="09:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1633" daytime="09:05" gender="M" number="33" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1634" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2821" />
                    <RANKING order="2" place="-1" resultid="2663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3801" />
                    <RANKING order="2" place="2" resultid="2833" />
                    <RANKING order="3" place="3" resultid="3969" />
                    <RANKING order="4" place="4" resultid="2829" />
                    <RANKING order="5" place="5" resultid="3164" />
                    <RANKING order="6" place="-1" resultid="3987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2810" />
                    <RANKING order="2" place="2" resultid="3435" />
                    <RANKING order="3" place="3" resultid="2716" />
                    <RANKING order="4" place="4" resultid="3820" />
                    <RANKING order="5" place="-1" resultid="2842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3900" />
                    <RANKING order="2" place="2" resultid="2791" />
                    <RANKING order="3" place="3" resultid="2706" />
                    <RANKING order="4" place="4" resultid="2526" />
                    <RANKING order="5" place="-1" resultid="3692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1638" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3491" />
                    <RANKING order="2" place="2" resultid="3806" />
                    <RANKING order="3" place="3" resultid="3151" />
                    <RANKING order="4" place="-1" resultid="3172" />
                    <RANKING order="5" place="-1" resultid="3813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1639" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3661" />
                    <RANKING order="2" place="2" resultid="1837" />
                    <RANKING order="3" place="3" resultid="3396" />
                    <RANKING order="4" place="4" resultid="1878" />
                    <RANKING order="5" place="5" resultid="3198" />
                    <RANKING order="6" place="6" resultid="3991" />
                    <RANKING order="7" place="7" resultid="3482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1640" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3029" />
                    <RANKING order="2" place="2" resultid="3863" />
                    <RANKING order="3" place="3" resultid="3757" />
                    <RANKING order="4" place="4" resultid="2857" />
                    <RANKING order="5" place="5" resultid="3704" />
                    <RANKING order="6" place="6" resultid="3881" />
                    <RANKING order="7" place="7" resultid="2246" />
                    <RANKING order="8" place="8" resultid="1931" />
                    <RANKING order="9" place="-1" resultid="2270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1641" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3191" />
                    <RANKING order="2" place="2" resultid="3444" />
                    <RANKING order="3" place="3" resultid="2508" />
                    <RANKING order="4" place="4" resultid="1951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1642" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1790" />
                    <RANKING order="2" place="2" resultid="2134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1643" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2394" />
                    <RANKING order="2" place="2" resultid="2366" />
                    <RANKING order="3" place="3" resultid="4001" />
                    <RANKING order="4" place="4" resultid="2161" />
                    <RANKING order="5" place="-1" resultid="2495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1644" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1645" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1918" />
                    <RANKING order="2" place="2" resultid="1986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1646" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1647" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1648" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1649" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4737" daytime="09:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4738" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4739" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4740" daytime="09:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4741" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4742" daytime="09:20" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1650" daytime="09:25" gender="F" number="34" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1651" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3777" />
                    <RANKING order="2" place="2" resultid="3259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1653" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3183" />
                    <RANKING order="2" place="2" resultid="2171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1654" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2635" />
                    <RANKING order="2" place="2" resultid="3143" />
                    <RANKING order="3" place="3" resultid="3411" />
                    <RANKING order="4" place="-1" resultid="3347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1655" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2120" />
                    <RANKING order="2" place="2" resultid="3654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1656" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2469" />
                    <RANKING order="2" place="2" resultid="2502" />
                    <RANKING order="3" place="3" resultid="2486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1657" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1909" />
                    <RANKING order="2" place="2" resultid="2518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1658" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1659" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3109" />
                    <RANKING order="2" place="-1" resultid="2597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1660" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1661" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1662" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1663" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1664" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1665" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1666" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4743" daytime="09:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4744" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4745" daytime="09:35" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1667" daytime="09:40" gender="M" number="35" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1668" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2816" />
                    <RANKING order="2" place="2" resultid="2536" />
                    <RANKING order="3" place="3" resultid="2679" />
                    <RANKING order="4" place="-1" resultid="3386" />
                    <RANKING order="5" place="-1" resultid="3988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1670" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2000" />
                    <RANKING order="2" place="-1" resultid="2351" />
                    <RANKING order="3" place="-1" resultid="4043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1671" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat" />
                <AGEGROUP agegroupid="1672" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3492" />
                    <RANKING order="2" place="2" resultid="3403" />
                    <RANKING order="3" place="3" resultid="2180" />
                    <RANKING order="4" place="-1" resultid="3173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1673" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3338" />
                    <RANKING order="2" place="2" resultid="3023" />
                    <RANKING order="3" place="3" resultid="2542" />
                    <RANKING order="4" place="4" resultid="3397" />
                    <RANKING order="5" place="5" resultid="3670" />
                    <RANKING order="6" place="6" resultid="2773" />
                    <RANKING order="7" place="7" resultid="2478" />
                    <RANKING order="8" place="-1" resultid="2318" />
                    <RANKING order="9" place="-1" resultid="3684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1674" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3758" />
                    <RANKING order="2" place="2" resultid="3923" />
                    <RANKING order="3" place="3" resultid="2606" />
                    <RANKING order="4" place="4" resultid="3846" />
                    <RANKING order="5" place="-1" resultid="1820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1675" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3796" />
                    <RANKING order="2" place="2" resultid="1971" />
                    <RANKING order="3" place="3" resultid="2188" />
                    <RANKING order="4" place="4" resultid="2972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1676" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3003" />
                    <RANKING order="2" place="2" resultid="3038" />
                    <RANKING order="3" place="3" resultid="3362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1677" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1888" />
                    <RANKING order="2" place="2" resultid="1808" />
                    <RANKING order="3" place="3" resultid="3931" />
                    <RANKING order="4" place="4" resultid="3735" />
                    <RANKING order="5" place="5" resultid="2127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1678" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3300" />
                    <RANKING order="2" place="2" resultid="2030" />
                    <RANKING order="3" place="3" resultid="3942" />
                    <RANKING order="4" place="4" resultid="3726" />
                    <RANKING order="5" place="-1" resultid="4807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1679" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2380" />
                    <RANKING order="2" place="2" resultid="2021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1680" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4018" />
                    <RANKING order="2" place="2" resultid="3619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1681" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1682" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1683" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4746" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4747" daytime="09:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4748" daytime="09:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4749" daytime="10:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4750" daytime="10:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1684" daytime="10:05" gender="F" number="36" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1685" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2651" />
                    <RANKING order="2" place="-1" resultid="3639" />
                    <RANKING order="3" place="-1" resultid="4012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1686" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3829" />
                    <RANKING order="2" place="2" resultid="3382" />
                    <RANKING order="3" place="3" resultid="1828" />
                    <RANKING order="4" place="4" resultid="3427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1687" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2258" />
                    <RANKING order="2" place="2" resultid="3178" />
                    <RANKING order="3" place="3" resultid="3594" />
                    <RANKING order="4" place="4" resultid="3333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1688" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2617" />
                    <RANKING order="2" place="2" resultid="3159" />
                    <RANKING order="3" place="3" resultid="3279" />
                    <RANKING order="4" place="-1" resultid="3611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1689" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2310" />
                    <RANKING order="2" place="2" resultid="2933" />
                    <RANKING order="3" place="3" resultid="2121" />
                    <RANKING order="4" place="4" resultid="3244" />
                    <RANKING order="5" place="5" resultid="4595" />
                    <RANKING order="6" place="6" resultid="2403" />
                    <RANKING order="7" place="-1" resultid="2410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1690" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2342" />
                    <RANKING order="2" place="2" resultid="3276" />
                    <RANKING order="3" place="3" resultid="3937" />
                    <RANKING order="4" place="4" resultid="2470" />
                    <RANKING order="5" place="5" resultid="2628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1691" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3375" />
                    <RANKING order="2" place="2" resultid="3496" />
                    <RANKING order="3" place="3" resultid="3784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1692" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2112" />
                    <RANKING order="2" place="2" resultid="3083" />
                    <RANKING order="3" place="3" resultid="3017" />
                    <RANKING order="4" place="4" resultid="3457" />
                    <RANKING order="5" place="5" resultid="2752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1693" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2420" />
                    <RANKING order="2" place="2" resultid="3110" />
                    <RANKING order="3" place="3" resultid="3121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1694" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1695" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3790" />
                    <RANKING order="2" place="2" resultid="2203" />
                    <RANKING order="3" place="3" resultid="1902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1696" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1697" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1698" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1699" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1700" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4751" daytime="10:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4752" daytime="10:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4753" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4754" daytime="10:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4755" daytime="10:15" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1701" daytime="10:15" gender="M" number="37" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1702" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2664" />
                    <RANKING order="2" place="-1" resultid="1961" />
                    <RANKING order="3" place="-1" resultid="2685" />
                    <RANKING order="4" place="-1" resultid="2942" />
                    <RANKING order="5" place="-1" resultid="3748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1703" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2785" />
                    <RANKING order="2" place="2" resultid="3048" />
                    <RANKING order="3" place="3" resultid="2817" />
                    <RANKING order="4" place="4" resultid="2834" />
                    <RANKING order="5" place="5" resultid="3978" />
                    <RANKING order="6" place="6" resultid="2642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1704" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2655" />
                    <RANKING order="2" place="2" resultid="3768" />
                    <RANKING order="3" place="3" resultid="3319" />
                    <RANKING order="4" place="4" resultid="2717" />
                    <RANKING order="5" place="5" resultid="3436" />
                    <RANKING order="6" place="6" resultid="3294" />
                    <RANKING order="7" place="7" resultid="3607" />
                    <RANKING order="8" place="-1" resultid="2843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1705" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2976" />
                    <RANKING order="2" place="2" resultid="3272" />
                    <RANKING order="3" place="3" resultid="3008" />
                    <RANKING order="4" place="4" resultid="2527" />
                    <RANKING order="5" place="-1" resultid="3062" />
                    <RANKING order="6" place="-1" resultid="3693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1706" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3152" />
                    <RANKING order="2" place="2" resultid="3644" />
                    <RANKING order="3" place="3" resultid="2322" />
                    <RANKING order="4" place="4" resultid="1855" />
                    <RANKING order="5" place="5" resultid="2698" />
                    <RANKING order="6" place="6" resultid="2325" />
                    <RANKING order="7" place="7" resultid="2008" />
                    <RANKING order="8" place="-1" resultid="4006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1707" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3251" />
                    <RANKING order="2" place="2" resultid="1879" />
                    <RANKING order="3" place="3" resultid="3676" />
                    <RANKING order="4" place="4" resultid="2543" />
                    <RANKING order="5" place="5" resultid="2848" />
                    <RANKING order="6" place="6" resultid="1832" />
                    <RANKING order="7" place="7" resultid="2252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1708" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3864" />
                    <RANKING order="2" place="2" resultid="3763" />
                    <RANKING order="3" place="3" resultid="2439" />
                    <RANKING order="4" place="-1" resultid="2862" />
                    <RANKING order="5" place="-1" resultid="3475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1709" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3450" />
                    <RANKING order="2" place="2" resultid="3503" />
                    <RANKING order="3" place="3" resultid="2509" />
                    <RANKING order="4" place="4" resultid="3207" />
                    <RANKING order="5" place="5" resultid="3000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1710" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3266" />
                    <RANKING order="2" place="2" resultid="1791" />
                    <RANKING order="3" place="3" resultid="2448" />
                    <RANKING order="4" place="4" resultid="2135" />
                    <RANKING order="5" place="-1" resultid="2361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1711" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2162" />
                    <RANKING order="2" place="2" resultid="2496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1712" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3285" />
                    <RANKING order="2" place="2" resultid="1863" />
                    <RANKING order="3" place="3" resultid="2867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1713" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2381" />
                    <RANKING order="2" place="2" resultid="2208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1714" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2197" />
                    <RANKING order="2" place="2" resultid="2142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1715" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1716" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1717" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4756" daytime="10:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4757" daytime="10:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4758" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4759" daytime="10:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4760" daytime="10:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4761" daytime="10:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4762" daytime="10:25" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1718" daytime="10:30" gender="X" number="38" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1735" agemax="-1" agemin="-1" name="&quot;0&quot; 0-99 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1736" agemax="119" agemin="100" name="&quot;A&quot; 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1737" agemax="159" agemin="120" name="&quot;B&quot; 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3311" />
                    <RANKING order="2" place="2" resultid="3508" />
                    <RANKING order="3" place="3" resultid="3312" />
                    <RANKING order="4" place="4" resultid="3111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1738" agemax="199" agemin="160" name="&quot;C&quot; 160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3510" />
                    <RANKING order="2" place="2" resultid="2946" />
                    <RANKING order="3" place="3" resultid="3313" />
                    <RANKING order="4" place="4" resultid="5400" />
                    <RANKING order="5" place="5" resultid="2563" />
                    <RANKING order="6" place="-1" resultid="3514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1739" agemax="239" agemin="200" name="&quot;D&quot; 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3310" />
                    <RANKING order="2" place="2" resultid="2554" />
                    <RANKING order="3" place="3" resultid="3116" />
                    <RANKING order="4" place="4" resultid="2562" />
                    <RANKING order="5" place="-1" resultid="3512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1740" agemax="279" agemin="240" name="&quot;E&quot; 240-279 lat " calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2561" />
                    <RANKING order="2" place="2" resultid="3945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1741" agemax="-1" agemin="280" name="&quot;F&quot; 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4763" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4764" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4765" daytime="10:35" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1742" daytime="10:40" gender="F" number="39" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1750" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2912" />
                    <RANKING order="2" place="2" resultid="3089" />
                    <RANKING order="3" place="3" resultid="3101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1751" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3428" />
                    <RANKING order="2" place="2" resultid="3954" />
                    <RANKING order="3" place="3" resultid="3830" />
                    <RANKING order="4" place="4" resultid="3071" />
                    <RANKING order="5" place="-1" resultid="3778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1752" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2172" />
                    <RANKING order="2" place="2" resultid="3699" />
                    <RANKING order="3" place="3" resultid="3236" />
                    <RANKING order="4" place="-1" resultid="3464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1753" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2636" />
                    <RANKING order="2" place="2" resultid="3217" />
                    <RANKING order="3" place="3" resultid="2915" />
                    <RANKING order="4" place="4" resultid="3144" />
                    <RANKING order="5" place="5" resultid="2618" />
                    <RANKING order="6" place="6" resultid="3418" />
                    <RANKING order="7" place="-1" resultid="3329" />
                    <RANKING order="8" place="-1" resultid="3348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1754" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1795" />
                    <RANKING order="2" place="2" resultid="2371" />
                    <RANKING order="3" place="3" resultid="3245" />
                    <RANKING order="4" place="4" resultid="2411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1755" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2336" />
                    <RANKING order="2" place="2" resultid="3095" />
                    <RANKING order="3" place="3" resultid="2533" />
                    <RANKING order="4" place="4" resultid="2487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1756" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1896" />
                    <RANKING order="2" place="2" resultid="3376" />
                    <RANKING order="3" place="3" resultid="2279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1757" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1758" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1759" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1760" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1761" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat" />
                <AGEGROUP agegroupid="1762" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat" />
                <AGEGROUP agegroupid="1763" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1764" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1765" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4791" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4792" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4793" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4794" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1766" daytime="11:10" gender="M" number="40" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1767" agemax="24" agemin="20" name="&quot;0&quot; 20-24 lat" />
                <AGEGROUP agegroupid="1768" agemax="29" agemin="25" name="&quot;A&quot; 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3970" />
                    <RANKING order="2" place="2" resultid="2830" />
                    <RANKING order="3" place="3" resultid="3850" />
                    <RANKING order="4" place="4" resultid="3979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1769" agemax="34" agemin="30" name="&quot;B&quot; 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3320" />
                    <RANKING order="2" place="2" resultid="3821" />
                    <RANKING order="3" place="3" resultid="2692" />
                    <RANKING order="4" place="4" resultid="1943" />
                    <RANKING order="5" place="5" resultid="2001" />
                    <RANKING order="6" place="6" resultid="1992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1770" agemax="39" agemin="35" name="&quot;C&quot; 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3391" />
                    <RANKING order="2" place="2" resultid="3901" />
                    <RANKING order="3" place="3" resultid="2792" />
                    <RANKING order="4" place="4" resultid="2707" />
                    <RANKING order="5" place="5" resultid="3063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1771" agemax="44" agemin="40" name="&quot;D&quot; 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2181" />
                    <RANKING order="2" place="2" resultid="3814" />
                    <RANKING order="3" place="3" resultid="4024" />
                    <RANKING order="4" place="4" resultid="3404" />
                    <RANKING order="5" place="5" resultid="1856" />
                    <RANKING order="6" place="6" resultid="2699" />
                    <RANKING order="7" place="7" resultid="2009" />
                    <RANKING order="8" place="-1" resultid="3807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1772" agemax="49" agemin="45" name="&quot;E&quot; 45-49 lat ">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3662" />
                    <RANKING order="2" place="2" resultid="3671" />
                    <RANKING order="3" place="3" resultid="2296" />
                    <RANKING order="4" place="4" resultid="3230" />
                    <RANKING order="5" place="5" resultid="1850" />
                    <RANKING order="6" place="6" resultid="3199" />
                    <RANKING order="7" place="7" resultid="3252" />
                    <RANKING order="8" place="8" resultid="2741" />
                    <RANKING order="9" place="9" resultid="3685" />
                    <RANKING order="10" place="10" resultid="2849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1773" agemax="54" agemin="50" name="&quot;F&quot; 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3030" />
                    <RANKING order="2" place="2" resultid="2799" />
                    <RANKING order="3" place="3" resultid="2858" />
                    <RANKING order="4" place="4" resultid="3705" />
                    <RANKING order="5" place="5" resultid="3882" />
                    <RANKING order="6" place="6" resultid="2607" />
                    <RANKING order="7" place="7" resultid="2440" />
                    <RANKING order="8" place="-1" resultid="2271" />
                    <RANKING order="9" place="-1" resultid="3476" />
                    <RANKING order="10" place="-1" resultid="3924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1774" agemax="59" agemin="55" name="&quot;G&quot; 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3192" />
                    <RANKING order="2" place="2" resultid="3626" />
                    <RANKING order="3" place="3" resultid="3445" />
                    <RANKING order="4" place="4" resultid="2189" />
                    <RANKING order="5" place="5" resultid="3208" />
                    <RANKING order="6" place="6" resultid="1952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1775" agemax="64" agemin="60" name="&quot;H&quot; 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3267" />
                    <RANKING order="2" place="2" resultid="2291" />
                    <RANKING order="3" place="3" resultid="2454" />
                    <RANKING order="4" place="4" resultid="3363" />
                    <RANKING order="5" place="5" resultid="1842" />
                    <RANKING order="6" place="6" resultid="3289" />
                    <RANKING order="7" place="-1" resultid="3039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1776" agemax="69" agemin="65" name="&quot;I&quot; 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1889" />
                    <RANKING order="2" place="2" resultid="3224" />
                    <RANKING order="3" place="3" resultid="3736" />
                    <RANKING order="4" place="4" resultid="2128" />
                    <RANKING order="5" place="-1" resultid="1809" />
                    <RANKING order="6" place="-1" resultid="2386" />
                    <RANKING order="7" place="-1" resultid="2395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1777" agemax="74" agemin="70" name="&quot;J&quot; 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2287" />
                    <RANKING order="2" place="2" resultid="3873" />
                    <RANKING order="3" place="3" resultid="2461" />
                    <RANKING order="4" place="4" resultid="5399" />
                    <RANKING order="5" place="5" resultid="3727" />
                    <RANKING order="6" place="-1" resultid="2868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1778" agemax="79" agemin="75" name="&quot;K&quot; 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3858" />
                    <RANKING order="2" place="2" resultid="1987" />
                    <RANKING order="3" place="-1" resultid="1919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1779" agemax="84" agemin="80" name="&quot;L&quot; 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2143" />
                    <RANKING order="2" place="2" resultid="3620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1780" agemax="89" agemin="85" name="&quot;M&quot; 85-89 lat" />
                <AGEGROUP agegroupid="1781" agemax="94" agemin="90" name="&quot;N&quot; 90-94 lat" />
                <AGEGROUP agegroupid="1782" agemax="99" agemin="95" name="&quot;O&quot; 95-99 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4795" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4796" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4797" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4798" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4799" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4800" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4801" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4802" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="STKAR" nation="POL" region="14" clubid="2906" name="St. Pływ. Sebastiana Karasia Łomianki" shortname="St. Pływ. Sebastiana Karasia">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Grabkowski" birthdate="1981-03-27" gender="M" nation="POL" athleteid="2921">
              <RESULTS>
                <RESULT eventid="1090" points="389" swimtime="00:00:31.76" resultid="2922" heatid="4610" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1320" points="362" swimtime="00:01:11.85" resultid="2923" heatid="4670" lane="9" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Diaby-Lipka" birthdate="1980-08-30" gender="F" nation="POL" athleteid="2919">
              <RESULTS>
                <RESULT eventid="1234" points="548" swimtime="00:00:36.19" resultid="2920" heatid="4643" lane="8" entrytime="00:00:35.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Karczewski" birthdate="1974-07-07" gender="M" nation="POL" athleteid="2934">
              <RESULTS>
                <RESULT comment="K7 - Pływak wykonał ruchy ramion nie w tej samej poziomej płaszczyźnie." eventid="1124" status="DSQ" swimtime="00:04:00.87" resultid="2935" heatid="4622" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.78" />
                    <SPLIT distance="100" swimtime="00:02:00.69" />
                    <SPLIT distance="150" swimtime="00:03:08.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Przekroczony limit czasu" eventid="1216" status="OTL" swimtime="00:29:17.86" resultid="2936" heatid="4638" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.25" />
                    <SPLIT distance="100" swimtime="00:01:48.80" />
                    <SPLIT distance="150" swimtime="00:02:47.12" />
                    <SPLIT distance="200" swimtime="00:03:45.82" />
                    <SPLIT distance="250" swimtime="00:04:44.27" />
                    <SPLIT distance="300" swimtime="00:05:42.36" />
                    <SPLIT distance="350" swimtime="00:06:40.68" />
                    <SPLIT distance="400" swimtime="00:07:39.68" />
                    <SPLIT distance="450" swimtime="00:08:37.81" />
                    <SPLIT distance="500" swimtime="00:09:35.27" />
                    <SPLIT distance="550" swimtime="00:10:34.01" />
                    <SPLIT distance="600" swimtime="00:11:32.44" />
                    <SPLIT distance="650" swimtime="00:12:32.37" />
                    <SPLIT distance="700" swimtime="00:13:31.02" />
                    <SPLIT distance="750" swimtime="00:14:30.47" />
                    <SPLIT distance="800" swimtime="00:15:27.77" />
                    <SPLIT distance="850" swimtime="00:16:26.39" />
                    <SPLIT distance="900" swimtime="00:17:24.05" />
                    <SPLIT distance="950" swimtime="00:18:22.51" />
                    <SPLIT distance="1000" swimtime="00:19:21.49" />
                    <SPLIT distance="1050" swimtime="00:20:22.02" />
                    <SPLIT distance="1100" swimtime="00:21:22.70" />
                    <SPLIT distance="1150" swimtime="00:22:23.69" />
                    <SPLIT distance="1200" swimtime="00:23:23.21" />
                    <SPLIT distance="1250" swimtime="00:24:21.76" />
                    <SPLIT distance="1300" swimtime="00:25:24.07" />
                    <SPLIT distance="1350" swimtime="00:26:25.72" />
                    <SPLIT distance="1400" swimtime="00:27:27.34" />
                    <SPLIT distance="1450" swimtime="00:28:25.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Karczewski" birthdate="1974-07-07" gender="M" nation="POL" athleteid="2924">
              <RESULTS>
                <RESULT eventid="1090" points="376" swimtime="00:00:32.62" resultid="2925" heatid="4609" lane="8" entrytime="00:00:32.40" />
                <RESULT eventid="1320" points="347" swimtime="00:01:14.33" resultid="2926" heatid="4667" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="298" swimtime="00:02:56.28" resultid="2927" heatid="4720" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:01:25.52" />
                    <SPLIT distance="150" swimtime="00:02:12.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Fuliński" birthdate="1982-03-06" gender="M" nation="POL" athleteid="2916">
              <RESULTS>
                <RESULT eventid="1090" points="638" swimtime="00:00:26.94" resultid="2917" heatid="4614" lane="4" entrytime="00:00:26.97" />
                <RESULT eventid="1320" points="625" swimtime="00:00:59.87" resultid="2918" heatid="4673" lane="4" entrytime="00:00:59.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Janicka" birthdate="1984-04-18" gender="F" nation="POL" athleteid="2913">
              <RESULTS>
                <RESULT eventid="1059" points="548" swimtime="00:00:31.74" resultid="2914" heatid="4601" lane="7" entrytime="00:00:30.17" />
                <RESULT eventid="1742" points="460" swimtime="00:05:44.65" resultid="2915" heatid="4792" lane="1" entrytime="00:05:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                    <SPLIT distance="150" swimtime="00:02:04.09" />
                    <SPLIT distance="200" swimtime="00:02:48.79" />
                    <SPLIT distance="250" swimtime="00:03:33.62" />
                    <SPLIT distance="300" swimtime="00:04:18.71" />
                    <SPLIT distance="350" swimtime="00:05:03.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kotarski" birthdate="2002-05-07" gender="M" nation="POL" athleteid="2937">
              <RESULTS>
                <RESULT eventid="1090" swimtime="00:00:25.03" resultid="2938" heatid="4617" lane="5" entrytime="00:00:24.00" />
                <RESULT eventid="1320" swimtime="00:00:54.43" resultid="2939" heatid="4675" lane="5" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" swimtime="00:00:27.03" resultid="2940" heatid="4705" lane="3" entrytime="00:00:25.50" />
                <RESULT eventid="1524" swimtime="00:02:06.81" resultid="2941" heatid="4725" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:03.49" />
                    <SPLIT distance="150" swimtime="00:01:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="2942" heatid="4762" lane="6" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Łukasiuk" birthdate="1980-01-02" gender="F" nation="POL" athleteid="2930">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="2931" heatid="4600" lane="9" entrytime="00:00:33.50" />
                <RESULT eventid="1404" points="438" swimtime="00:01:35.17" resultid="2932" heatid="4687" lane="6" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="460" swimtime="00:00:41.99" resultid="2933" heatid="4754" lane="8" entrytime="00:00:42.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Witek" birthdate="1984-09-22" gender="M" nation="POL" athleteid="2928">
              <RESULTS>
                <RESULT eventid="1090" points="496" swimtime="00:00:28.74" resultid="2929" heatid="4614" lane="8" entrytime="00:00:27.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Borys" birthdate="2000-05-01" gender="F" nation="POL" athleteid="2907">
              <RESULTS>
                <RESULT eventid="1234" swimtime="00:00:33.96" resultid="2908" heatid="4643" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1473" swimtime="00:01:13.33" resultid="2909" heatid="4708" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" swimtime="00:02:26.15" resultid="2910" heatid="4717" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:47.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" swimtime="00:02:38.77" resultid="2911" heatid="4745" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:16.53" />
                    <SPLIT distance="150" swimtime="00:01:57.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" swimtime="00:05:06.81" resultid="2912" heatid="4791" lane="7" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:12.95" />
                    <SPLIT distance="150" swimtime="00:01:52.11" />
                    <SPLIT distance="200" swimtime="00:02:31.08" />
                    <SPLIT distance="250" swimtime="00:03:09.77" />
                    <SPLIT distance="300" swimtime="00:03:48.93" />
                    <SPLIT distance="350" swimtime="00:04:28.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="508" swimtime="00:01:58.93" resultid="2943" heatid="4727" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                    <SPLIT distance="100" swimtime="00:00:54.95" />
                    <SPLIT distance="150" swimtime="00:01:27.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2916" number="1" />
                    <RELAYPOSITION athleteid="2928" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2924" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="2921" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="396" swimtime="00:02:23.57" resultid="2944" heatid="4683" lane="8">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:51.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2924" number="1" />
                    <RELAYPOSITION athleteid="2916" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2928" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="2921" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1141" points="545" swimtime="00:02:05.13" resultid="2945" heatid="4629" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.90" />
                    <SPLIT distance="100" swimtime="00:00:57.95" />
                    <SPLIT distance="150" swimtime="00:01:26.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2916" number="1" />
                    <RELAYPOSITION athleteid="2913" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2928" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2930" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1718" points="572" swimtime="00:02:16.41" resultid="2946" heatid="4764" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:18.22" />
                    <SPLIT distance="150" swimtime="00:01:50.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2919" number="1" />
                    <RELAYPOSITION athleteid="2930" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="2928" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2916" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SPGRO" nation="POL" region="14" clubid="2311" name="UKS SPARTA Grodzisk Mazowiecki" shortname="SPARTA Grodzisk Mazowiecki">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Głowa" birthdate="1979-10-08" gender="M" nation="POL" athleteid="2312">
              <RESULTS>
                <RESULT eventid="1320" points="569" swimtime="00:01:01.77" resultid="2313" heatid="4672" lane="9" entrytime="00:01:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="485" swimtime="00:02:24.56" resultid="2314" heatid="4723" lane="0" entrytime="00:02:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                    <SPLIT distance="150" swimtime="00:01:47.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Płotnicki" birthdate="1982-10-08" gender="M" nation="POL" athleteid="2323">
              <RESULTS>
                <RESULT eventid="1422" points="331" swimtime="00:01:31.87" resultid="2324" heatid="4692" lane="8" entrytime="00:01:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="364" swimtime="00:00:40.38" resultid="2325" heatid="4759" lane="0" entrytime="00:00:40.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Zieliński" birthdate="1980-05-18" gender="M" nation="POL" athleteid="2319">
              <RESULTS>
                <RESULT eventid="1286" points="454" swimtime="00:03:00.23" resultid="2320" heatid="4657" lane="5" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:26.48" />
                    <SPLIT distance="150" swimtime="00:02:12.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="444" swimtime="00:01:23.34" resultid="2321" heatid="4692" lane="2" entrytime="00:01:21.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="508" swimtime="00:00:36.14" resultid="2322" heatid="4760" lane="1" entrytime="00:00:37.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Plich" birthdate="1978-06-21" gender="M" nation="POL" athleteid="2315">
              <RESULTS>
                <RESULT eventid="1252" points="396" swimtime="00:00:37.59" resultid="2316" heatid="4648" lane="9" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1490" points="418" swimtime="00:01:20.39" resultid="2317" heatid="4711" lane="5" entrytime="00:01:22.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" status="DNS" swimtime="00:00:00.00" resultid="2318" heatid="4748" lane="3" entrytime="00:03:10.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="455" swimtime="00:02:17.03" resultid="2326" heatid="4684" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:50.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2315" number="1" />
                    <RELAYPOSITION athleteid="2319" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="2323" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2312" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="480" swimtime="00:02:01.16" resultid="2327" heatid="4727" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="100" swimtime="00:00:59.91" />
                    <SPLIT distance="150" swimtime="00:01:34.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2315" number="1" />
                    <RELAYPOSITION athleteid="2319" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="2323" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="2312" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="05806" nation="POL" region="06" clubid="3710" name="IKS DRUGA STRONA SPORTU Kraków" shortname="DRUGA STRONA SPORTU Kraków">
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Rupp" birthdate="1956-03-06" gender="F" nation="POL" license="505806600021" athleteid="3711">
              <RESULTS>
                <RESULT eventid="1059" points="176" swimtime="00:00:51.91" resultid="3712" heatid="4597" lane="1" entrytime="00:00:53.24" />
                <RESULT eventid="1107" points="169" swimtime="00:05:10.16" resultid="3713" heatid="4618" lane="5" entrytime="00:04:57.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.46" />
                    <SPLIT distance="100" swimtime="00:02:32.59" />
                    <SPLIT distance="150" swimtime="00:04:01.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="160" swimtime="00:01:01.77" resultid="3714" heatid="4640" lane="5" entrytime="00:01:02.00" />
                <RESULT eventid="1303" points="147" swimtime="00:02:02.87" resultid="3715" heatid="4659" lane="6" entrytime="00:02:01.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="63" swimtime="00:01:22.55" resultid="3716" heatid="4694" lane="6" entrytime="00:01:12.12" />
                <RESULT eventid="1473" points="171" swimtime="00:02:14.18" resultid="3717" heatid="4706" lane="6" entrytime="00:02:15.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="58" swimtime="00:03:09.77" resultid="3718" heatid="4735" lane="1" entrytime="00:02:56.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="199" swimtime="00:04:47.15" resultid="3719" heatid="4743" lane="5" entrytime="00:04:42.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.83" />
                    <SPLIT distance="100" swimtime="00:02:22.50" />
                    <SPLIT distance="150" swimtime="00:03:36.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogdan" lastname="Szczurek" birthdate="1952-02-07" gender="M" nation="POL" license="105806700037" athleteid="3720">
              <RESULTS>
                <RESULT eventid="1090" points="162" swimtime="00:00:50.73" resultid="3721" heatid="4605" lane="0" entrytime="00:00:49.18" />
                <RESULT eventid="1252" points="179" swimtime="00:00:59.48" resultid="3722" heatid="4646" lane="0" entrytime="00:00:58.11" />
                <RESULT eventid="1320" points="140" swimtime="00:02:01.72" resultid="3723" heatid="4665" lane="7" entrytime="00:01:53.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="187" swimtime="00:02:08.36" resultid="3724" heatid="4709" lane="5" entrytime="00:02:04.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="137" swimtime="00:04:37.78" resultid="3725" heatid="4718" lane="4" entrytime="00:04:21.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.54" />
                    <SPLIT distance="100" swimtime="00:02:11.19" />
                    <SPLIT distance="150" swimtime="00:03:24.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="186" swimtime="00:04:40.39" resultid="3726" heatid="4747" lane="9" entrytime="00:04:26.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.66" />
                    <SPLIT distance="100" swimtime="00:02:18.51" />
                    <SPLIT distance="150" swimtime="00:03:31.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="142" swimtime="00:09:41.76" resultid="3727" heatid="4801" lane="9" entrytime="00:08:58.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.13" />
                    <SPLIT distance="100" swimtime="00:02:13.78" />
                    <SPLIT distance="150" swimtime="00:03:26.05" />
                    <SPLIT distance="200" swimtime="00:04:41.03" />
                    <SPLIT distance="250" swimtime="00:05:56.06" />
                    <SPLIT distance="300" swimtime="00:07:14.00" />
                    <SPLIT distance="350" swimtime="00:08:29.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01914" nation="POL" region="14" clubid="1920" name="UŚKS Ostrołęka" shortname="UŚKS OStrołęka">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="Janczewski" birthdate="1990-12-06" gender="M" nation="POL" athleteid="2353">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="2354" heatid="4615" lane="4" entrytime="00:00:25.70" />
                <RESULT eventid="1124" points="662" swimtime="00:02:20.12" resultid="2355" heatid="4628" lane="2" entrytime="00:02:25.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                    <SPLIT distance="100" swimtime="00:01:05.52" />
                    <SPLIT distance="150" swimtime="00:01:46.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="521" swimtime="00:10:06.77" resultid="2356" heatid="4636" lane="1" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:11.11" />
                    <SPLIT distance="150" swimtime="00:01:48.95" />
                    <SPLIT distance="200" swimtime="00:02:27.42" />
                    <SPLIT distance="250" swimtime="00:03:06.04" />
                    <SPLIT distance="300" swimtime="00:03:45.09" />
                    <SPLIT distance="350" swimtime="00:04:24.00" />
                    <SPLIT distance="400" swimtime="00:05:03.16" />
                    <SPLIT distance="450" swimtime="00:05:41.70" />
                    <SPLIT distance="500" swimtime="00:06:20.40" />
                    <SPLIT distance="550" swimtime="00:06:59.04" />
                    <SPLIT distance="600" swimtime="00:07:37.16" />
                    <SPLIT distance="650" swimtime="00:08:15.52" />
                    <SPLIT distance="700" swimtime="00:08:53.58" />
                    <SPLIT distance="750" swimtime="00:09:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Ambroziak" birthdate="1964-01-01" gender="M" nation="POL" athleteid="1921">
              <RESULTS>
                <RESULT eventid="1124" points="248" swimtime="00:03:43.78" resultid="1922" heatid="4624" lane="7" entrytime="00:03:44.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                    <SPLIT distance="100" swimtime="00:01:51.73" />
                    <SPLIT distance="150" swimtime="00:02:55.56" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Przekroczony limit czasu" eventid="1216" status="OTL" swimtime="00:27:16.37" resultid="1923" heatid="4639" lane="9" entrytime="00:26:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                    <SPLIT distance="100" swimtime="00:01:33.67" />
                    <SPLIT distance="150" swimtime="00:02:25.51" />
                    <SPLIT distance="200" swimtime="00:03:20.20" />
                    <SPLIT distance="250" swimtime="00:04:15.33" />
                    <SPLIT distance="300" swimtime="00:05:10.35" />
                    <SPLIT distance="350" swimtime="00:06:05.38" />
                    <SPLIT distance="400" swimtime="00:07:01.29" />
                    <SPLIT distance="450" swimtime="00:07:57.29" />
                    <SPLIT distance="500" swimtime="00:08:53.17" />
                    <SPLIT distance="550" swimtime="00:09:49.08" />
                    <SPLIT distance="600" swimtime="00:10:44.84" />
                    <SPLIT distance="650" swimtime="00:11:40.07" />
                    <SPLIT distance="700" swimtime="00:12:35.50" />
                    <SPLIT distance="750" swimtime="00:13:30.79" />
                    <SPLIT distance="800" swimtime="00:14:26.30" />
                    <SPLIT distance="850" swimtime="00:15:21.91" />
                    <SPLIT distance="900" swimtime="00:16:16.27" />
                    <SPLIT distance="950" swimtime="00:17:11.97" />
                    <SPLIT distance="1000" swimtime="00:18:06.14" />
                    <SPLIT distance="1050" swimtime="00:19:02.27" />
                    <SPLIT distance="1100" swimtime="00:19:56.89" />
                    <SPLIT distance="1150" swimtime="00:20:52.94" />
                    <SPLIT distance="1200" swimtime="00:21:47.31" />
                    <SPLIT distance="1250" swimtime="00:22:42.45" />
                    <SPLIT distance="1300" swimtime="00:23:37.56" />
                    <SPLIT distance="1350" swimtime="00:24:32.81" />
                    <SPLIT distance="1400" swimtime="00:25:28.44" />
                    <SPLIT distance="1450" swimtime="00:26:24.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="319" swimtime="00:01:21.91" resultid="4044" heatid="4669" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02016" nation="POL" region="16" clubid="3728" name="Koszalińskie TKKF">
          <ATHLETES>
            <ATHLETE firstname="Marian" lastname="Lasowy" birthdate="1955-07-15" gender="M" nation="POL" license="502016700001" athleteid="3729">
              <RESULTS>
                <RESULT eventid="1216" points="349" swimtime="00:27:45.92" resultid="3730" heatid="4638" lane="3" entrytime="00:27:04.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.37" />
                    <SPLIT distance="100" swimtime="00:01:40.62" />
                    <SPLIT distance="150" swimtime="00:02:36.05" />
                    <SPLIT distance="200" swimtime="00:03:31.65" />
                    <SPLIT distance="250" swimtime="00:04:27.63" />
                    <SPLIT distance="300" swimtime="00:05:21.56" />
                    <SPLIT distance="350" swimtime="00:06:17.24" />
                    <SPLIT distance="400" swimtime="00:07:12.97" />
                    <SPLIT distance="450" swimtime="00:08:07.33" />
                    <SPLIT distance="500" swimtime="00:09:03.82" />
                    <SPLIT distance="550" swimtime="00:09:58.33" />
                    <SPLIT distance="600" swimtime="00:10:54.49" />
                    <SPLIT distance="650" swimtime="00:11:53.11" />
                    <SPLIT distance="700" swimtime="00:12:47.58" />
                    <SPLIT distance="750" swimtime="00:13:43.73" />
                    <SPLIT distance="800" swimtime="00:14:40.33" />
                    <SPLIT distance="850" swimtime="00:15:36.32" />
                    <SPLIT distance="900" swimtime="00:16:34.01" />
                    <SPLIT distance="950" swimtime="00:17:30.94" />
                    <SPLIT distance="1000" swimtime="00:18:26.37" />
                    <SPLIT distance="1050" swimtime="00:19:22.88" />
                    <SPLIT distance="1100" swimtime="00:20:19.38" />
                    <SPLIT distance="1150" swimtime="00:21:16.03" />
                    <SPLIT distance="1200" swimtime="00:22:11.48" />
                    <SPLIT distance="1250" swimtime="00:23:08.00" />
                    <SPLIT distance="1300" swimtime="00:24:06.16" />
                    <SPLIT distance="1350" swimtime="00:24:55.70" />
                    <SPLIT distance="1400" swimtime="00:25:57.32" />
                    <SPLIT distance="1450" swimtime="00:26:53.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="213" swimtime="00:04:30.12" resultid="3731" heatid="4655" lane="3" entrytime="00:04:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.13" />
                    <SPLIT distance="100" swimtime="00:02:06.00" />
                    <SPLIT distance="150" swimtime="00:03:19.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="290" swimtime="00:01:29.78" resultid="3732" heatid="4667" lane="9" entrytime="00:01:29.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="195" swimtime="00:01:57.43" resultid="3733" heatid="4709" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="250" swimtime="00:03:25.24" resultid="3734" heatid="4719" lane="4" entrytime="00:03:20.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                    <SPLIT distance="100" swimtime="00:01:41.18" />
                    <SPLIT distance="150" swimtime="00:02:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="201" swimtime="00:04:18.73" resultid="3735" heatid="4746" lane="4" entrytime="00:04:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.96" />
                    <SPLIT distance="100" swimtime="00:02:08.26" />
                    <SPLIT distance="150" swimtime="00:03:14.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="259" swimtime="00:07:15.23" resultid="3736" heatid="4800" lane="0" entrytime="00:07:02.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.16" />
                    <SPLIT distance="100" swimtime="00:01:44.34" />
                    <SPLIT distance="150" swimtime="00:02:40.33" />
                    <SPLIT distance="200" swimtime="00:03:36.39" />
                    <SPLIT distance="250" swimtime="00:04:31.94" />
                    <SPLIT distance="300" swimtime="00:05:27.36" />
                    <SPLIT distance="350" swimtime="00:06:24.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00309" nation="POL" region="09" clubid="1783" name="MKS JUVENIA Białystok" shortname="JUVENIA Białystok">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Michalik" birthdate="1979-01-01" gender="F" nation="POL" license="500309600228" athleteid="1792">
              <RESULTS>
                <RESULT eventid="1199" points="557" swimtime="00:21:15.46" resultid="1793" heatid="4637" lane="4" entrytime="00:20:24.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:16.96" />
                    <SPLIT distance="150" swimtime="00:01:57.50" />
                    <SPLIT distance="200" swimtime="00:02:39.65" />
                    <SPLIT distance="250" swimtime="00:03:21.87" />
                    <SPLIT distance="300" swimtime="00:04:04.78" />
                    <SPLIT distance="350" swimtime="00:04:46.82" />
                    <SPLIT distance="400" swimtime="00:05:28.96" />
                    <SPLIT distance="450" swimtime="00:06:11.53" />
                    <SPLIT distance="500" swimtime="00:06:54.70" />
                    <SPLIT distance="550" swimtime="00:07:37.81" />
                    <SPLIT distance="600" swimtime="00:08:21.41" />
                    <SPLIT distance="650" swimtime="00:09:04.07" />
                    <SPLIT distance="700" swimtime="00:09:46.76" />
                    <SPLIT distance="750" swimtime="00:10:29.66" />
                    <SPLIT distance="800" swimtime="00:11:13.18" />
                    <SPLIT distance="850" swimtime="00:11:56.08" />
                    <SPLIT distance="900" swimtime="00:12:39.30" />
                    <SPLIT distance="950" swimtime="00:13:22.24" />
                    <SPLIT distance="1000" swimtime="00:14:05.99" />
                    <SPLIT distance="1050" swimtime="00:14:49.15" />
                    <SPLIT distance="1100" swimtime="00:15:33.33" />
                    <SPLIT distance="1150" swimtime="00:16:16.55" />
                    <SPLIT distance="1200" swimtime="00:17:00.55" />
                    <SPLIT distance="1250" swimtime="00:17:44.04" />
                    <SPLIT distance="1300" swimtime="00:18:28.22" />
                    <SPLIT distance="1350" swimtime="00:19:11.21" />
                    <SPLIT distance="1400" swimtime="00:19:54.83" />
                    <SPLIT distance="1450" swimtime="00:20:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="687" swimtime="00:02:26.45" resultid="1794" heatid="4717" lane="2" entrytime="00:02:22.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:11.24" />
                    <SPLIT distance="150" swimtime="00:01:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="571" swimtime="00:05:16.78" resultid="1795" heatid="4791" lane="4" entrytime="00:05:03.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                    <SPLIT distance="150" swimtime="00:01:54.24" />
                    <SPLIT distance="200" swimtime="00:02:34.41" />
                    <SPLIT distance="250" swimtime="00:03:15.17" />
                    <SPLIT distance="300" swimtime="00:03:56.03" />
                    <SPLIT distance="350" swimtime="00:04:37.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Wasilewicz" birthdate="1959-01-01" gender="F" nation="POL" license="500309600230" athleteid="1796">
              <RESULTS>
                <RESULT eventid="1059" points="421" swimtime="00:00:38.55" resultid="1797" heatid="4598" lane="6" entrytime="00:00:38.53" />
                <RESULT eventid="1303" points="360" swimtime="00:01:29.71" resultid="1798" heatid="4660" lane="2" entrytime="00:01:29.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="300" swimtime="00:03:30.61" resultid="1799" heatid="4715" lane="0" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:41.28" />
                    <SPLIT distance="150" swimtime="00:02:38.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Żmiejko" birthdate="1963-01-01" gender="M" nation="POL" license="500309700377" athleteid="1784">
              <RESULTS>
                <RESULT eventid="1090" points="630" swimtime="00:00:29.43" resultid="1785" heatid="4612" lane="9" entrytime="00:00:29.85" />
                <RESULT eventid="1124" points="632" swimtime="00:02:45.37" resultid="1786" heatid="4626" lane="4" entrytime="00:02:48.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:02:07.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="708" swimtime="00:01:04.69" resultid="1787" heatid="4671" lane="6" entrytime="00:01:05.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1456" points="701" swimtime="00:00:31.12" resultid="1788" heatid="4702" lane="1" entrytime="00:00:31.45" />
                <RESULT eventid="1490" points="576" swimtime="00:01:19.41" resultid="1789" heatid="4712" lane="9" entrytime="00:01:21.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1633" points="627" swimtime="00:01:12.42" resultid="1790" heatid="4740" lane="7" entrytime="00:01:13.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="599" swimtime="00:00:37.89" resultid="1791" heatid="4760" lane="9" entrytime="00:00:37.85" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00706" nation="POL" region="06" clubid="1800" name="UKS SP8 Chrzanów" shortname="SP8 Chrzanów">
          <ATHLETES>
            <ATHLETE firstname="Alfred" lastname="Zabrzański" birthdate="1954-05-12" gender="M" nation="POL" athleteid="1801">
              <RESULTS>
                <RESULT eventid="1090" points="464" swimtime="00:00:33.85" resultid="1802" heatid="4607" lane="5" entrytime="00:00:34.31" entrycourse="LCM" />
                <RESULT eventid="1182" points="316" swimtime="00:14:43.04" resultid="1803" heatid="4634" lane="8" entrytime="00:13:58.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:02:26.44" />
                    <SPLIT distance="200" swimtime="00:03:23.15" />
                    <SPLIT distance="250" swimtime="00:04:18.84" />
                    <SPLIT distance="300" swimtime="00:05:17.98" />
                    <SPLIT distance="350" swimtime="00:06:15.20" />
                    <SPLIT distance="400" swimtime="00:07:12.85" />
                    <SPLIT distance="450" swimtime="00:08:08.90" />
                    <SPLIT distance="500" swimtime="00:09:03.59" />
                    <SPLIT distance="550" swimtime="00:09:59.92" />
                    <SPLIT distance="600" swimtime="00:10:57.41" />
                    <SPLIT distance="650" swimtime="00:11:53.08" />
                    <SPLIT distance="700" swimtime="00:12:50.68" />
                    <SPLIT distance="750" swimtime="00:13:47.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="1804" heatid="4647" lane="8" entrytime="00:00:44.93" entrycourse="LCM" />
                <RESULT eventid="1320" points="430" swimtime="00:01:18.79" resultid="1805" heatid="4668" lane="2" entrytime="00:01:17.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" status="DNS" swimtime="00:00:00.00" resultid="1806" heatid="4710" lane="2" entrytime="00:01:43.70" entrycourse="LCM" />
                <RESULT eventid="1524" points="321" swimtime="00:03:08.84" resultid="1807" heatid="4721" lane="0" entrytime="00:02:59.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:28.06" />
                    <SPLIT distance="150" swimtime="00:02:19.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="255" swimtime="00:03:58.91" resultid="1808" heatid="4747" lane="6" entrytime="00:03:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.44" />
                    <SPLIT distance="100" swimtime="00:01:57.09" />
                    <SPLIT distance="150" swimtime="00:03:00.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="1809" heatid="4800" lane="3" entrytime="00:06:38.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MALOD" nation="POL" region="05" clubid="2254" name="MASTERS Łódź">
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Grzeszczuk" birthdate="1991-02-25" gender="F" nation="POL" license="503605600035" athleteid="2255">
              <RESULTS>
                <RESULT eventid="1404" points="657" swimtime="00:01:20.61" resultid="2256" heatid="4688" lane="3" entrytime="00:01:18.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="599" swimtime="00:00:32.59" resultid="2257" heatid="4696" lane="4" entrytime="00:00:32.40" />
                <RESULT eventid="1684" points="748" swimtime="00:00:35.48" resultid="2258" heatid="4755" lane="5" entrytime="00:00:35.11" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06306" nation="POL" region="06" clubid="2105" name="KS KORONA 1919 Kraków" shortname="KORONA 1919 Kraków">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Toporski" birthdate="1959-10-20" gender="M" nation="POL" license="506306700060" athleteid="2129">
              <RESULTS>
                <RESULT eventid="1286" points="402" swimtime="00:03:35.99" resultid="2130" heatid="4656" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.41" />
                    <SPLIT distance="100" swimtime="00:01:46.95" />
                    <SPLIT distance="150" swimtime="00:02:42.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="194" swimtime="00:04:07.52" resultid="2131" heatid="4679" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.10" />
                    <SPLIT distance="100" swimtime="00:01:56.95" />
                    <SPLIT distance="150" swimtime="00:03:04.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="358" swimtime="00:01:40.83" resultid="2132" heatid="4690" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="251" swimtime="00:08:08.18" resultid="2133" heatid="4788" lane="9" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.44" />
                    <SPLIT distance="100" swimtime="00:01:57.12" />
                    <SPLIT distance="150" swimtime="00:03:13.67" />
                    <SPLIT distance="200" swimtime="00:04:27.18" />
                    <SPLIT distance="250" swimtime="00:05:28.43" />
                    <SPLIT distance="300" swimtime="00:06:25.88" />
                    <SPLIT distance="350" swimtime="00:07:20.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="163" swimtime="00:01:53.40" resultid="2134" heatid="4738" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="289" swimtime="00:00:48.27" resultid="2135" heatid="4757" lane="1" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariola" lastname="Kuliś" birthdate="1966-07-27" gender="F" nation="POL" license="506306600043" athleteid="2106">
              <RESULTS>
                <RESULT eventid="1059" points="693" swimtime="00:00:31.91" resultid="2107" heatid="4600" lane="6" entrytime="00:00:31.50" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1107" points="586" swimtime="00:03:00.98" resultid="2108" heatid="4620" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:23.37" />
                    <SPLIT distance="150" swimtime="00:02:17.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="590" swimtime="00:00:38.12" resultid="2109" heatid="4642" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1303" points="604" swimtime="00:01:13.37" resultid="2110" heatid="4662" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="673" swimtime="00:01:31.14" resultid="2111" heatid="4687" lane="3" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="734" swimtime="00:00:39.84" resultid="2112" heatid="4754" lane="3" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" license="506306600048" athleteid="2144">
              <RESULTS>
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="2147" heatid="4647" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1107" points="545" swimtime="00:03:21.43" resultid="2591" heatid="4620" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="100" swimtime="00:01:37.59" />
                    <SPLIT distance="150" swimtime="00:02:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1158" points="498" swimtime="00:13:00.27" resultid="2592" heatid="4632" lane="0" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                    <SPLIT distance="100" swimtime="00:01:28.68" />
                    <SPLIT distance="150" swimtime="00:02:16.67" />
                    <SPLIT distance="200" swimtime="00:03:06.48" />
                    <SPLIT distance="250" swimtime="00:03:56.32" />
                    <SPLIT distance="300" swimtime="00:04:46.18" />
                    <SPLIT distance="350" swimtime="00:05:36.40" />
                    <SPLIT distance="400" swimtime="00:06:26.41" />
                    <SPLIT distance="450" swimtime="00:07:15.95" />
                    <SPLIT distance="500" swimtime="00:08:06.05" />
                    <SPLIT distance="550" swimtime="00:08:56.08" />
                    <SPLIT distance="600" swimtime="00:09:45.68" />
                    <SPLIT distance="650" swimtime="00:10:35.53" />
                    <SPLIT distance="700" swimtime="00:11:25.42" />
                    <SPLIT distance="750" swimtime="00:12:14.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="464" swimtime="00:00:43.66" resultid="2593" heatid="4642" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="1337" points="430" swimtime="00:03:33.33" resultid="2594" heatid="4677" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                    <SPLIT distance="100" swimtime="00:01:40.89" />
                    <SPLIT distance="150" swimtime="00:02:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="485" swimtime="00:02:59.40" resultid="2595" heatid="4716" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:26.10" />
                    <SPLIT distance="150" swimtime="00:02:13.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="517" swimtime="00:07:14.67" resultid="2596" heatid="4786" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="100" swimtime="00:01:41.75" />
                    <SPLIT distance="150" swimtime="00:02:40.85" />
                    <SPLIT distance="200" swimtime="00:03:35.81" />
                    <SPLIT distance="250" swimtime="00:04:38.62" />
                    <SPLIT distance="300" swimtime="00:05:41.51" />
                    <SPLIT distance="350" swimtime="00:06:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" status="DNS" swimtime="00:00:00.00" resultid="2597" heatid="4744" lane="5" entrytime="00:03:25.00" />
                <RESULT eventid="1742" status="DNS" swimtime="00:00:00.00" resultid="2598" heatid="4793" lane="4" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Waga" birthdate="1940-07-04" gender="M" nation="POL" license="506306700064" athleteid="2136">
              <RESULTS>
                <RESULT eventid="1090" points="203" swimtime="00:00:54.36" resultid="2137" heatid="4604" lane="4" entrytime="00:00:51.00" />
                <RESULT eventid="1182" points="196" swimtime="00:20:20.52" resultid="2138" heatid="4633" lane="7" entrytime="00:19:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.80" />
                    <SPLIT distance="100" swimtime="00:02:22.93" />
                    <SPLIT distance="150" swimtime="00:03:42.42" />
                    <SPLIT distance="200" swimtime="00:05:00.19" />
                    <SPLIT distance="250" swimtime="00:06:22.45" />
                    <SPLIT distance="300" swimtime="00:07:38.92" />
                    <SPLIT distance="350" swimtime="00:08:55.23" />
                    <SPLIT distance="400" swimtime="00:10:12.51" />
                    <SPLIT distance="450" swimtime="00:11:32.07" />
                    <SPLIT distance="500" swimtime="00:12:47.41" />
                    <SPLIT distance="550" swimtime="00:14:05.80" />
                    <SPLIT distance="600" swimtime="00:15:20.68" />
                    <SPLIT distance="650" swimtime="00:16:38.05" />
                    <SPLIT distance="700" swimtime="00:17:55.13" />
                    <SPLIT distance="750" swimtime="00:19:08.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="193" swimtime="00:02:04.11" resultid="2139" heatid="4665" lane="6" entrytime="00:01:52.00" />
                <RESULT eventid="1422" points="135" swimtime="00:03:03.65" resultid="2140" heatid="4689" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="176" swimtime="00:04:45.89" resultid="2141" heatid="4719" lane="9" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.13" />
                    <SPLIT distance="100" swimtime="00:02:19.30" />
                    <SPLIT distance="150" swimtime="00:03:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="194" swimtime="00:01:11.98" resultid="2142" heatid="4757" lane="0" entrytime="00:01:20.00" />
                <RESULT eventid="1766" points="185" swimtime="00:10:05.65" resultid="2143" heatid="4802" lane="5" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.60" />
                    <SPLIT distance="100" swimtime="00:02:25.14" />
                    <SPLIT distance="150" swimtime="00:03:44.00" />
                    <SPLIT distance="200" swimtime="00:05:05.27" />
                    <SPLIT distance="250" swimtime="00:06:21.20" />
                    <SPLIT distance="300" swimtime="00:07:38.94" />
                    <SPLIT distance="350" swimtime="00:08:54.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogusław" lastname="Kwiatkowski" birthdate="1956-07-24" gender="M" nation="POL" license="506306700044" athleteid="2122">
              <RESULTS>
                <RESULT eventid="1090" points="163" swimtime="00:00:47.95" resultid="2123" heatid="4605" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="1252" points="126" swimtime="00:01:01.60" resultid="2124" heatid="4645" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1320" points="141" swimtime="00:01:54.21" resultid="2125" heatid="4665" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="107" swimtime="00:02:37.12" resultid="2126" heatid="4690" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="140" swimtime="00:04:51.53" resultid="2127" heatid="4746" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.83" />
                    <SPLIT distance="100" swimtime="00:02:18.53" />
                    <SPLIT distance="150" swimtime="00:03:36.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="137" swimtime="00:08:57.39" resultid="2128" heatid="4801" lane="0" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.92" />
                    <SPLIT distance="100" swimtime="00:02:06.29" />
                    <SPLIT distance="150" swimtime="00:03:16.02" />
                    <SPLIT distance="200" swimtime="00:04:25.83" />
                    <SPLIT distance="250" swimtime="00:05:34.61" />
                    <SPLIT distance="300" swimtime="00:06:44.56" />
                    <SPLIT distance="350" swimtime="00:07:52.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Leńczowska" birthdate="1982-01-15" gender="F" nation="POL" license="506306600071" athleteid="2113">
              <RESULTS>
                <RESULT eventid="1059" points="522" swimtime="00:00:32.82" resultid="2114" heatid="4601" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1107" points="524" swimtime="00:02:59.84" resultid="2115" heatid="4620" lane="6" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:24.85" />
                    <SPLIT distance="150" swimtime="00:02:18.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="442" swimtime="00:00:38.86" resultid="2116" heatid="4642" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1303" points="467" swimtime="00:01:14.79" resultid="2117" heatid="4661" lane="1" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="517" swimtime="00:00:35.32" resultid="2118" heatid="4696" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1473" points="412" swimtime="00:01:26.95" resultid="2119" heatid="4708" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="447" swimtime="00:03:07.23" resultid="2120" heatid="4745" lane="1" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                    <SPLIT distance="100" swimtime="00:01:32.27" />
                    <SPLIT distance="150" swimtime="00:02:20.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="427" swimtime="00:00:43.05" resultid="2121" heatid="4753" lane="2" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Baranik" birthdate="1969-06-29" gender="M" nation="POL" license="506306700027" athleteid="3759">
              <RESULTS>
                <RESULT eventid="1090" points="682" swimtime="00:00:27.35" resultid="3760" heatid="4604" lane="8" />
                <RESULT eventid="1320" points="672" swimtime="00:01:01.80" resultid="3761" heatid="4664" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="645" swimtime="00:00:29.94" resultid="3762" heatid="4698" lane="0" />
                <RESULT eventid="1701" points="557" swimtime="00:00:36.33" resultid="3763" heatid="4756" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03311" nation="POL" region="11" clubid="2357" name="UKS WODNIK 29 Katowice" shortname="WODNIK 29 Katowice">
          <ATHLETES>
            <ATHLETE firstname="Jerzy" lastname="Mrożiński" birthdate="1959-12-28" gender="M" nation="POL" athleteid="2358">
              <RESULTS>
                <RESULT eventid="1286" points="547" swimtime="00:03:14.95" resultid="2359" heatid="4657" lane="2" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                    <SPLIT distance="100" swimtime="00:01:33.98" />
                    <SPLIT distance="150" swimtime="00:02:24.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="585" swimtime="00:01:25.62" resultid="2360" heatid="4692" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="2361" heatid="4760" lane="7" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Mróz" birthdate="1979-06-09" gender="F" nation="POL" athleteid="2367">
              <RESULTS>
                <RESULT eventid="1234" points="413" swimtime="00:00:39.77" resultid="2368" heatid="4642" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1303" points="443" swimtime="00:01:16.09" resultid="2369" heatid="4662" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="469" swimtime="00:02:46.31" resultid="2370" heatid="4716" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:03.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="445" swimtime="00:05:44.07" resultid="2371" heatid="4791" lane="9" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:21.38" />
                    <SPLIT distance="150" swimtime="00:02:04.96" />
                    <SPLIT distance="200" swimtime="00:02:49.30" />
                    <SPLIT distance="250" swimtime="00:03:33.38" />
                    <SPLIT distance="300" swimtime="00:04:17.93" />
                    <SPLIT distance="350" swimtime="00:05:01.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Wilczek" birthdate="1958-03-01" gender="M" nation="POL" athleteid="2362">
              <RESULTS>
                <RESULT eventid="1090" points="588" swimtime="00:00:31.27" resultid="2363" heatid="4611" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1320" points="472" swimtime="00:01:16.36" resultid="2364" heatid="4669" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="569" swimtime="00:00:34.24" resultid="2365" heatid="4700" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1633" points="430" swimtime="00:01:27.17" resultid="2366" heatid="4739" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="07611" nation="POL" region="11" clubid="2674" name="UKS DRAGON Sosnowiec" shortname="DRAGON Sosnowiec">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Jankowski" birthdate="1995-01-01" gender="M" nation="POL" athleteid="2673">
              <RESULTS>
                <RESULT eventid="1090" points="728" swimtime="00:00:24.78" resultid="2675" heatid="4617" lane="1" entrytime="00:00:24.50" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1252" points="814" swimtime="00:00:27.24" resultid="2676" heatid="4651" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1320" points="837" swimtime="00:00:53.53" resultid="2677" heatid="4675" lane="6" entrytime="00:00:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="748" swimtime="00:01:00.68" resultid="2678" heatid="4713" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1667" points="465" swimtime="00:02:38.38" resultid="2679" heatid="4750" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.07" />
                    <SPLIT distance="100" swimtime="00:01:12.19" />
                    <SPLIT distance="150" swimtime="00:01:55.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04501" nation="POL" region="01" clubid="2337" name="MKS SWIM ACADEMY Termy Jakuba Oława" shortname="SWIM ACADEMY Oława">
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Chorąży" birthdate="1978-09-27" gender="F" nation="POL" license="104501600044" athleteid="2338">
              <RESULTS>
                <RESULT eventid="1269" status="DNS" swimtime="00:00:00.00" resultid="2339" heatid="4654" lane="0" entrytime="00:03:10.50" />
                <RESULT eventid="1404" points="549" swimtime="00:01:28.32" resultid="2340" heatid="4688" lane="1" entrytime="00:01:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="550" swimtime="00:00:34.65" resultid="2341" heatid="4696" lane="6" entrytime="00:00:33.90" />
                <RESULT eventid="1684" points="648" swimtime="00:00:38.78" resultid="2342" heatid="4755" lane="8" entrytime="00:00:37.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LEWAR" nation="POL" region="14" clubid="3585" name="LEGIA Warszawa" />
        <CLUB type="CLUB" code="MABIA" nation="POL" region="09" clubid="2182" name="MASTERS Białystok">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Twarowski" birthdate="1965-05-24" gender="M" nation="POL" athleteid="2183">
              <RESULTS>
                <RESULT comment="Przekroczony limit czasu" eventid="1216" status="OTL" swimtime="00:27:07.80" resultid="2184" heatid="4638" lane="4" entrytime="00:26:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:42.54" />
                    <SPLIT distance="150" swimtime="00:02:36.54" />
                    <SPLIT distance="200" swimtime="00:03:31.47" />
                    <SPLIT distance="250" swimtime="00:04:26.92" />
                    <SPLIT distance="300" swimtime="00:05:21.45" />
                    <SPLIT distance="350" swimtime="00:06:16.54" />
                    <SPLIT distance="400" swimtime="00:07:11.69" />
                    <SPLIT distance="450" swimtime="00:08:05.29" />
                    <SPLIT distance="500" swimtime="00:09:00.29" />
                    <SPLIT distance="550" swimtime="00:09:53.26" />
                    <SPLIT distance="600" swimtime="00:10:47.63" />
                    <SPLIT distance="650" swimtime="00:11:41.96" />
                    <SPLIT distance="700" swimtime="00:12:37.27" />
                    <SPLIT distance="750" swimtime="00:13:32.27" />
                    <SPLIT distance="800" swimtime="00:14:27.31" />
                    <SPLIT distance="850" swimtime="00:15:20.62" />
                    <SPLIT distance="900" swimtime="00:16:15.37" />
                    <SPLIT distance="950" swimtime="00:17:09.53" />
                    <SPLIT distance="1000" swimtime="00:18:05.17" />
                    <SPLIT distance="1050" swimtime="00:18:59.17" />
                    <SPLIT distance="1100" swimtime="00:19:54.20" />
                    <SPLIT distance="1150" swimtime="00:20:48.43" />
                    <SPLIT distance="1200" swimtime="00:21:44.02" />
                    <SPLIT distance="1250" swimtime="00:22:38.59" />
                    <SPLIT distance="1300" swimtime="00:23:33.95" />
                    <SPLIT distance="1350" swimtime="00:24:27.08" />
                    <SPLIT distance="1400" swimtime="00:25:22.29" />
                    <SPLIT distance="1450" swimtime="00:26:16.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="355" swimtime="00:00:40.99" resultid="2185" heatid="4648" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1490" points="329" swimtime="00:01:31.98" resultid="2186" heatid="4710" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" status="DNS" swimtime="00:00:00.00" resultid="2187" heatid="4720" lane="7" entrytime="00:03:19.00" />
                <RESULT eventid="1667" points="311" swimtime="00:03:27.73" resultid="2188" heatid="4747" lane="4" entrytime="00:03:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.82" />
                    <SPLIT distance="100" swimtime="00:01:42.28" />
                    <SPLIT distance="150" swimtime="00:02:36.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="247" swimtime="00:06:57.94" resultid="2189" heatid="4800" lane="6" entrytime="00:06:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.96" />
                    <SPLIT distance="100" swimtime="00:01:40.82" />
                    <SPLIT distance="150" swimtime="00:02:34.75" />
                    <SPLIT distance="200" swimtime="00:03:29.41" />
                    <SPLIT distance="250" swimtime="00:04:23.98" />
                    <SPLIT distance="300" swimtime="00:05:18.21" />
                    <SPLIT distance="350" swimtime="00:06:10.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZSUW" nation="POL" region="14" clubid="2805" name="KU AZS UW Warszawa" shortname="AZS UW Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Gralewski" birthdate="1994-01-11" gender="M" nation="POL" athleteid="2824">
              <RESULTS>
                <RESULT eventid="1090" points="630" swimtime="00:00:26.01" resultid="2825" heatid="4614" lane="2" entrytime="00:00:27.49" entrycourse="LCM" />
                <RESULT eventid="1124" points="602" swimtime="00:02:26.36" resultid="2826" heatid="4628" lane="7" entrytime="00:02:25.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                    <SPLIT distance="100" swimtime="00:01:08.24" />
                    <SPLIT distance="150" swimtime="00:01:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="731" swimtime="00:00:55.99" resultid="2827" heatid="4673" lane="3" entrytime="00:00:59.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="641" swimtime="00:02:08.40" resultid="2828" heatid="4725" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:01.30" />
                    <SPLIT distance="150" swimtime="00:01:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="547" swimtime="00:01:04.88" resultid="2829" heatid="4742" lane="0" entrytime="00:01:04.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="605" swimtime="00:04:44.86" resultid="2830" heatid="4795" lane="5" entrytime="00:04:29.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="100" swimtime="00:01:06.25" />
                    <SPLIT distance="150" swimtime="00:01:42.22" />
                    <SPLIT distance="200" swimtime="00:02:18.18" />
                    <SPLIT distance="250" swimtime="00:02:54.17" />
                    <SPLIT distance="300" swimtime="00:03:30.43" />
                    <SPLIT distance="350" swimtime="00:04:07.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Szafarczyk" birthdate="1997-06-22" gender="M" nation="POL" athleteid="2811">
              <RESULTS>
                <RESULT eventid="1124" points="687" swimtime="00:02:20.04" resultid="2812" heatid="4628" lane="6" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                    <SPLIT distance="150" swimtime="00:01:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="597" swimtime="00:02:36.49" resultid="2813" heatid="4658" lane="5" entrytime="00:02:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:18.07" />
                    <SPLIT distance="150" swimtime="00:01:57.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="624" swimtime="00:01:10.66" resultid="2814" heatid="4693" lane="8" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="604" swimtime="00:05:19.42" resultid="2815" heatid="4787" lane="4" entrytime="00:04:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:11.84" />
                    <SPLIT distance="150" swimtime="00:01:55.00" />
                    <SPLIT distance="200" swimtime="00:02:37.25" />
                    <SPLIT distance="250" swimtime="00:03:21.04" />
                    <SPLIT distance="300" swimtime="00:04:05.04" />
                    <SPLIT distance="350" swimtime="00:04:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="590" swimtime="00:02:26.36" resultid="2816" heatid="4750" lane="8" entrytime="00:02:32.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:11.62" />
                    <SPLIT distance="150" swimtime="00:01:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="600" swimtime="00:00:32.25" resultid="2817" heatid="4762" lane="8" entrytime="00:00:31.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Kaźmierczak" birthdate="1997-07-06" gender="M" nation="POL" athleteid="2835" />
            <ATHLETE firstname="Eugeniusz" lastname="Puzan" birthdate="1995-06-05" gender="M" nation="POL" athleteid="2831">
              <RESULTS>
                <RESULT eventid="1456" points="697" swimtime="00:00:26.74" resultid="2832" heatid="4705" lane="1" entrytime="00:00:26.00" entrycourse="LCM" />
                <RESULT eventid="1633" points="734" swimtime="00:00:58.85" resultid="2833" heatid="4742" lane="4" entrytime="00:00:58.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="476" swimtime="00:00:34.84" resultid="2834" heatid="4761" lane="0" entrytime="00:00:35.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Mordzonek" birthdate="2001-08-13" gender="M" nation="POL" athleteid="2818">
              <RESULTS>
                <RESULT eventid="1354" swimtime="00:02:44.43" resultid="2819" heatid="4681" lane="7" entrytime="00:02:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:03.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" swimtime="00:02:17.08" resultid="2820" heatid="4724" lane="5" entrytime="00:02:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="150" swimtime="00:01:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" swimtime="00:01:09.76" resultid="2821" heatid="4741" lane="3" entrytime="00:01:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Micorek" birthdate="1993-08-25" gender="M" nation="POL" athleteid="2837">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="2838" heatid="4614" lane="9" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="2839" heatid="4650" lane="2" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2840" heatid="4673" lane="7" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1456" points="588" swimtime="00:00:27.76" resultid="2841" heatid="4703" lane="5" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1633" status="DNS" swimtime="00:00:00.00" resultid="2842" heatid="4742" lane="3" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="2843" heatid="4761" lane="5" entrytime="00:00:33.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rębas" birthdate="1989-12-11" gender="M" nation="POL" athleteid="2806">
              <RESULTS>
                <RESULT eventid="1090" points="624" swimtime="00:00:25.89" resultid="2807" heatid="4613" lane="6" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1320" points="702" swimtime="00:00:56.01" resultid="2808" heatid="4673" lane="2" entrytime="00:00:59.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="655" swimtime="00:00:26.77" resultid="2809" heatid="4704" lane="3" entrytime="00:00:27.05" entrycourse="LCM" />
                <RESULT eventid="1633" points="710" swimtime="00:00:59.51" resultid="2810" heatid="4742" lane="2" entrytime="00:01:00.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Pachowski" birthdate="1997-05-06" gender="M" nation="POL" athleteid="2822">
              <RESULTS>
                <RESULT eventid="1182" points="595" swimtime="00:09:59.54" resultid="2823" heatid="4636" lane="4" entrytime="00:09:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:02.64" />
                    <SPLIT distance="150" swimtime="00:01:38.40" />
                    <SPLIT distance="200" swimtime="00:02:15.04" />
                    <SPLIT distance="250" swimtime="00:02:52.71" />
                    <SPLIT distance="300" swimtime="00:03:30.86" />
                    <SPLIT distance="350" swimtime="00:04:09.72" />
                    <SPLIT distance="400" swimtime="00:04:48.49" />
                    <SPLIT distance="450" swimtime="00:05:27.38" />
                    <SPLIT distance="500" swimtime="00:06:06.62" />
                    <SPLIT distance="550" swimtime="00:06:46.39" />
                    <SPLIT distance="600" swimtime="00:07:25.47" />
                    <SPLIT distance="650" swimtime="00:08:04.38" />
                    <SPLIT distance="700" swimtime="00:08:42.52" />
                    <SPLIT distance="750" swimtime="00:09:21.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="765" swimtime="00:01:40.53" resultid="2836" heatid="4728" lane="4" entrytime="00:01:37.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.12" />
                    <SPLIT distance="100" swimtime="00:00:50.99" />
                    <SPLIT distance="150" swimtime="00:01:15.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2822" number="1" />
                    <RELAYPOSITION athleteid="2837" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="2806" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2831" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NIUK" nation="UKR" clubid="4035" name="Niezrzeszony - Kijów">
          <ATHLETES>
            <ATHLETE firstname="Serhii" lastname="Chernov" birthdate="1950-07-15" gender="M" nation="UKR" athleteid="2102">
              <RESULTS>
                <RESULT eventid="1090" points="117" swimtime="00:00:56.59" resultid="2103" heatid="4604" lane="3" entrytime="00:00:55.97" entrycourse="SCM" />
                <RESULT eventid="1320" points="106" swimtime="00:02:13.50" resultid="2104" heatid="4665" lane="1" entrytime="00:02:14.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="3138" name="WARSAW MASTERS TEAM Warszawa" shortname="WMT Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Leszek" lastname="Rąpała" birthdate="1962-12-05" gender="M" nation="POL" athleteid="3286">
              <RESULTS>
                <RESULT eventid="1456" points="189" swimtime="00:00:48.16" resultid="3287" heatid="4698" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1524" points="191" swimtime="00:03:41.36" resultid="3288" heatid="4719" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.39" />
                    <SPLIT distance="100" swimtime="00:01:45.01" />
                    <SPLIT distance="150" swimtime="00:02:45.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="192" swimtime="00:07:56.47" resultid="3289" heatid="4800" lane="8" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                    <SPLIT distance="100" swimtime="00:01:47.05" />
                    <SPLIT distance="150" swimtime="00:02:48.25" />
                    <SPLIT distance="200" swimtime="00:03:50.64" />
                    <SPLIT distance="250" swimtime="00:04:54.29" />
                    <SPLIT distance="300" swimtime="00:05:58.66" />
                    <SPLIT distance="350" swimtime="00:07:01.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Giejsztowt" birthdate="1978-06-13" gender="M" nation="POL" athleteid="3225">
              <RESULTS>
                <RESULT eventid="1216" points="518" swimtime="00:20:43.51" resultid="3226" heatid="4639" lane="6" entrytime="00:20:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:14.47" />
                    <SPLIT distance="150" swimtime="00:01:54.18" />
                    <SPLIT distance="200" swimtime="00:02:34.30" />
                    <SPLIT distance="250" swimtime="00:03:15.39" />
                    <SPLIT distance="300" swimtime="00:03:56.61" />
                    <SPLIT distance="350" swimtime="00:04:37.14" />
                    <SPLIT distance="400" swimtime="00:05:19.24" />
                    <SPLIT distance="450" swimtime="00:05:59.79" />
                    <SPLIT distance="500" swimtime="00:06:41.38" />
                    <SPLIT distance="550" swimtime="00:07:22.18" />
                    <SPLIT distance="600" swimtime="00:08:04.14" />
                    <SPLIT distance="650" swimtime="00:08:46.59" />
                    <SPLIT distance="700" swimtime="00:09:28.96" />
                    <SPLIT distance="750" swimtime="00:10:11.04" />
                    <SPLIT distance="800" swimtime="00:10:53.63" />
                    <SPLIT distance="850" swimtime="00:11:35.87" />
                    <SPLIT distance="900" swimtime="00:12:19.03" />
                    <SPLIT distance="950" swimtime="00:13:01.17" />
                    <SPLIT distance="1000" swimtime="00:13:43.73" />
                    <SPLIT distance="1050" swimtime="00:14:25.86" />
                    <SPLIT distance="1100" swimtime="00:15:09.25" />
                    <SPLIT distance="1150" swimtime="00:15:52.46" />
                    <SPLIT distance="1200" swimtime="00:16:35.72" />
                    <SPLIT distance="1250" swimtime="00:17:18.56" />
                    <SPLIT distance="1300" swimtime="00:18:00.39" />
                    <SPLIT distance="1350" swimtime="00:18:41.46" />
                    <SPLIT distance="1400" swimtime="00:19:23.40" />
                    <SPLIT distance="1450" swimtime="00:20:05.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="601" swimtime="00:01:01.88" resultid="3227" heatid="4672" lane="2" entrytime="00:01:02.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="569" swimtime="00:00:30.45" resultid="3228" heatid="4702" lane="8" entrytime="00:00:31.50" />
                <RESULT eventid="1524" points="617" swimtime="00:02:18.24" resultid="3229" heatid="4724" lane="0" entrytime="00:02:18.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:07.34" />
                    <SPLIT distance="150" swimtime="00:01:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="586" swimtime="00:05:00.01" resultid="3230" heatid="4796" lane="7" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:49.41" />
                    <SPLIT distance="200" swimtime="00:02:28.12" />
                    <SPLIT distance="250" swimtime="00:03:06.43" />
                    <SPLIT distance="300" swimtime="00:03:45.18" />
                    <SPLIT distance="350" swimtime="00:04:23.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marlena" lastname="Dobrasiewicz" birthdate="1988-05-24" gender="F" nation="POL" athleteid="3277">
              <RESULTS>
                <RESULT eventid="1404" points="546" swimtime="00:01:26.19" resultid="3278" heatid="4687" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="487" swimtime="00:00:39.82" resultid="3279" heatid="4754" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Matlak" birthdate="1984-05-04" gender="F" nation="POL" athleteid="3214">
              <RESULTS>
                <RESULT eventid="1439" points="490" swimtime="00:00:34.81" resultid="3215" heatid="4695" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1507" points="440" swimtime="00:02:45.60" resultid="3216" heatid="4715" lane="4" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:17.39" />
                    <SPLIT distance="150" swimtime="00:02:01.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="461" swimtime="00:05:44.49" resultid="3217" heatid="4792" lane="0" entrytime="00:05:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                    <SPLIT distance="150" swimtime="00:02:03.63" />
                    <SPLIT distance="200" swimtime="00:02:48.43" />
                    <SPLIT distance="250" swimtime="00:03:33.12" />
                    <SPLIT distance="300" swimtime="00:04:18.72" />
                    <SPLIT distance="350" swimtime="00:05:02.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Skośkiewicz" birthdate="1966-05-05" gender="M" nation="POL" athleteid="3184">
              <RESULTS>
                <RESULT eventid="1090" points="643" swimtime="00:00:28.32" resultid="3185" heatid="4612" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1124" points="705" swimtime="00:02:38.04" resultid="3186" heatid="4627" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:02:02.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="646" swimtime="00:00:33.58" resultid="3187" heatid="4650" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1320" points="734" swimtime="00:01:02.06" resultid="3188" heatid="4672" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="640" swimtime="00:00:30.81" resultid="3189" heatid="4703" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1524" points="732" swimtime="00:02:17.57" resultid="3190" heatid="4723" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:07.87" />
                    <SPLIT distance="150" swimtime="00:01:43.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="601" swimtime="00:01:11.73" resultid="3191" heatid="4740" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="599" swimtime="00:05:11.34" resultid="3192" heatid="4796" lane="2" entrytime="00:04:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:13.85" />
                    <SPLIT distance="150" swimtime="00:01:53.44" />
                    <SPLIT distance="200" swimtime="00:02:33.92" />
                    <SPLIT distance="250" swimtime="00:03:13.44" />
                    <SPLIT distance="300" swimtime="00:03:53.28" />
                    <SPLIT distance="350" swimtime="00:04:33.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Mikołajków" birthdate="1992-11-28" gender="M" nation="POL" athleteid="3290">
              <RESULTS>
                <RESULT eventid="1090" points="400" swimtime="00:00:30.03" resultid="3291" heatid="4610" lane="6" entrytime="00:00:30.62" />
                <RESULT eventid="1422" points="402" swimtime="00:01:22.98" resultid="3292" heatid="4690" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="341" swimtime="00:00:33.27" resultid="3293" heatid="4700" lane="7" entrytime="00:00:36.12" />
                <RESULT eventid="1701" points="433" swimtime="00:00:36.65" resultid="3294" heatid="4760" lane="0" entrytime="00:00:37.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" athleteid="3246">
              <RESULTS>
                <RESULT eventid="1090" points="658" swimtime="00:00:27.07" resultid="3247" heatid="4614" lane="7" entrytime="00:00:27.50" />
                <RESULT eventid="1320" points="626" swimtime="00:01:01.04" resultid="3248" heatid="4673" lane="0" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="639" swimtime="00:01:15.17" resultid="3249" heatid="4692" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="590" swimtime="00:00:30.08" resultid="3250" heatid="4702" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1701" points="762" swimtime="00:00:31.99" resultid="3251" heatid="4761" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1766" points="415" swimtime="00:05:36.39" resultid="3252" heatid="4797" lane="9" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                    <SPLIT distance="150" swimtime="00:01:58.90" />
                    <SPLIT distance="200" swimtime="00:02:41.66" />
                    <SPLIT distance="250" swimtime="00:03:25.33" />
                    <SPLIT distance="300" swimtime="00:04:08.99" />
                    <SPLIT distance="350" swimtime="00:04:53.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Rogosz" birthdate="1976-04-28" gender="M" nation="POL" athleteid="3193">
              <RESULTS>
                <RESULT eventid="1090" points="522" swimtime="00:00:29.24" resultid="3194" heatid="4611" lane="4" entrytime="00:00:29.90" />
                <RESULT eventid="1124" points="574" swimtime="00:02:36.49" resultid="3195" heatid="4627" lane="1" entrytime="00:02:40.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:02:01.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="552" swimtime="00:02:49.96" resultid="3196" heatid="4658" lane="9" entrytime="00:02:54.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:23.66" />
                    <SPLIT distance="150" swimtime="00:02:07.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="595" swimtime="00:05:37.27" resultid="3197" heatid="4787" lane="8" entrytime="00:05:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:20.11" />
                    <SPLIT distance="150" swimtime="00:02:05.03" />
                    <SPLIT distance="200" swimtime="00:02:50.95" />
                    <SPLIT distance="250" swimtime="00:03:35.92" />
                    <SPLIT distance="300" swimtime="00:04:22.88" />
                    <SPLIT distance="350" swimtime="00:05:00.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="438" swimtime="00:01:14.83" resultid="3198" heatid="4740" lane="9" entrytime="00:01:17.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="497" swimtime="00:05:16.82" resultid="3199" heatid="4797" lane="1" entrytime="00:05:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                    <SPLIT distance="100" swimtime="00:01:18.63" />
                    <SPLIT distance="150" swimtime="00:01:59.30" />
                    <SPLIT distance="200" swimtime="00:02:40.91" />
                    <SPLIT distance="250" swimtime="00:03:20.87" />
                    <SPLIT distance="300" swimtime="00:04:01.22" />
                    <SPLIT distance="350" swimtime="00:04:39.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leszek" lastname="Madej" birthdate="1960-06-17" gender="M" nation="POL" athleteid="3260">
              <RESULTS>
                <RESULT eventid="1090" points="655" swimtime="00:00:29.04" resultid="3261" heatid="4612" lane="0" entrytime="00:00:29.54" />
                <RESULT eventid="1182" points="639" swimtime="00:10:51.15" resultid="3262" heatid="4635" lane="1" entrytime="00:11:29.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:17.98" />
                    <SPLIT distance="150" swimtime="00:01:59.84" />
                    <SPLIT distance="200" swimtime="00:02:41.47" />
                    <SPLIT distance="250" swimtime="00:03:23.50" />
                    <SPLIT distance="300" swimtime="00:04:05.09" />
                    <SPLIT distance="350" swimtime="00:04:46.63" />
                    <SPLIT distance="400" swimtime="00:05:27.67" />
                    <SPLIT distance="450" swimtime="00:06:08.61" />
                    <SPLIT distance="500" swimtime="00:06:49.71" />
                    <SPLIT distance="550" swimtime="00:07:30.39" />
                    <SPLIT distance="600" swimtime="00:08:11.23" />
                    <SPLIT distance="650" swimtime="00:08:51.67" />
                    <SPLIT distance="700" swimtime="00:09:31.90" />
                    <SPLIT distance="750" swimtime="00:10:11.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="769" swimtime="00:01:02.92" resultid="3263" heatid="4671" lane="4" entrytime="00:01:03.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="602" swimtime="00:01:24.82" resultid="3264" heatid="4692" lane="7" entrytime="00:01:23.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="718" swimtime="00:02:22.54" resultid="3265" heatid="4723" lane="6" entrytime="00:02:21.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:11.61" />
                    <SPLIT distance="150" swimtime="00:01:47.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="625" swimtime="00:00:37.35" resultid="3266" heatid="4760" lane="8" entrytime="00:00:37.11" />
                <RESULT eventid="1766" points="711" swimtime="00:05:07.95" resultid="3267" heatid="4797" lane="5" entrytime="00:05:15.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:01:56.24" />
                    <SPLIT distance="200" swimtime="00:02:36.21" />
                    <SPLIT distance="250" swimtime="00:03:15.36" />
                    <SPLIT distance="300" swimtime="00:03:53.81" />
                    <SPLIT distance="350" swimtime="00:04:31.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Dargas-Miszczak" birthdate="1981-09-06" gender="F" nation="POL" athleteid="3237">
              <RESULTS>
                <RESULT eventid="1059" points="495" swimtime="00:00:33.42" resultid="3238" heatid="4599" lane="4" entrytime="00:00:33.50" />
                <RESULT eventid="1158" points="385" swimtime="00:12:20.36" resultid="3239" heatid="4631" lane="2" entrytime="00:13:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                    <SPLIT distance="150" swimtime="00:02:11.01" />
                    <SPLIT distance="200" swimtime="00:02:57.27" />
                    <SPLIT distance="250" swimtime="00:03:44.70" />
                    <SPLIT distance="300" swimtime="00:04:32.07" />
                    <SPLIT distance="350" swimtime="00:05:18.83" />
                    <SPLIT distance="400" swimtime="00:06:05.62" />
                    <SPLIT distance="450" swimtime="00:06:53.92" />
                    <SPLIT distance="500" swimtime="00:07:41.02" />
                    <SPLIT distance="550" swimtime="00:08:28.65" />
                    <SPLIT distance="600" swimtime="00:09:16.90" />
                    <SPLIT distance="650" swimtime="00:10:02.63" />
                    <SPLIT distance="700" swimtime="00:10:50.41" />
                    <SPLIT distance="750" swimtime="00:11:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="453" swimtime="00:01:15.53" resultid="3240" heatid="4662" lane="9" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1337" points="257" swimtime="00:03:47.70" resultid="3241" heatid="4676" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                    <SPLIT distance="100" swimtime="00:01:45.04" />
                    <SPLIT distance="150" swimtime="00:02:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="470" swimtime="00:00:36.47" resultid="3242" heatid="4696" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1507" points="458" swimtime="00:02:47.63" resultid="3243" heatid="4716" lane="1" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:21.09" />
                    <SPLIT distance="150" swimtime="00:02:05.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="378" swimtime="00:00:44.83" resultid="3244" heatid="4753" lane="3" entrytime="00:00:46.80" />
                <RESULT eventid="1742" points="397" swimtime="00:05:57.44" resultid="3245" heatid="4793" lane="3" entrytime="00:06:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:22.82" />
                    <SPLIT distance="150" swimtime="00:02:08.83" />
                    <SPLIT distance="200" swimtime="00:02:54.39" />
                    <SPLIT distance="250" swimtime="00:03:41.76" />
                    <SPLIT distance="300" swimtime="00:04:28.85" />
                    <SPLIT distance="350" swimtime="00:05:15.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zenon" lastname="Kuliś" birthdate="1954-06-04" gender="M" nation="POL" athleteid="3218">
              <RESULTS>
                <RESULT eventid="1090" points="254" swimtime="00:00:41.34" resultid="3219" heatid="4605" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1182" points="288" swimtime="00:15:10.99" resultid="3220" heatid="4633" lane="3" entrytime="00:15:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.10" />
                    <SPLIT distance="100" swimtime="00:01:46.88" />
                    <SPLIT distance="150" swimtime="00:02:45.19" />
                    <SPLIT distance="200" swimtime="00:03:43.22" />
                    <SPLIT distance="250" swimtime="00:04:42.98" />
                    <SPLIT distance="300" swimtime="00:05:39.56" />
                    <SPLIT distance="350" swimtime="00:06:36.53" />
                    <SPLIT distance="400" swimtime="00:07:34.47" />
                    <SPLIT distance="450" swimtime="00:08:32.71" />
                    <SPLIT distance="500" swimtime="00:09:30.37" />
                    <SPLIT distance="550" swimtime="00:10:27.66" />
                    <SPLIT distance="600" swimtime="00:11:24.62" />
                    <SPLIT distance="650" swimtime="00:12:21.34" />
                    <SPLIT distance="700" swimtime="00:13:18.45" />
                    <SPLIT distance="750" swimtime="00:14:15.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="3221" heatid="4646" lane="2" entrytime="00:00:53.00" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3222" heatid="4666" lane="7" entrytime="00:01:35.00" />
                <RESULT eventid="1524" points="247" swimtime="00:03:25.98" resultid="3223" heatid="4719" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                    <SPLIT distance="100" swimtime="00:01:40.13" />
                    <SPLIT distance="150" swimtime="00:02:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="268" swimtime="00:07:10.46" resultid="3224" heatid="4801" lane="2" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                    <SPLIT distance="100" swimtime="00:01:43.66" />
                    <SPLIT distance="150" swimtime="00:02:39.67" />
                    <SPLIT distance="200" swimtime="00:03:35.00" />
                    <SPLIT distance="250" swimtime="00:04:29.81" />
                    <SPLIT distance="300" swimtime="00:05:24.27" />
                    <SPLIT distance="350" swimtime="00:06:18.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Sołtan" birthdate="1975-12-02" gender="M" nation="POL" athleteid="3273" />
            <ATHLETE firstname="Zbigniew" lastname="Paluszak" birthdate="1967-02-17" gender="M" nation="POL" athleteid="3200">
              <RESULTS>
                <RESULT eventid="1090" points="208" swimtime="00:00:41.26" resultid="3201" heatid="4605" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1124" points="273" swimtime="00:03:36.80" resultid="3202" heatid="4624" lane="1" entrytime="00:03:44.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                    <SPLIT distance="100" swimtime="00:01:43.19" />
                    <SPLIT distance="150" swimtime="00:02:44.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="229" swimtime="00:00:47.41" resultid="3203" heatid="4646" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1320" points="204" swimtime="00:01:35.05" resultid="3204" heatid="4666" lane="5" entrytime="00:01:31.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="214" swimtime="00:00:44.34" resultid="3205" heatid="4698" lane="5" entrytime="00:00:42.58" />
                <RESULT eventid="1524" points="223" swimtime="00:03:24.27" resultid="3206" heatid="4719" lane="6" entrytime="00:03:33.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                    <SPLIT distance="100" swimtime="00:01:40.69" />
                    <SPLIT distance="150" swimtime="00:02:35.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="253" swimtime="00:00:47.42" resultid="3207" heatid="4757" lane="4" entrytime="00:00:48.25" />
                <RESULT eventid="1766" points="227" swimtime="00:07:09.67" resultid="3208" heatid="4801" lane="4" entrytime="00:07:19.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                    <SPLIT distance="100" swimtime="00:01:39.27" />
                    <SPLIT distance="150" swimtime="00:02:33.93" />
                    <SPLIT distance="200" swimtime="00:03:29.48" />
                    <SPLIT distance="250" swimtime="00:04:25.00" />
                    <SPLIT distance="300" swimtime="00:05:20.46" />
                    <SPLIT distance="350" swimtime="00:06:16.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Warchoł" birthdate="1953-08-30" gender="M" nation="POL" athleteid="3295">
              <RESULTS>
                <RESULT eventid="1090" points="612" swimtime="00:00:32.63" resultid="3296" heatid="4610" lane="2" entrytime="00:00:30.95" />
                <RESULT eventid="1124" points="618" swimtime="00:03:11.28" resultid="3297" heatid="4626" lane="9" entrytime="00:02:55.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                    <SPLIT distance="100" swimtime="00:01:30.58" />
                    <SPLIT distance="150" swimtime="00:02:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="702" swimtime="00:01:11.24" resultid="3298" heatid="4670" lane="7" entrytime="00:01:10.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1490" points="700" swimtime="00:01:22.75" resultid="3299" heatid="4711" lane="3" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1667" points="754" swimtime="00:02:56.06" resultid="3300" heatid="4749" lane="8" entrytime="00:02:52.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="100" swimtime="00:01:24.19" />
                    <SPLIT distance="150" swimtime="00:02:10.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Szemberg" birthdate="1949-07-26" gender="F" nation="POL" athleteid="3209">
              <RESULTS>
                <RESULT eventid="1059" points="177" swimtime="00:00:54.64" resultid="3210" heatid="4597" lane="0" entrytime="00:00:56.05" />
                <RESULT eventid="1199" points="260" swimtime="00:34:53.81" resultid="3211" heatid="4637" lane="7" entrytime="00:36:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.95" />
                    <SPLIT distance="100" swimtime="00:02:11.30" />
                    <SPLIT distance="150" swimtime="00:03:21.46" />
                    <SPLIT distance="200" swimtime="00:04:32.63" />
                    <SPLIT distance="250" swimtime="00:05:43.06" />
                    <SPLIT distance="300" swimtime="00:06:53.03" />
                    <SPLIT distance="350" swimtime="00:08:04.20" />
                    <SPLIT distance="400" swimtime="00:09:15.60" />
                    <SPLIT distance="450" swimtime="00:10:24.34" />
                    <SPLIT distance="500" swimtime="00:11:34.19" />
                    <SPLIT distance="550" swimtime="00:12:43.12" />
                    <SPLIT distance="600" swimtime="00:13:52.90" />
                    <SPLIT distance="650" swimtime="00:15:02.00" />
                    <SPLIT distance="700" swimtime="00:16:13.03" />
                    <SPLIT distance="750" swimtime="00:17:23.03" />
                    <SPLIT distance="800" swimtime="00:18:32.86" />
                    <SPLIT distance="850" swimtime="00:19:43.56" />
                    <SPLIT distance="900" swimtime="00:20:52.91" />
                    <SPLIT distance="950" swimtime="00:22:02.63" />
                    <SPLIT distance="1000" swimtime="00:23:12.35" />
                    <SPLIT distance="1050" swimtime="00:24:23.34" />
                    <SPLIT distance="1100" swimtime="00:25:33.17" />
                    <SPLIT distance="1150" swimtime="00:26:45.60" />
                    <SPLIT distance="1200" swimtime="00:27:56.02" />
                    <SPLIT distance="1250" swimtime="00:29:06.84" />
                    <SPLIT distance="1300" swimtime="00:30:17.34" />
                    <SPLIT distance="1350" swimtime="00:31:28.17" />
                    <SPLIT distance="1400" swimtime="00:32:38.43" />
                    <SPLIT distance="1450" swimtime="00:33:48.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="181" swimtime="00:04:24.27" resultid="3212" heatid="4714" lane="3" entrytime="00:04:34.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.84" />
                    <SPLIT distance="100" swimtime="00:02:07.73" />
                    <SPLIT distance="150" swimtime="00:03:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="209" swimtime="00:09:00.85" resultid="3213" heatid="4794" lane="3" entrytime="00:08:59.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.72" />
                    <SPLIT distance="100" swimtime="00:02:09.64" />
                    <SPLIT distance="150" swimtime="00:03:19.72" />
                    <SPLIT distance="200" swimtime="00:04:29.94" />
                    <SPLIT distance="250" swimtime="00:05:38.36" />
                    <SPLIT distance="300" swimtime="00:06:46.91" />
                    <SPLIT distance="350" swimtime="00:07:54.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Bielecka" birthdate="1988-04-07" gender="F" nation="POL" athleteid="3153">
              <RESULTS>
                <RESULT eventid="1107" points="544" swimtime="00:02:52.76" resultid="3154" heatid="4621" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:21.06" />
                    <SPLIT distance="150" swimtime="00:02:10.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1337" points="409" swimtime="00:03:08.77" resultid="3155" heatid="4677" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:29.01" />
                    <SPLIT distance="150" swimtime="00:02:18.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="494" swimtime="00:00:34.73" resultid="3156" heatid="4696" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1573" points="507" swimtime="00:06:15.60" resultid="3157" heatid="4785" lane="7" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:29.34" />
                    <SPLIT distance="150" swimtime="00:02:17.77" />
                    <SPLIT distance="200" swimtime="00:03:04.03" />
                    <SPLIT distance="250" swimtime="00:03:55.46" />
                    <SPLIT distance="300" swimtime="00:04:47.22" />
                    <SPLIT distance="350" swimtime="00:05:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="465" swimtime="00:01:20.07" resultid="3158" heatid="4736" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="494" swimtime="00:00:39.64" resultid="3159" heatid="4754" lane="4" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Kośla" birthdate="1993-01-05" gender="F" nation="POL" athleteid="3179">
              <RESULTS>
                <RESULT eventid="1059" points="555" swimtime="00:00:31.31" resultid="3180" heatid="4601" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1234" points="572" swimtime="00:00:34.40" resultid="3181" heatid="4643" lane="6" entrytime="00:00:33.50" />
                <RESULT eventid="1473" points="565" swimtime="00:01:14.73" resultid="3182" heatid="4708" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="585" swimtime="00:02:44.47" resultid="3183" heatid="4745" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                    <SPLIT distance="100" swimtime="00:01:19.86" />
                    <SPLIT distance="150" swimtime="00:02:02.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Dziedzic" birthdate="1986-01-20" gender="F" nation="POL" athleteid="3139">
              <RESULTS>
                <RESULT eventid="1107" points="440" swimtime="00:03:05.41" resultid="3140" heatid="4618" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:28.23" />
                    <SPLIT distance="150" swimtime="00:02:21.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="457" swimtime="00:11:51.68" resultid="3141" heatid="4632" lane="7" entrytime="00:11:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:19.90" />
                    <SPLIT distance="150" swimtime="00:02:02.78" />
                    <SPLIT distance="200" swimtime="00:02:47.03" />
                    <SPLIT distance="250" swimtime="00:03:31.30" />
                    <SPLIT distance="300" swimtime="00:04:15.87" />
                    <SPLIT distance="350" swimtime="00:05:00.57" />
                    <SPLIT distance="400" swimtime="00:05:45.98" />
                    <SPLIT distance="450" swimtime="00:06:31.99" />
                    <SPLIT distance="500" swimtime="00:07:18.24" />
                    <SPLIT distance="550" swimtime="00:08:04.41" />
                    <SPLIT distance="600" swimtime="00:08:50.63" />
                    <SPLIT distance="650" swimtime="00:09:36.76" />
                    <SPLIT distance="700" swimtime="00:10:22.81" />
                    <SPLIT distance="750" swimtime="00:11:07.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="366" swimtime="00:00:38.37" resultid="3142" heatid="4696" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1650" points="382" swimtime="00:03:10.31" resultid="3143" heatid="4745" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                    <SPLIT distance="100" swimtime="00:01:31.68" />
                    <SPLIT distance="150" swimtime="00:02:21.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="442" swimtime="00:05:49.25" resultid="3144" heatid="4792" lane="6" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:21.39" />
                    <SPLIT distance="150" swimtime="00:02:05.84" />
                    <SPLIT distance="200" swimtime="00:02:50.68" />
                    <SPLIT distance="250" swimtime="00:03:34.92" />
                    <SPLIT distance="300" swimtime="00:04:20.61" />
                    <SPLIT distance="350" swimtime="00:05:05.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olga" lastname="Krysiak" birthdate="1991-06-07" gender="F" nation="POL" athleteid="3231">
              <RESULTS>
                <RESULT eventid="1059" points="617" swimtime="00:00:30.23" resultid="3232" heatid="4601" lane="6" entrytime="00:00:29.50" />
                <RESULT eventid="1158" points="478" swimtime="00:11:13.29" resultid="3233" heatid="4632" lane="2" entrytime="00:10:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:18.30" />
                    <SPLIT distance="150" swimtime="00:02:00.03" />
                    <SPLIT distance="200" swimtime="00:02:42.40" />
                    <SPLIT distance="250" swimtime="00:03:25.70" />
                    <SPLIT distance="300" swimtime="00:04:08.67" />
                    <SPLIT distance="350" swimtime="00:04:52.18" />
                    <SPLIT distance="400" swimtime="00:05:35.78" />
                    <SPLIT distance="450" swimtime="00:06:18.00" />
                    <SPLIT distance="500" swimtime="00:07:01.06" />
                    <SPLIT distance="550" swimtime="00:07:43.99" />
                    <SPLIT distance="600" swimtime="00:08:26.45" />
                    <SPLIT distance="650" swimtime="00:09:09.12" />
                    <SPLIT distance="700" swimtime="00:09:51.91" />
                    <SPLIT distance="750" swimtime="00:10:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="565" swimtime="00:01:06.81" resultid="3234" heatid="4663" lane="8" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="557" swimtime="00:02:28.69" resultid="3235" heatid="4717" lane="7" entrytime="00:02:26.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:12.03" />
                    <SPLIT distance="150" swimtime="00:01:50.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="566" swimtime="00:05:12.65" resultid="3236" heatid="4791" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:14.94" />
                    <SPLIT distance="150" swimtime="00:01:55.30" />
                    <SPLIT distance="200" swimtime="00:02:35.76" />
                    <SPLIT distance="250" swimtime="00:03:15.74" />
                    <SPLIT distance="300" swimtime="00:03:55.74" />
                    <SPLIT distance="350" swimtime="00:04:35.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Porada" birthdate="1983-10-06" gender="M" nation="POL" athleteid="3145">
              <RESULTS>
                <RESULT eventid="1090" points="550" swimtime="00:00:28.30" resultid="3146" heatid="4613" lane="2" entrytime="00:00:28.10" />
                <RESULT eventid="1124" points="581" swimtime="00:02:36.46" resultid="3147" heatid="4628" lane="9" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                    <SPLIT distance="100" swimtime="00:01:16.27" />
                    <SPLIT distance="150" swimtime="00:02:00.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="537" swimtime="00:02:50.43" resultid="3148" heatid="4658" lane="0" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:01:21.69" />
                    <SPLIT distance="150" swimtime="00:02:06.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="528" swimtime="00:01:18.65" resultid="3149" heatid="4693" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="548" swimtime="00:00:29.71" resultid="3150" heatid="4703" lane="7" entrytime="00:00:29.90" />
                <RESULT eventid="1633" points="543" swimtime="00:01:08.83" resultid="3151" heatid="4741" lane="0" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="601" swimtime="00:00:34.16" resultid="3152" heatid="4761" lane="6" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Jarecka-Skorykow" birthdate="1974-01-30" gender="F" nation="POL" athleteid="3274">
              <RESULTS>
                <RESULT eventid="1404" points="426" swimtime="00:01:36.07" resultid="3275" heatid="4686" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="481" swimtime="00:00:42.83" resultid="3276" heatid="4753" lane="1" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Pfitzner" birthdate="1986-05-24" gender="M" nation="POL" athleteid="3268">
              <RESULTS>
                <RESULT eventid="1252" points="478" swimtime="00:00:33.46" resultid="3269" heatid="4650" lane="5" entrytime="00:00:31.80" />
                <RESULT eventid="1320" points="539" swimtime="00:01:02.38" resultid="3270" heatid="4673" lane="6" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" status="DNS" swimtime="00:00:00.00" resultid="3271" heatid="4712" lane="3" entrytime="00:01:12.00" />
                <RESULT eventid="1701" points="448" swimtime="00:00:37.04" resultid="3272" heatid="4759" lane="6" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Saienko" birthdate="1994-08-03" gender="M" nation="POL" athleteid="3160">
              <RESULTS>
                <RESULT eventid="1090" points="626" swimtime="00:00:26.06" resultid="3161" heatid="4615" lane="3" entrytime="00:00:26.01" />
                <RESULT eventid="1320" points="659" swimtime="00:00:57.97" resultid="3162" heatid="4674" lane="2" entrytime="00:00:57.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="581" swimtime="00:00:28.41" resultid="3163" heatid="4704" lane="1" entrytime="00:00:28.01" />
                <RESULT eventid="1633" points="531" swimtime="00:01:05.56" resultid="3164" heatid="4742" lane="8" entrytime="00:01:04.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Burdelak" birthdate="1991-07-06" gender="F" nation="POL" athleteid="3174">
              <RESULTS>
                <RESULT eventid="1059" points="664" swimtime="00:00:29.50" resultid="3175" heatid="4602" lane="1" entrytime="00:00:28.60" />
                <RESULT eventid="1269" points="472" swimtime="00:03:11.19" resultid="3176" heatid="4654" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                    <SPLIT distance="100" swimtime="00:01:33.64" />
                    <SPLIT distance="150" swimtime="00:02:23.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="628" swimtime="00:01:21.84" resultid="3177" heatid="4688" lane="6" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="649" swimtime="00:00:37.21" resultid="3178" heatid="4755" lane="7" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Nowak" birthdate="1952-12-17" gender="M" nation="POL" athleteid="3280">
              <RESULTS>
                <RESULT eventid="1124" points="495" swimtime="00:03:25.89" resultid="3281" heatid="4625" lane="8" entrytime="00:03:28.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                    <SPLIT distance="100" swimtime="00:01:42.64" />
                    <SPLIT distance="150" swimtime="00:02:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="646" swimtime="00:03:33.76" resultid="3282" heatid="4656" lane="4" entrytime="00:03:32.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.08" />
                    <SPLIT distance="100" swimtime="00:01:41.44" />
                    <SPLIT distance="150" swimtime="00:02:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="698" swimtime="00:01:32.40" resultid="3283" heatid="4691" lane="6" entrytime="00:01:31.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="436" swimtime="00:07:49.24" resultid="3284" heatid="4789" lane="6" entrytime="00:08:02.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.81" />
                    <SPLIT distance="100" swimtime="00:01:59.82" />
                    <SPLIT distance="200" swimtime="00:04:03.28" />
                    <SPLIT distance="250" swimtime="00:05:04.22" />
                    <SPLIT distance="300" swimtime="00:06:07.44" />
                    <SPLIT distance="350" swimtime="00:06:59.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="760" swimtime="00:00:39.67" resultid="3285" heatid="4759" lane="2" entrytime="00:00:39.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szymańśki" birthdate="1981-11-04" gender="M" nation="POL" athleteid="3165">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="3166" heatid="4612" lane="4" entrytime="00:00:28.50" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="3167" heatid="4626" lane="7" entrytime="00:02:50.00" />
                <RESULT eventid="1252" points="500" swimtime="00:00:34.16" resultid="3168" heatid="4649" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1320" points="453" swimtime="00:01:06.63" resultid="3169" heatid="4670" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="495" swimtime="00:00:30.73" resultid="3170" heatid="4702" lane="3" entrytime="00:00:30.50" />
                <RESULT eventid="1490" status="DNS" swimtime="00:00:00.00" resultid="3171" heatid="4712" lane="0" entrytime="00:01:20.00" />
                <RESULT eventid="1633" status="DNS" swimtime="00:00:00.00" resultid="3172" heatid="4740" lane="0" entrytime="00:01:16.00" />
                <RESULT eventid="1667" status="DNS" swimtime="00:00:00.00" resultid="3173" heatid="4749" lane="9" entrytime="00:02:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Petryszyn" birthdate="1994-07-31" gender="F" nation="POL" athleteid="3253">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="3254" heatid="4602" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1234" points="569" swimtime="00:00:34.26" resultid="3255" heatid="4643" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1303" points="623" swimtime="00:01:06.67" resultid="3256" heatid="4663" lane="2" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="571" swimtime="00:00:31.71" resultid="3257" heatid="4697" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1473" points="530" swimtime="00:01:16.11" resultid="3258" heatid="4708" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="483" swimtime="00:02:49.65" resultid="3259" heatid="4745" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:01:24.20" />
                    <SPLIT distance="150" swimtime="00:02:07.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="564" swimtime="00:02:03.81" resultid="3305" heatid="4684" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:07.88" />
                    <SPLIT distance="150" swimtime="00:01:36.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3165" number="1" />
                    <RELAYPOSITION athleteid="3246" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="3160" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="3268" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="709" swimtime="00:01:46.43" resultid="3308" heatid="4728" lane="7" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                    <SPLIT distance="100" swimtime="00:00:53.44" />
                    <SPLIT distance="150" swimtime="00:01:18.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3246" number="1" />
                    <RELAYPOSITION athleteid="3273" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="3160" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3268" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1565" points="403" swimtime="00:02:08.45" resultid="3309" heatid="4727" lane="5" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="100" swimtime="00:00:57.58" />
                    <SPLIT distance="150" swimtime="00:01:40.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3165" number="1" />
                    <RELAYPOSITION athleteid="3290" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="3200" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="3145" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1371" points="782" swimtime="00:02:12.79" resultid="3303" heatid="4682" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:43.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3179" number="1" />
                    <RELAYPOSITION athleteid="3174" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3253" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="3231" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1541" points="770" swimtime="00:01:58.95" resultid="3306" heatid="4726" lane="4" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                    <SPLIT distance="100" swimtime="00:00:58.60" />
                    <SPLIT distance="150" swimtime="00:01:28.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3231" number="1" />
                    <RELAYPOSITION athleteid="3253" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="3179" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="3174" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1371" points="577" swimtime="00:02:26.88" resultid="3304" heatid="4682" lane="3" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:01:53.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3153" number="1" />
                    <RELAYPOSITION athleteid="3277" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3139" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="3237" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1541" points="529" swimtime="00:02:14.07" resultid="3307" heatid="4726" lane="3" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:05.59" />
                    <SPLIT distance="150" swimtime="00:01:39.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3214" number="1" />
                    <RELAYPOSITION athleteid="3277" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="3274" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3139" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1141" points="723" swimtime="00:01:51.54" resultid="3301" heatid="4630" lane="5" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                    <SPLIT distance="100" swimtime="00:00:52.82" />
                    <SPLIT distance="150" swimtime="00:01:22.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3160" number="1" />
                    <RELAYPOSITION athleteid="3246" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3231" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3174" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1718" points="566" swimtime="00:02:25.03" resultid="3310" heatid="4765" lane="8" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:14.08" />
                    <SPLIT distance="150" swimtime="00:01:50.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3184" number="1" />
                    <RELAYPOSITION athleteid="3280" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="3237" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3274" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1141" points="622" swimtime="00:01:59.77" resultid="3302" heatid="4630" lane="2" entrytime="00:02:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.23" />
                    <SPLIT distance="150" swimtime="00:01:29.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3273" number="1" />
                    <RELAYPOSITION athleteid="3237" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3193" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3179" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1718" points="713" swimtime="00:02:03.95" resultid="3311" heatid="4765" lane="6" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:06.93" />
                    <SPLIT distance="150" swimtime="00:01:34.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3253" number="1" />
                    <RELAYPOSITION athleteid="3246" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="3160" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3174" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1718" points="592" swimtime="00:02:11.90" resultid="3312" heatid="4765" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:09.35" />
                    <SPLIT distance="150" swimtime="00:01:43.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3179" number="1" />
                    <RELAYPOSITION athleteid="3145" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3153" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3268" number="4" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1718" points="553" swimtime="00:02:17.92" resultid="3313" heatid="4765" lane="1" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:16.18" />
                    <SPLIT distance="150" swimtime="00:01:46.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3139" number="1" />
                    <RELAYPOSITION athleteid="3193" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3273" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3277" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="06711" nation="POL" region="11" clubid="3892" name="UKS  DRAGON Będzin" shortname="DRAGON Będzin">
          <ATHLETES>
            <ATHLETE firstname="Emil" lastname="Strumiński" birthdate="1988-05-18" gender="M" nation="POL" license="306711700032" athleteid="3893">
              <RESULTS>
                <RESULT eventid="1090" points="660" swimtime="00:00:26.13" resultid="3894" heatid="4615" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="1124" points="605" swimtime="00:02:28.49" resultid="3895" heatid="4627" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                    <SPLIT distance="150" swimtime="00:01:57.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="711" swimtime="00:00:56.87" resultid="3896" heatid="4674" lane="4" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="471" swimtime="00:02:37.44" resultid="3897" heatid="4681" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                    <SPLIT distance="150" swimtime="00:01:54.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="672" swimtime="00:00:27.55" resultid="3898" heatid="4704" lane="6" entrytime="00:00:27.50" />
                <RESULT eventid="1524" points="656" swimtime="00:02:09.85" resultid="3899" heatid="4725" lane="1" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:04.01" />
                    <SPLIT distance="150" swimtime="00:01:38.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="623" swimtime="00:01:02.80" resultid="3900" heatid="4742" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="641" swimtime="00:04:45.18" resultid="3901" heatid="4802" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="100" swimtime="00:01:07.75" />
                    <SPLIT distance="150" swimtime="00:01:44.54" />
                    <SPLIT distance="200" swimtime="00:02:22.04" />
                    <SPLIT distance="250" swimtime="00:02:59.45" />
                    <SPLIT distance="300" swimtime="00:03:36.77" />
                    <SPLIT distance="350" swimtime="00:04:12.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00111" nation="POL" region="11" clubid="2343" name="UKS TRÓJKA Częstochowa" shortname="TRÓJKA Częstochowa">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Gajda" birthdate="1995-04-23" gender="M" nation="POL" license="100111700062" athleteid="3962">
              <RESULTS>
                <RESULT eventid="1090" points="701" swimtime="00:00:25.10" resultid="3963" heatid="4616" lane="5" entrytime="00:00:24.98" />
                <RESULT eventid="1182" points="622" swimtime="00:09:50.75" resultid="3964" heatid="4636" lane="6" entrytime="00:09:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:08.56" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                    <SPLIT distance="200" swimtime="00:02:24.01" />
                    <SPLIT distance="250" swimtime="00:03:02.30" />
                    <SPLIT distance="300" swimtime="00:03:40.75" />
                    <SPLIT distance="350" swimtime="00:04:19.29" />
                    <SPLIT distance="400" swimtime="00:04:57.57" />
                    <SPLIT distance="450" swimtime="00:05:30.73" />
                    <SPLIT distance="500" swimtime="00:06:14.44" />
                    <SPLIT distance="550" swimtime="00:06:52.22" />
                    <SPLIT distance="600" swimtime="00:07:29.75" />
                    <SPLIT distance="650" swimtime="00:08:06.23" />
                    <SPLIT distance="700" swimtime="00:08:42.59" />
                    <SPLIT distance="750" swimtime="00:09:17.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="702" swimtime="00:00:56.75" resultid="3965" heatid="4675" lane="1" entrytime="00:00:55.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="533" swimtime="00:02:28.88" resultid="3966" heatid="4681" lane="5" entrytime="00:02:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="150" swimtime="00:01:48.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="694" swimtime="00:00:26.77" resultid="3967" heatid="4705" lane="8" entrytime="00:00:26.30" />
                <RESULT eventid="1524" points="629" swimtime="00:02:09.25" resultid="3968" heatid="4725" lane="6" entrytime="00:02:06.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:03.11" />
                    <SPLIT distance="150" swimtime="00:01:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="670" swimtime="00:01:00.66" resultid="3969" heatid="4742" lane="6" entrytime="00:01:00.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="630" swimtime="00:04:41.07" resultid="3970" heatid="4795" lane="7" entrytime="00:04:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:05.65" />
                    <SPLIT distance="150" swimtime="00:01:41.98" />
                    <SPLIT distance="200" swimtime="00:02:18.98" />
                    <SPLIT distance="250" swimtime="00:02:55.77" />
                    <SPLIT distance="300" swimtime="00:03:32.09" />
                    <SPLIT distance="350" swimtime="00:04:08.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Szczypiński" birthdate="1990-11-28" gender="M" nation="POL" athleteid="2344">
              <RESULTS>
                <RESULT eventid="1090" points="373" swimtime="00:00:30.73" resultid="2345" heatid="4613" lane="0" entrytime="00:00:28.47" />
                <RESULT eventid="1124" points="343" swimtime="00:02:54.53" resultid="2346" heatid="4627" lane="4" entrytime="00:02:38.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:18.11" />
                    <SPLIT distance="150" swimtime="00:02:11.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="378" swimtime="00:00:35.91" resultid="2347" heatid="4650" lane="1" entrytime="00:00:32.90" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2348" heatid="4671" lane="5" entrytime="00:01:04.25" />
                <RESULT eventid="1456" points="365" swimtime="00:00:32.54" resultid="2349" heatid="4702" lane="0" entrytime="00:00:31.69" />
                <RESULT eventid="1490" points="346" swimtime="00:01:19.61" resultid="2350" heatid="4712" lane="4" entrytime="00:01:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" status="DNS" swimtime="00:00:00.00" resultid="2351" heatid="4750" lane="9" entrytime="00:02:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Musik" birthdate="1997-08-04" gender="F" nation="POL" license="100111600053" athleteid="3955">
              <RESULTS>
                <RESULT eventid="1059" points="750" swimtime="00:00:27.97" resultid="3956" heatid="4602" lane="2" entrytime="00:00:28.40" />
                <RESULT eventid="1107" points="741" swimtime="00:02:35.48" resultid="3957" heatid="4621" lane="3" entrytime="00:02:36.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:59.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="790" swimtime="00:01:01.61" resultid="3958" heatid="4663" lane="3" entrytime="00:01:01.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1337" points="543" swimtime="00:02:45.41" resultid="3959" heatid="4677" lane="5" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:02:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="625" swimtime="00:00:30.78" resultid="3960" heatid="4697" lane="8" entrytime="00:00:30.40" />
                <RESULT eventid="1507" points="688" swimtime="00:02:21.06" resultid="3961" heatid="4717" lane="3" entrytime="00:02:18.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:07.23" />
                    <SPLIT distance="150" swimtime="00:01:44.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sonia" lastname="Nowak" birthdate="1996-05-23" gender="F" nation="POL" license="100111600092" athleteid="3946">
              <RESULTS>
                <RESULT eventid="1059" points="520" swimtime="00:00:31.61" resultid="3947" heatid="4600" lane="7" entrytime="00:00:32.20" />
                <RESULT eventid="1158" points="545" swimtime="00:10:43.43" resultid="3948" heatid="4632" lane="5" entrytime="00:10:22.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:16.66" />
                    <SPLIT distance="150" swimtime="00:01:57.09" />
                    <SPLIT distance="200" swimtime="00:02:37.44" />
                    <SPLIT distance="250" swimtime="00:03:17.95" />
                    <SPLIT distance="300" swimtime="00:03:58.51" />
                    <SPLIT distance="350" swimtime="00:04:39.21" />
                    <SPLIT distance="400" swimtime="00:05:19.79" />
                    <SPLIT distance="450" swimtime="00:06:00.20" />
                    <SPLIT distance="500" swimtime="00:06:40.92" />
                    <SPLIT distance="550" swimtime="00:07:21.82" />
                    <SPLIT distance="600" swimtime="00:08:02.75" />
                    <SPLIT distance="650" swimtime="00:08:43.54" />
                    <SPLIT distance="700" swimtime="00:09:24.08" />
                    <SPLIT distance="750" swimtime="00:10:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="604" swimtime="00:01:07.37" resultid="3949" heatid="4663" lane="7" entrytime="00:01:06.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1337" points="538" swimtime="00:02:46.00" resultid="3950" heatid="4677" lane="3" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:19.80" />
                    <SPLIT distance="150" swimtime="00:02:02.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="473" swimtime="00:00:33.76" resultid="3951" heatid="4696" lane="3" entrytime="00:00:33.89" />
                <RESULT eventid="1507" points="619" swimtime="00:02:26.13" resultid="3952" heatid="4717" lane="1" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="520" swimtime="00:01:14.60" resultid="3953" heatid="4736" lane="3" entrytime="00:01:12.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="568" swimtime="00:05:12.20" resultid="3954" heatid="4791" lane="2" entrytime="00:05:08.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:17.11" />
                    <SPLIT distance="150" swimtime="00:01:56.93" />
                    <SPLIT distance="200" swimtime="00:02:36.32" />
                    <SPLIT distance="250" swimtime="00:03:15.65" />
                    <SPLIT distance="300" swimtime="00:03:54.98" />
                    <SPLIT distance="350" swimtime="00:04:34.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Warwas" birthdate="1995-07-13" gender="M" nation="POL" license="100111700100" athleteid="3980">
              <RESULTS>
                <RESULT eventid="1090" points="663" swimtime="00:00:25.57" resultid="3981" heatid="4616" lane="6" entrytime="00:00:25.50" />
                <RESULT comment="Przekroczony limit czasu" eventid="1182" status="OTL" swimtime="00:11:16.93" resultid="3982" heatid="4636" lane="8" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="100" swimtime="00:01:09.59" />
                    <SPLIT distance="150" swimtime="00:01:48.16" />
                    <SPLIT distance="200" swimtime="00:02:27.39" />
                    <SPLIT distance="250" swimtime="00:03:08.11" />
                    <SPLIT distance="300" swimtime="00:03:49.71" />
                    <SPLIT distance="350" swimtime="00:04:31.98" />
                    <SPLIT distance="400" swimtime="00:05:15.58" />
                    <SPLIT distance="450" swimtime="00:05:59.58" />
                    <SPLIT distance="500" swimtime="00:06:44.43" />
                    <SPLIT distance="550" swimtime="00:07:29.36" />
                    <SPLIT distance="600" swimtime="00:08:15.28" />
                    <SPLIT distance="650" swimtime="00:09:00.51" />
                    <SPLIT distance="700" swimtime="00:09:46.28" />
                    <SPLIT distance="750" swimtime="00:10:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="541" swimtime="00:00:31.21" resultid="3983" heatid="4650" lane="3" entrytime="00:00:31.90" />
                <RESULT eventid="1320" points="687" swimtime="00:00:57.16" resultid="3984" heatid="4674" lane="1" entrytime="00:00:58.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="609" swimtime="00:00:27.96" resultid="3985" heatid="4704" lane="7" entrytime="00:00:27.66" />
                <RESULT eventid="1490" points="506" swimtime="00:01:09.09" resultid="3986" heatid="4713" lane="7" entrytime="00:01:06.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" status="DNS" swimtime="00:00:00.00" resultid="3987" heatid="4742" lane="9" entrytime="00:01:04.50" />
                <RESULT eventid="1667" status="DNS" swimtime="00:00:00.00" resultid="3988" heatid="4750" lane="5" entrytime="00:02:19.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kurek" birthdate="1994-07-11" gender="M" nation="POL" license="100111700097" athleteid="3971">
              <RESULTS>
                <RESULT eventid="1090" points="484" swimtime="00:00:28.40" resultid="3972" heatid="4614" lane="1" entrytime="00:00:27.70" />
                <RESULT comment="Przekroczony limit czasu" eventid="1182" status="OTL" swimtime="00:11:20.35" resultid="3973" heatid="4636" lane="0" entrytime="00:10:40.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:14.21" />
                    <SPLIT distance="150" swimtime="00:01:55.05" />
                    <SPLIT distance="200" swimtime="00:02:37.33" />
                    <SPLIT distance="250" swimtime="00:03:19.96" />
                    <SPLIT distance="300" swimtime="00:04:03.79" />
                    <SPLIT distance="350" swimtime="00:04:47.69" />
                    <SPLIT distance="400" swimtime="00:05:31.91" />
                    <SPLIT distance="450" swimtime="00:06:16.70" />
                    <SPLIT distance="500" swimtime="00:07:01.89" />
                    <SPLIT distance="550" swimtime="00:07:46.35" />
                    <SPLIT distance="600" swimtime="00:08:31.20" />
                    <SPLIT distance="650" swimtime="00:09:14.85" />
                    <SPLIT distance="700" swimtime="00:09:58.16" />
                    <SPLIT distance="750" swimtime="00:10:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="389" swimtime="00:03:00.48" resultid="3974" heatid="4658" lane="1" entrytime="00:02:40.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                    <SPLIT distance="150" swimtime="00:02:12.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="483" swimtime="00:01:04.27" resultid="3975" heatid="4672" lane="7" entrytime="00:01:02.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="394" swimtime="00:00:32.32" resultid="3976" heatid="4701" lane="4" entrytime="00:00:32.44" />
                <RESULT eventid="1524" points="436" swimtime="00:02:25.96" resultid="3977" heatid="4724" lane="8" entrytime="00:02:18.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:10.58" />
                    <SPLIT distance="150" swimtime="00:01:48.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="406" swimtime="00:00:36.73" resultid="3978" heatid="4761" lane="9" entrytime="00:00:35.50" />
                <RESULT eventid="1766" points="374" swimtime="00:05:34.29" resultid="3979" heatid="4796" lane="9" entrytime="00:05:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:14.68" />
                    <SPLIT distance="150" swimtime="00:01:55.73" />
                    <SPLIT distance="200" swimtime="00:02:38.68" />
                    <SPLIT distance="250" swimtime="00:03:23.03" />
                    <SPLIT distance="300" swimtime="00:04:08.08" />
                    <SPLIT distance="350" swimtime="00:04:53.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="528" swimtime="00:02:05.92" resultid="4038" heatid="4683" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:40.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2344" number="1" />
                    <RELAYPOSITION athleteid="3971" number="2" reactiontime="+24" />
                    <RELAYPOSITION athleteid="3962" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="3980" number="4" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="600" swimtime="00:01:48.97" resultid="4039" heatid="4727" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                    <SPLIT distance="100" swimtime="00:00:58.69" />
                    <SPLIT distance="150" swimtime="00:01:24.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3971" number="1" />
                    <RELAYPOSITION athleteid="2344" number="2" reactiontime="+9" />
                    <RELAYPOSITION athleteid="3980" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3962" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1141" points="814" swimtime="00:01:48.36" resultid="4037" heatid="4629" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.58" />
                    <SPLIT distance="100" swimtime="00:00:55.97" />
                    <SPLIT distance="150" swimtime="00:01:23.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3980" number="1" />
                    <RELAYPOSITION athleteid="3946" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3955" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="3962" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="14814" nation="POL" region="14" clubid="3865" name="St. Pływackie LEGIA Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Bogdan" lastname="Dubiński" birthdate="1953-05-05" gender="M" nation="POL" license="514814700003" athleteid="3866">
              <RESULTS>
                <RESULT eventid="1090" points="500" swimtime="00:00:34.89" resultid="3867" heatid="4603" lane="5" />
                <RESULT eventid="1182" points="393" swimtime="00:14:30.41" resultid="3868" heatid="4633" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.49" />
                    <SPLIT distance="100" swimtime="00:01:33.70" />
                    <SPLIT distance="150" swimtime="00:02:28.22" />
                    <SPLIT distance="200" swimtime="00:03:23.68" />
                    <SPLIT distance="250" swimtime="00:04:18.92" />
                    <SPLIT distance="300" swimtime="00:05:15.86" />
                    <SPLIT distance="350" swimtime="00:06:12.18" />
                    <SPLIT distance="400" swimtime="00:07:09.64" />
                    <SPLIT distance="450" swimtime="00:08:05.40" />
                    <SPLIT distance="500" swimtime="00:09:02.06" />
                    <SPLIT distance="550" swimtime="00:09:57.90" />
                    <SPLIT distance="600" swimtime="00:10:53.96" />
                    <SPLIT distance="650" swimtime="00:11:49.40" />
                    <SPLIT distance="700" swimtime="00:12:45.52" />
                    <SPLIT distance="750" swimtime="00:13:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="443" swimtime="00:00:44.05" resultid="3869" heatid="4644" lane="4" />
                <RESULT eventid="1320" points="491" swimtime="00:01:20.22" resultid="3870" heatid="4664" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="434" swimtime="00:03:09.17" resultid="3871" heatid="4718" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:27.02" />
                    <SPLIT distance="150" swimtime="00:02:18.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" status="DNS" swimtime="00:00:00.00" resultid="3872" heatid="4790" lane="3" />
                <RESULT eventid="1766" points="399" swimtime="00:06:52.33" resultid="3873" heatid="4802" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:01:32.86" />
                    <SPLIT distance="150" swimtime="00:02:25.50" />
                    <SPLIT distance="200" swimtime="00:03:18.61" />
                    <SPLIT distance="250" swimtime="00:04:15.46" />
                    <SPLIT distance="300" swimtime="00:05:09.15" />
                    <SPLIT distance="350" swimtime="00:06:02.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Certa" birthdate="1993-03-23" gender="F" nation="POL" athleteid="3586">
              <RESULTS>
                <RESULT eventid="1439" points="773" swimtime="00:00:29.94" resultid="3587" heatid="4696" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1615" points="575" swimtime="00:01:10.69" resultid="3588" heatid="4736" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Grzelak" birthdate="1970-06-24" gender="M" nation="POL" license="514814700011" athleteid="3874">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="3875" heatid="4603" lane="3" />
                <RESULT eventid="1124" points="249" swimtime="00:03:28.32" resultid="3876" heatid="4622" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:43.11" />
                    <SPLIT distance="150" swimtime="00:02:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3877" heatid="4665" lane="9" />
                <RESULT eventid="1354" points="240" swimtime="00:03:34.15" resultid="3878" heatid="4678" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                    <SPLIT distance="100" swimtime="00:01:41.93" />
                    <SPLIT distance="150" swimtime="00:02:38.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" status="DNS" swimtime="00:00:00.00" resultid="3879" heatid="4718" lane="7" />
                <RESULT eventid="1597" points="260" swimtime="00:07:26.98" resultid="3880" heatid="4790" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:37.55" />
                    <SPLIT distance="150" swimtime="00:02:44.75" />
                    <SPLIT distance="200" swimtime="00:03:53.25" />
                    <SPLIT distance="250" swimtime="00:04:52.96" />
                    <SPLIT distance="300" swimtime="00:05:54.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="267" swimtime="00:01:28.78" resultid="3881" heatid="4737" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="330" swimtime="00:06:10.29" resultid="3882" heatid="4802" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:02:14.97" />
                    <SPLIT distance="200" swimtime="00:03:02.88" />
                    <SPLIT distance="250" swimtime="00:03:51.48" />
                    <SPLIT distance="300" swimtime="00:04:40.50" />
                    <SPLIT distance="350" swimtime="00:05:27.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Urbańska" birthdate="1992-03-04" gender="F" nation="POL" athleteid="3589">
              <RESULTS>
                <RESULT eventid="1107" points="580" swimtime="00:02:40.52" resultid="3590" heatid="4621" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:15.85" />
                    <SPLIT distance="150" swimtime="00:02:02.55" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1234" points="682" swimtime="00:00:32.45" resultid="3591" heatid="4643" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1404" points="606" swimtime="00:01:22.80" resultid="3592" heatid="4687" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="590" swimtime="00:01:13.65" resultid="3593" heatid="4707" lane="4" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="570" swimtime="00:00:38.85" resultid="3594" heatid="4754" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X">
              <RESULTS>
                <RESULT eventid="1718" points="479" swimtime="00:02:24.67" resultid="5400" heatid="4764" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:01:21.65" />
                    <SPLIT distance="150" swimtime="00:01:51.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3866" number="1" />
                    <RELAYPOSITION athleteid="3586" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="3589" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3874" number="4" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01709" nation="POL" region="09" clubid="2859" name="iSWIM Białystok">
          <ATHLETES>
            <ATHLETE firstname="Dawid" lastname="Perkowski" birthdate="1996-06-10" gender="M" nation="POL" license="117/09700023" athleteid="2871">
              <RESULTS>
                <RESULT eventid="1090" points="596" swimtime="00:00:26.49" resultid="2872" heatid="4615" lane="6" entrytime="00:00:26.20" />
                <RESULT eventid="1320" points="668" swimtime="00:00:57.70" resultid="2873" heatid="4674" lane="8" entrytime="00:00:58.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Gawryluk" birthdate="1953-10-13" gender="M" nation="POL" license="501709700264" athleteid="2863">
              <RESULTS>
                <RESULT eventid="1090" points="177" swimtime="00:00:49.27" resultid="2864" heatid="4605" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1320" points="144" swimtime="00:02:00.75" resultid="2865" heatid="4665" lane="4" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="239" swimtime="00:02:11.92" resultid="2866" heatid="4690" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="202" swimtime="00:01:01.70" resultid="2867" heatid="4757" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="2868" heatid="4802" lane="4" entrytime="00:09:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Iwaniuk-Mróz" birthdate="1979-07-17" gender="F" nation="POL" license="117/09600024" athleteid="2883">
              <RESULTS>
                <RESULT eventid="1059" points="581" swimtime="00:00:31.67" resultid="2884" heatid="4600" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1303" points="521" swimtime="00:01:12.09" resultid="2885" heatid="4662" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="572" swimtime="00:00:34.15" resultid="2886" heatid="4696" lane="2" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Uściłko" birthdate="1995-07-13" gender="M" nation="POL" license="101709700260" athleteid="2869">
              <RESULTS>
                <RESULT eventid="1524" points="702" swimtime="00:02:04.58" resultid="2870" heatid="4725" lane="3" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                    <SPLIT distance="100" swimtime="00:01:01.01" />
                    <SPLIT distance="150" swimtime="00:01:33.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Daszuta" birthdate="1973-03-12" gender="M" nation="POL" license="117/09700012" athleteid="2860">
              <RESULTS>
                <RESULT eventid="1456" status="DNS" swimtime="00:00:00.00" resultid="2861" heatid="4703" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="2862" heatid="4761" lane="1" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Świderski" birthdate="1979-02-13" gender="M" nation="POL" license="517/09700108" athleteid="2881">
              <RESULTS>
                <RESULT eventid="1456" points="551" swimtime="00:00:29.66" resultid="2882" heatid="4702" lane="6" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elżbieta" lastname="Piwowarczyk" birthdate="1966-01-06" gender="F" nation="POL" license="501709600257" athleteid="2874">
              <RESULTS>
                <RESULT eventid="1059" points="494" swimtime="00:00:35.73" resultid="2875" heatid="4599" lane="8" entrytime="00:00:34.90" />
                <RESULT eventid="1234" points="402" swimtime="00:00:43.33" resultid="2876" heatid="4641" lane="3" entrytime="00:00:44.80" />
                <RESULT eventid="1303" points="482" swimtime="00:01:19.05" resultid="2877" heatid="4660" lane="4" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="414" swimtime="00:01:33.47" resultid="2878" heatid="4707" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="457" swimtime="00:02:56.86" resultid="2879" heatid="4715" lane="2" entrytime="00:02:56.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="419" swimtime="00:03:22.69" resultid="2880" heatid="4744" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.44" />
                    <SPLIT distance="100" swimtime="00:01:37.91" />
                    <SPLIT distance="150" swimtime="00:02:31.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" status="DNS" swimtime="00:00:00.00" resultid="2887" heatid="4684" lane="3" entrytime="00:01:57.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2860" number="1" />
                    <RELAYPOSITION athleteid="2871" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2881" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2869" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" status="DNS" swimtime="00:00:00.00" resultid="2888" heatid="4728" lane="3" entrytime="00:01:45.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2860" number="1" />
                    <RELAYPOSITION athleteid="2871" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2869" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2881" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="BM469" nation="POL" region="08" clubid="2288" name="ORION TEAM Rzeszów">
          <ATHLETES>
            <ATHLETE firstname="Mariusz" lastname="Faff" birthdate="1963-11-15" gender="M" nation="POL" license="bm862" athleteid="2289">
              <RESULTS>
                <RESULT eventid="1090" points="619" swimtime="00:00:29.60" resultid="2290" heatid="4611" lane="5" entrytime="00:00:29.94" />
                <RESULT eventid="1766" points="526" swimtime="00:05:40.49" resultid="2291" heatid="4798" lane="4" entrytime="00:05:32.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:18.51" />
                    <SPLIT distance="150" swimtime="00:02:03.46" />
                    <SPLIT distance="200" swimtime="00:02:48.59" />
                    <SPLIT distance="250" swimtime="00:03:32.70" />
                    <SPLIT distance="300" swimtime="00:04:17.64" />
                    <SPLIT distance="350" swimtime="00:05:01.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="491" swimtime="00:02:41.74" resultid="2292" heatid="4722" lane="1" entrytime="00:02:37.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:16.81" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="623" swimtime="00:00:32.36" resultid="2293" heatid="4701" lane="0" entrytime="00:00:33.79" />
                <RESULT eventid="1320" points="631" swimtime="00:01:07.22" resultid="2294" heatid="4671" lane="1" entrytime="00:01:07.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Sarna" birthdate="1975-10-31" gender="M" nation="POL" license="bm842" athleteid="2295">
              <RESULTS>
                <RESULT eventid="1766" points="589" swimtime="00:04:59.38" resultid="2296" heatid="4795" lane="1" entrytime="00:04:43.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:09.05" />
                    <SPLIT distance="150" swimtime="00:01:46.73" />
                    <SPLIT distance="200" swimtime="00:02:25.17" />
                    <SPLIT distance="250" swimtime="00:03:04.24" />
                    <SPLIT distance="300" swimtime="00:03:43.30" />
                    <SPLIT distance="350" swimtime="00:04:22.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="629" swimtime="00:02:17.37" resultid="2297" heatid="4724" lane="4" entrytime="00:02:13.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:07.07" />
                    <SPLIT distance="150" swimtime="00:01:43.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="599" swimtime="00:01:01.95" resultid="2298" heatid="4673" lane="1" entrytime="00:01:00.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="551" swimtime="00:02:38.59" resultid="2299" heatid="4622" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:10.94" />
                    <SPLIT distance="150" swimtime="00:02:00.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="604" swimtime="00:00:27.85" resultid="2300" heatid="4614" lane="3" entrytime="00:00:27.41" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="3842" name="MKS ASTORIA Bydgoszcz" shortname="ASTORIA Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" license="102202700126" athleteid="3843">
              <RESULTS>
                <RESULT eventid="1252" points="197" swimtime="00:00:49.08" resultid="3844" heatid="4645" lane="6" />
                <RESULT eventid="1490" points="160" swimtime="00:01:53.35" resultid="3845" heatid="4709" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="169" swimtime="00:04:03.03" resultid="3846" heatid="4746" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.99" />
                    <SPLIT distance="100" swimtime="00:01:58.45" />
                    <SPLIT distance="150" swimtime="00:03:00.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Krasicki" birthdate="1995-02-17" gender="M" nation="POL" license="102202700140" athleteid="3847">
              <RESULTS>
                <RESULT eventid="1252" points="579" swimtime="00:00:30.51" resultid="3848" heatid="4645" lane="7" />
                <RESULT eventid="1524" points="605" swimtime="00:02:10.90" resultid="3849" heatid="4718" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="100" swimtime="00:01:02.82" />
                    <SPLIT distance="150" swimtime="00:01:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="596" swimtime="00:04:46.31" resultid="3850" heatid="4802" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:05.91" />
                    <SPLIT distance="150" swimtime="00:01:42.46" />
                    <SPLIT distance="200" swimtime="00:02:19.44" />
                    <SPLIT distance="250" swimtime="00:02:56.76" />
                    <SPLIT distance="300" swimtime="00:03:34.15" />
                    <SPLIT distance="350" swimtime="00:04:11.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="IKKON" nation="POL" region="14" clubid="2844" name="IKS Konstancin">
          <ATHLETES>
            <ATHLETE firstname="Rafal" lastname="Juchno" birthdate="1976-10-03" gender="M" nation="POL" license="103714700079" athleteid="2845">
              <RESULTS>
                <RESULT eventid="1090" points="484" swimtime="00:00:29.98" resultid="2846" heatid="4611" lane="1" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1182" points="292" swimtime="00:13:04.50" resultid="2847" heatid="4635" lane="0" entrytime="00:12:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:23.45" />
                    <SPLIT distance="150" swimtime="00:02:11.29" />
                    <SPLIT distance="200" swimtime="00:03:01.26" />
                    <SPLIT distance="250" swimtime="00:03:51.15" />
                    <SPLIT distance="300" swimtime="00:04:42.14" />
                    <SPLIT distance="350" swimtime="00:05:33.19" />
                    <SPLIT distance="400" swimtime="00:06:24.47" />
                    <SPLIT distance="450" swimtime="00:07:16.04" />
                    <SPLIT distance="500" swimtime="00:08:07.26" />
                    <SPLIT distance="550" swimtime="00:08:58.63" />
                    <SPLIT distance="600" swimtime="00:09:49.54" />
                    <SPLIT distance="650" swimtime="00:10:40.26" />
                    <SPLIT distance="700" swimtime="00:11:29.91" />
                    <SPLIT distance="750" swimtime="00:12:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="368" swimtime="00:00:40.74" resultid="2848" heatid="4759" lane="8" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1766" points="341" swimtime="00:05:59.33" resultid="2849" heatid="4798" lane="0" entrytime="00:05:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:18.42" />
                    <SPLIT distance="150" swimtime="00:02:04.36" />
                    <SPLIT distance="200" swimtime="00:02:52.78" />
                    <SPLIT distance="250" swimtime="00:03:40.79" />
                    <SPLIT distance="300" swimtime="00:04:29.67" />
                    <SPLIT distance="350" swimtime="00:05:17.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Obiedziński" birthdate="1969-04-11" gender="M" nation="POL" athleteid="2850">
              <RESULTS>
                <RESULT eventid="1090" points="570" swimtime="00:00:29.04" resultid="2851" heatid="4612" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1124" points="477" swimtime="00:02:47.77" resultid="2852" heatid="4627" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:02:09.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="628" swimtime="00:01:03.21" resultid="2853" heatid="4672" lane="0" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="335" swimtime="00:03:11.84" resultid="2854" heatid="4680" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:28.03" />
                    <SPLIT distance="150" swimtime="00:02:17.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="554" swimtime="00:00:31.51" resultid="2855" heatid="4701" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1524" points="571" swimtime="00:02:22.93" resultid="2856" heatid="4724" lane="7" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:07.58" />
                    <SPLIT distance="150" swimtime="00:01:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="414" swimtime="00:01:16.76" resultid="2857" heatid="4740" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="521" swimtime="00:05:17.98" resultid="2858" heatid="4796" lane="0" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:12.95" />
                    <SPLIT distance="150" swimtime="00:01:53.47" />
                    <SPLIT distance="200" swimtime="00:02:34.43" />
                    <SPLIT distance="250" swimtime="00:03:15.36" />
                    <SPLIT distance="300" swimtime="00:03:56.72" />
                    <SPLIT distance="350" swimtime="00:04:38.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="08" clubid="1871" name="UKS DELFIN MASTERS Tarnobrzeg" shortname="DELFIN MASTERS Tarnobrzeg">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Ślęczka" birthdate="1974-10-23" gender="M" nation="POL" license="500408700205" athleteid="1872">
              <RESULTS>
                <RESULT eventid="1090" points="602" swimtime="00:00:27.89" resultid="1873" heatid="4611" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1124" points="566" swimtime="00:02:37.18" resultid="1874" heatid="4627" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:59.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="589" swimtime="00:01:02.29" resultid="1875" heatid="4671" lane="7" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="561" swimtime="00:01:18.51" resultid="1876" heatid="4692" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="623" swimtime="00:02:17.82" resultid="1877" heatid="4723" lane="5" entrytime="00:02:20.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:06.34" />
                    <SPLIT distance="150" swimtime="00:01:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="520" swimtime="00:01:10.69" resultid="1878" heatid="4740" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="586" swimtime="00:00:34.91" resultid="1879" heatid="4760" lane="5" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TORLT" nation="LTU" clubid="4036" name="Marijampoles TORPEDOS">
          <ATHLETES>
            <ATHLETE firstname="Stasys" lastname="Grigas" birthdate="1941-01-01" gender="M" nation="LTU" athleteid="3612">
              <RESULTS>
                <RESULT eventid="1090" points="140" swimtime="00:01:01.44" resultid="3613" heatid="4604" lane="6" entrytime="00:01:08.24" />
                <RESULT comment="O2 - Pływak nie miał kontaktu ze ścianą podczas nawrotu" eventid="1182" status="DSQ" swimtime="00:00:00.00" resultid="3614" heatid="4633" lane="1" entrytime="00:22:10.00" />
                <RESULT eventid="1252" points="148" swimtime="00:01:12.07" resultid="3615" heatid="4645" lane="3" entrytime="00:01:16.85" />
                <RESULT eventid="1320" points="96" swimtime="00:02:36.54" resultid="3616" heatid="4665" lane="8" entrytime="00:02:49.45" />
                <RESULT eventid="1490" points="162" swimtime="00:02:38.29" resultid="3617" heatid="4709" lane="2" entrytime="00:02:41.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="85" swimtime="00:06:04.34" resultid="3618" heatid="4718" lane="3" entrytime="00:06:09.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.29" />
                    <SPLIT distance="100" swimtime="00:02:56.42" />
                    <SPLIT distance="150" swimtime="00:04:33.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="156" swimtime="00:05:57.80" resultid="3619" heatid="4746" lane="3" entrytime="00:06:12.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.45" />
                    <SPLIT distance="100" swimtime="00:02:57.18" />
                    <SPLIT distance="150" swimtime="00:04:30.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="88" swimtime="00:12:55.18" resultid="3620" heatid="4802" lane="6" entrytime="00:12:13.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vilmantas" lastname="Krasauskas" birthdate="1964-01-01" gender="M" nation="LTU" athleteid="3621">
              <RESULTS>
                <RESULT eventid="1090" points="534" swimtime="00:00:30.13" resultid="3622" heatid="4611" lane="0" entrytime="00:00:30.02" />
                <RESULT eventid="1182" points="538" swimtime="00:11:03.68" resultid="3623" heatid="4635" lane="5" entrytime="00:11:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:01.65" />
                    <SPLIT distance="200" swimtime="00:02:43.82" />
                    <SPLIT distance="250" swimtime="00:03:26.08" />
                    <SPLIT distance="300" swimtime="00:04:08.22" />
                    <SPLIT distance="350" swimtime="00:04:50.37" />
                    <SPLIT distance="400" swimtime="00:05:32.71" />
                    <SPLIT distance="450" swimtime="00:06:14.74" />
                    <SPLIT distance="500" swimtime="00:06:56.94" />
                    <SPLIT distance="550" swimtime="00:07:38.93" />
                    <SPLIT distance="600" swimtime="00:08:21.05" />
                    <SPLIT distance="650" swimtime="00:09:02.91" />
                    <SPLIT distance="700" swimtime="00:09:45.15" />
                    <SPLIT distance="750" swimtime="00:10:26.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="619" swimtime="00:01:05.69" resultid="3624" heatid="4671" lane="2" entrytime="00:01:05.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="604" swimtime="00:02:26.68" resultid="3625" heatid="4723" lane="9" entrytime="00:02:26.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:11.88" />
                    <SPLIT distance="150" swimtime="00:01:49.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="574" swimtime="00:05:15.80" resultid="3626" heatid="4797" lane="6" entrytime="00:05:18.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="150" swimtime="00:01:56.54" />
                    <SPLIT distance="200" swimtime="00:02:37.28" />
                    <SPLIT distance="250" swimtime="00:03:17.49" />
                    <SPLIT distance="300" swimtime="00:03:58.08" />
                    <SPLIT distance="350" swimtime="00:04:37.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="07914" nation="POL" region="14" clubid="1843" name="St. Pł. SWIMMERS Warszawa" shortname="SWIMMERS Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Remigiusz" lastname="Gołębiowski" birthdate="1976-07-07" gender="M" nation="POL" license="507914700017" athleteid="1844">
              <RESULTS>
                <RESULT eventid="1090" points="638" swimtime="00:00:27.35" resultid="1845" heatid="4613" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1182" points="515" swimtime="00:10:49.70" resultid="1846" heatid="4636" lane="5" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:09.78" />
                    <SPLIT distance="150" swimtime="00:01:47.81" />
                    <SPLIT distance="200" swimtime="00:02:26.72" />
                    <SPLIT distance="250" swimtime="00:03:06.37" />
                    <SPLIT distance="300" swimtime="00:03:45.85" />
                    <SPLIT distance="350" swimtime="00:04:26.04" />
                    <SPLIT distance="400" swimtime="00:05:06.38" />
                    <SPLIT distance="450" swimtime="00:05:48.35" />
                    <SPLIT distance="500" swimtime="00:06:32.10" />
                    <SPLIT distance="550" swimtime="00:07:15.10" />
                    <SPLIT distance="600" swimtime="00:07:57.72" />
                    <SPLIT distance="650" swimtime="00:08:40.81" />
                    <SPLIT distance="700" swimtime="00:09:24.51" />
                    <SPLIT distance="750" swimtime="00:10:07.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="630" swimtime="00:01:00.92" resultid="1847" heatid="4674" lane="9" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="649" swimtime="00:00:29.15" resultid="1848" heatid="4702" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1524" points="601" swimtime="00:02:19.49" resultid="1849" heatid="4724" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:08.83" />
                    <SPLIT distance="150" swimtime="00:01:45.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="562" swimtime="00:05:04.20" resultid="1850" heatid="4796" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:12.46" />
                    <SPLIT distance="150" swimtime="00:01:51.70" />
                    <SPLIT distance="200" swimtime="00:02:31.01" />
                    <SPLIT distance="250" swimtime="00:03:10.18" />
                    <SPLIT distance="300" swimtime="00:03:49.02" />
                    <SPLIT distance="350" swimtime="00:04:27.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Lis" birthdate="1979-01-23" gender="M" nation="POL" license="507914700028" athleteid="1851">
              <RESULTS>
                <RESULT eventid="1090" points="432" swimtime="00:00:30.68" resultid="1852" heatid="4610" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="1456" points="358" swimtime="00:00:34.23" resultid="1853" heatid="4700" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1524" points="354" swimtime="00:02:40.65" resultid="1854" heatid="4721" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:16.97" />
                    <SPLIT distance="150" swimtime="00:02:00.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="395" swimtime="00:00:39.30" resultid="1855" heatid="4759" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1766" points="330" swimtime="00:05:57.01" resultid="1856" heatid="4798" lane="8" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:23.05" />
                    <SPLIT distance="150" swimtime="00:02:08.10" />
                    <SPLIT distance="200" swimtime="00:02:54.28" />
                    <SPLIT distance="250" swimtime="00:03:41.09" />
                    <SPLIT distance="300" swimtime="00:04:27.91" />
                    <SPLIT distance="350" swimtime="00:05:14.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01012" nation="POL" region="12" clubid="3851" name="MOSiR Ostrowiec Św.">
          <ATHLETES>
            <ATHLETE firstname="Józef" lastname="Różalski" birthdate="1945-03-28" gender="M" nation="POL" license="501012700001" athleteid="3852">
              <RESULTS>
                <RESULT eventid="1090" points="339" swimtime="00:00:41.85" resultid="3853" heatid="4603" lane="4" />
                <RESULT comment="Przekroczony limit czasu" eventid="1182" status="OTL" swimtime="00:20:12.68" resultid="3854" heatid="4633" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.48" />
                    <SPLIT distance="100" swimtime="00:02:09.63" />
                    <SPLIT distance="150" swimtime="00:03:25.04" />
                    <SPLIT distance="200" swimtime="00:04:43.44" />
                    <SPLIT distance="250" swimtime="00:06:01.49" />
                    <SPLIT distance="300" swimtime="00:07:20.72" />
                    <SPLIT distance="350" swimtime="00:08:39.03" />
                    <SPLIT distance="400" swimtime="00:09:58.66" />
                    <SPLIT distance="450" swimtime="00:11:16.62" />
                    <SPLIT distance="500" swimtime="00:12:35.57" />
                    <SPLIT distance="550" swimtime="00:13:53.68" />
                    <SPLIT distance="600" swimtime="00:15:11.87" />
                    <SPLIT distance="650" swimtime="00:16:27.55" />
                    <SPLIT distance="700" swimtime="00:17:44.22" />
                    <SPLIT distance="750" swimtime="00:19:00.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="198" swimtime="00:00:59.06" resultid="3855" heatid="4645" lane="2" />
                <RESULT eventid="1320" points="228" swimtime="00:01:48.55" resultid="3856" heatid="4664" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="173" swimtime="00:04:21.23" resultid="3857" heatid="4720" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.24" />
                    <SPLIT distance="150" swimtime="00:03:13.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="170" swimtime="00:09:32.59" resultid="3858" heatid="4802" lane="0">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:09.34" />
                    <SPLIT distance="150" swimtime="00:03:22.62" />
                    <SPLIT distance="200" swimtime="00:04:36.14" />
                    <SPLIT distance="250" swimtime="00:05:50.36" />
                    <SPLIT distance="300" swimtime="00:07:07.02" />
                    <SPLIT distance="350" swimtime="00:08:21.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NOTU" nation="GER" clubid="2328" name="NORDER TURNVEREIN Von 1861">
          <ATHLETES>
            <ATHLETE firstname="Katarzyna" lastname="Szwagiel" birthdate="1976-03-14" gender="F" nation="GER" athleteid="2329">
              <RESULTS>
                <RESULT eventid="1107" points="513" swimtime="00:02:56.52" resultid="2330" heatid="4620" lane="4" entrytime="00:02:54.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:26.63" />
                    <SPLIT distance="150" swimtime="00:02:15.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="465" swimtime="00:11:51.63" resultid="2331" heatid="4632" lane="1" entrytime="00:11:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:21.78" />
                    <SPLIT distance="150" swimtime="00:02:06.41" />
                    <SPLIT distance="200" swimtime="00:02:51.61" />
                    <SPLIT distance="250" swimtime="00:03:36.42" />
                    <SPLIT distance="300" swimtime="00:04:21.24" />
                    <SPLIT distance="350" swimtime="00:05:05.90" />
                    <SPLIT distance="400" swimtime="00:05:51.09" />
                    <SPLIT distance="450" swimtime="00:06:36.21" />
                    <SPLIT distance="500" swimtime="00:07:21.31" />
                    <SPLIT distance="550" swimtime="00:08:07.16" />
                    <SPLIT distance="600" swimtime="00:08:53.15" />
                    <SPLIT distance="650" swimtime="00:09:37.92" />
                    <SPLIT distance="700" swimtime="00:10:23.21" />
                    <SPLIT distance="750" swimtime="00:11:08.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="619" swimtime="00:03:12.07" resultid="2332" heatid="4654" lane="1" entrytime="00:03:08.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                    <SPLIT distance="100" swimtime="00:01:33.45" />
                    <SPLIT distance="150" swimtime="00:02:23.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1337" points="405" swimtime="00:03:15.09" resultid="2333" heatid="4677" lane="2" entrytime="00:03:11.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:01:32.59" />
                    <SPLIT distance="150" swimtime="00:02:24.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="471" swimtime="00:01:32.97" resultid="2334" heatid="4687" lane="5" entrytime="00:01:30.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="510" swimtime="00:06:32.71" resultid="2335" heatid="4785" lane="6" entrytime="00:06:11.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:32.15" />
                    <SPLIT distance="150" swimtime="00:02:24.54" />
                    <SPLIT distance="200" swimtime="00:03:15.60" />
                    <SPLIT distance="250" swimtime="00:04:07.24" />
                    <SPLIT distance="300" swimtime="00:04:59.61" />
                    <SPLIT distance="350" swimtime="00:05:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="475" swimtime="00:05:48.50" resultid="2336" heatid="4792" lane="4" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:22.50" />
                    <SPLIT distance="150" swimtime="00:02:06.59" />
                    <SPLIT distance="200" swimtime="00:02:51.09" />
                    <SPLIT distance="250" swimtime="00:03:35.52" />
                    <SPLIT distance="300" swimtime="00:04:20.75" />
                    <SPLIT distance="350" swimtime="00:05:05.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMSZC" nation="POL" region="16" clubid="3040" name="SMT Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Stępień-Gielo" birthdate="1961-05-03" gender="F" nation="POL" athleteid="3102">
              <RESULTS>
                <RESULT eventid="1059" points="479" swimtime="00:00:36.93" resultid="3103" heatid="4598" lane="2" entrytime="00:00:38.70" />
                <RESULT eventid="1158" points="326" swimtime="00:14:58.93" resultid="3104" heatid="4631" lane="1" entrytime="00:15:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.17" />
                    <SPLIT distance="100" swimtime="00:01:42.88" />
                    <SPLIT distance="150" swimtime="00:02:38.54" />
                    <SPLIT distance="200" swimtime="00:03:33.93" />
                    <SPLIT distance="250" swimtime="00:04:30.56" />
                    <SPLIT distance="300" swimtime="00:05:27.40" />
                    <SPLIT distance="350" swimtime="00:06:24.78" />
                    <SPLIT distance="400" swimtime="00:07:22.09" />
                    <SPLIT distance="450" swimtime="00:08:19.49" />
                    <SPLIT distance="500" swimtime="00:09:16.37" />
                    <SPLIT distance="550" swimtime="00:10:13.42" />
                    <SPLIT distance="600" swimtime="00:11:10.75" />
                    <SPLIT distance="650" swimtime="00:12:09.62" />
                    <SPLIT distance="700" swimtime="00:13:07.06" />
                    <SPLIT distance="750" swimtime="00:14:04.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="367" swimtime="00:00:47.21" resultid="3105" heatid="4641" lane="1" entrytime="00:00:48.50" />
                <RESULT eventid="1269" points="505" swimtime="00:03:51.17" resultid="3106" heatid="4653" lane="8" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.36" />
                    <SPLIT distance="100" swimtime="00:01:50.28" />
                    <SPLIT distance="150" swimtime="00:02:50.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="522" swimtime="00:01:43.14" resultid="3107" heatid="4687" lane="9" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="306" swimtime="00:01:50.18" resultid="3108" heatid="4707" lane="9" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="290" swimtime="00:04:03.79" resultid="3109" heatid="4744" lane="1" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.55" />
                    <SPLIT distance="100" swimtime="00:02:02.04" />
                    <SPLIT distance="150" swimtime="00:03:04.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="569" swimtime="00:00:45.16" resultid="3110" heatid="4753" lane="5" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Zając" birthdate="1966-06-30" gender="M" nation="POL" athleteid="3049">
              <RESULTS>
                <RESULT eventid="1090" points="456" swimtime="00:00:31.75" resultid="3050" heatid="4610" lane="9" entrytime="00:00:31.18" />
                <RESULT eventid="1320" points="419" swimtime="00:01:14.83" resultid="3051" heatid="4669" lane="9" entrytime="00:01:15.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="442" swimtime="00:00:34.86" resultid="3052" heatid="4700" lane="4" entrytime="00:00:34.28" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rachel" lastname="Jankowski" birthdate="1999-09-21" gender="F" nation="POL" athleteid="3084">
              <RESULTS>
                <RESULT eventid="1107" swimtime="00:03:07.02" resultid="3085" heatid="4620" lane="0" entrytime="00:03:10.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                    <SPLIT distance="100" swimtime="00:01:35.18" />
                    <SPLIT distance="150" swimtime="00:02:24.47" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Przekroczony limit czasu" eventid="1158" status="OTL" swimtime="00:12:47.12" resultid="3086" heatid="4632" lane="8" entrytime="00:12:02.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="100" swimtime="00:01:23.27" />
                    <SPLIT distance="150" swimtime="00:02:09.57" />
                    <SPLIT distance="200" swimtime="00:02:57.24" />
                    <SPLIT distance="250" swimtime="00:03:45.40" />
                    <SPLIT distance="300" swimtime="00:04:34.18" />
                    <SPLIT distance="350" swimtime="00:05:22.99" />
                    <SPLIT distance="400" swimtime="00:06:12.25" />
                    <SPLIT distance="450" swimtime="00:07:01.66" />
                    <SPLIT distance="500" swimtime="00:07:51.63" />
                    <SPLIT distance="550" swimtime="00:08:41.33" />
                    <SPLIT distance="600" swimtime="00:09:31.72" />
                    <SPLIT distance="650" swimtime="00:10:21.51" />
                    <SPLIT distance="700" swimtime="00:11:11.45" />
                    <SPLIT distance="750" swimtime="00:12:00.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" swimtime="00:03:17.56" resultid="3087" heatid="4653" lane="5" entrytime="00:03:17.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:32.08" />
                    <SPLIT distance="150" swimtime="00:02:22.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" swimtime="00:02:49.19" resultid="3088" heatid="4716" lane="5" entrytime="00:02:40.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:03.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" swimtime="00:06:04.08" resultid="3089" heatid="4792" lane="7" entrytime="00:05:50.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:10.62" />
                    <SPLIT distance="200" swimtime="00:02:57.89" />
                    <SPLIT distance="250" swimtime="00:03:45.37" />
                    <SPLIT distance="300" swimtime="00:04:32.75" />
                    <SPLIT distance="350" swimtime="00:05:18.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iwona" lastname="Damljanović-Wacławik" birthdate="1965-04-21" gender="F" nation="POL" athleteid="3076">
              <RESULTS>
                <RESULT eventid="1107" points="378" swimtime="00:03:29.41" resultid="3077" heatid="4619" lane="6" entrytime="00:03:35.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:40.12" />
                    <SPLIT distance="150" swimtime="00:02:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="362" swimtime="00:13:39.99" resultid="3078" heatid="4631" lane="7" entrytime="00:14:04.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                    <SPLIT distance="100" swimtime="00:01:34.31" />
                    <SPLIT distance="150" swimtime="00:02:25.92" />
                    <SPLIT distance="200" swimtime="00:03:17.70" />
                    <SPLIT distance="250" swimtime="00:04:10.00" />
                    <SPLIT distance="300" swimtime="00:05:01.63" />
                    <SPLIT distance="350" swimtime="00:05:53.70" />
                    <SPLIT distance="400" swimtime="00:06:45.82" />
                    <SPLIT distance="450" swimtime="00:07:37.65" />
                    <SPLIT distance="500" swimtime="00:08:29.29" />
                    <SPLIT distance="550" swimtime="00:09:21.29" />
                    <SPLIT distance="600" swimtime="00:10:13.20" />
                    <SPLIT distance="650" swimtime="00:11:05.68" />
                    <SPLIT distance="700" swimtime="00:11:57.74" />
                    <SPLIT distance="750" swimtime="00:12:49.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="515" swimtime="00:03:42.98" resultid="3079" heatid="4653" lane="1" entrytime="00:03:48.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.47" />
                    <SPLIT distance="100" swimtime="00:01:49.03" />
                    <SPLIT distance="150" swimtime="00:02:47.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="440" swimtime="00:01:45.01" resultid="3080" heatid="4687" lane="0" entrytime="00:01:43.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="409" swimtime="00:00:41.11" resultid="3081" heatid="4695" lane="0" entrytime="00:00:42.07" />
                <RESULT eventid="1615" points="243" swimtime="00:01:50.13" resultid="3082" heatid="4735" lane="3" entrytime="00:01:44.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="443" swimtime="00:00:47.14" resultid="3083" heatid="4753" lane="6" entrytime="00:00:46.86" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Zieliński" birthdate="1992-09-02" gender="M" nation="POL" athleteid="3064">
              <RESULTS>
                <RESULT eventid="1090" points="713" swimtime="00:00:24.77" resultid="3065" heatid="4617" lane="9" entrytime="00:00:24.78" />
                <RESULT eventid="1456" points="620" swimtime="00:00:27.27" resultid="3066" heatid="4705" lane="0" entrytime="00:00:26.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Kramek" birthdate="1992-02-04" gender="M" nation="POL" athleteid="3041">
              <RESULTS>
                <RESULT eventid="1090" points="672" swimtime="00:00:25.26" resultid="3042" heatid="4615" lane="1" entrytime="00:00:26.42" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3043" heatid="4674" lane="0" entrytime="00:00:58.83" />
                <RESULT eventid="1456" points="567" swimtime="00:00:28.10" resultid="3044" heatid="4703" lane="4" entrytime="00:00:28.91" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Szponder" birthdate="1970-08-22" gender="M" nation="POL" athleteid="3053">
              <RESULTS>
                <RESULT eventid="1090" points="184" swimtime="00:00:42.30" resultid="3054" heatid="4605" lane="6" entrytime="00:00:40.52" />
                <RESULT eventid="1320" points="132" swimtime="00:01:46.11" resultid="3055" heatid="4665" lane="2" entrytime="00:01:52.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="272" swimtime="00:01:41.97" resultid="3056" heatid="4690" lane="4" entrytime="00:01:58.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tyberiusz" lastname="Frymus" birthdate="1995-01-13" gender="M" nation="POL" athleteid="3045">
              <RESULTS>
                <RESULT eventid="1090" points="609" swimtime="00:00:26.30" resultid="3046" heatid="4616" lane="1" entrytime="00:00:25.59" />
                <RESULT eventid="1422" points="582" swimtime="00:01:12.33" resultid="3047" heatid="4693" lane="6" entrytime="00:01:08.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="609" swimtime="00:00:32.10" resultid="3048" heatid="4762" lane="2" entrytime="00:00:30.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Kowalczyk" birthdate="1976-01-31" gender="F" nation="POL" athleteid="3090">
              <RESULTS>
                <RESULT eventid="1059" points="471" swimtime="00:00:34.17" resultid="3091" heatid="4599" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1158" points="399" swimtime="00:12:28.65" resultid="3092" heatid="4631" lane="4" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                    <SPLIT distance="100" swimtime="00:01:28.55" />
                    <SPLIT distance="150" swimtime="00:02:16.59" />
                    <SPLIT distance="200" swimtime="00:03:04.81" />
                    <SPLIT distance="250" swimtime="00:03:53.28" />
                    <SPLIT distance="300" swimtime="00:04:41.46" />
                    <SPLIT distance="350" swimtime="00:05:29.09" />
                    <SPLIT distance="400" swimtime="00:06:17.08" />
                    <SPLIT distance="450" swimtime="00:07:04.94" />
                    <SPLIT distance="500" swimtime="00:07:52.04" />
                    <SPLIT distance="550" swimtime="00:08:39.15" />
                    <SPLIT distance="600" swimtime="00:09:26.13" />
                    <SPLIT distance="650" swimtime="00:10:13.28" />
                    <SPLIT distance="700" swimtime="00:11:00.23" />
                    <SPLIT distance="750" swimtime="00:11:46.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="445" swimtime="00:01:15.15" resultid="3093" heatid="4661" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="435" swimtime="00:02:51.67" resultid="3094" heatid="4716" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:23.63" />
                    <SPLIT distance="150" swimtime="00:02:08.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="430" swimtime="00:06:00.21" resultid="3095" heatid="4792" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:26.08" />
                    <SPLIT distance="150" swimtime="00:02:13.27" />
                    <SPLIT distance="200" swimtime="00:03:00.43" />
                    <SPLIT distance="250" swimtime="00:03:47.22" />
                    <SPLIT distance="300" swimtime="00:04:33.74" />
                    <SPLIT distance="350" swimtime="00:05:19.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Usewicz" birthdate="1994-08-12" gender="F" nation="POL" athleteid="3067">
              <RESULTS>
                <RESULT eventid="1059" points="416" swimtime="00:00:34.03" resultid="3068" heatid="4600" lane="1" entrytime="00:00:32.90" />
                <RESULT eventid="1303" points="416" swimtime="00:01:16.27" resultid="3069" heatid="4661" lane="8" entrytime="00:01:18.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="356" swimtime="00:02:55.63" resultid="3070" heatid="4715" lane="6" entrytime="00:02:56.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                    <SPLIT distance="100" swimtime="00:01:22.85" />
                    <SPLIT distance="150" swimtime="00:02:11.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="302" swimtime="00:06:25.19" resultid="3071" heatid="4793" lane="1" entrytime="00:06:40.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                    <SPLIT distance="100" swimtime="00:01:26.97" />
                    <SPLIT distance="150" swimtime="00:02:15.02" />
                    <SPLIT distance="200" swimtime="00:03:04.65" />
                    <SPLIT distance="250" swimtime="00:03:55.02" />
                    <SPLIT distance="300" swimtime="00:04:45.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grażyna" lastname="Kudra" birthdate="1959-11-24" gender="F" nation="POL" athleteid="3072">
              <RESULTS>
                <RESULT eventid="1059" points="170" swimtime="00:00:52.13" resultid="3119" heatid="4597" lane="6" entrytime="00:00:49.20" />
                <RESULT eventid="1404" points="315" swimtime="00:02:01.97" resultid="3120" heatid="4686" lane="2" entrytime="00:01:55.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="332" swimtime="00:00:54.02" resultid="3121" heatid="4753" lane="9" entrytime="00:00:49.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Moskalenko" birthdate="2000-12-01" gender="F" nation="POL" athleteid="3096">
              <RESULTS>
                <RESULT eventid="1059" swimtime="00:00:34.25" resultid="3097" heatid="4599" lane="7" entrytime="00:00:34.12" />
                <RESULT comment="Przekroczony limit czasu" eventid="1158" status="OTL" swimtime="00:13:08.03" resultid="3098" heatid="4631" lane="5" entrytime="00:13:05.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:28.34" />
                    <SPLIT distance="150" swimtime="00:02:16.00" />
                    <SPLIT distance="200" swimtime="00:03:04.10" />
                    <SPLIT distance="250" swimtime="00:03:53.41" />
                    <SPLIT distance="300" swimtime="00:04:42.83" />
                    <SPLIT distance="350" swimtime="00:05:33.34" />
                    <SPLIT distance="400" swimtime="00:06:24.59" />
                    <SPLIT distance="450" swimtime="00:07:15.90" />
                    <SPLIT distance="500" swimtime="00:08:06.80" />
                    <SPLIT distance="550" swimtime="00:08:58.57" />
                    <SPLIT distance="600" swimtime="00:09:49.76" />
                    <SPLIT distance="650" swimtime="00:10:40.74" />
                    <SPLIT distance="700" swimtime="00:11:31.79" />
                    <SPLIT distance="750" swimtime="00:12:22.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" swimtime="00:01:15.93" resultid="3099" heatid="4661" lane="5" entrytime="00:01:16.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" swimtime="00:02:55.24" resultid="3100" heatid="4715" lane="3" entrytime="00:02:55.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:24.47" />
                    <SPLIT distance="150" swimtime="00:02:11.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" swimtime="00:06:10.41" resultid="3101" heatid="4793" lane="2" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:25.93" />
                    <SPLIT distance="150" swimtime="00:02:12.84" />
                    <SPLIT distance="200" swimtime="00:03:00.00" />
                    <SPLIT distance="250" swimtime="00:03:47.63" />
                    <SPLIT distance="300" swimtime="00:04:36.08" />
                    <SPLIT distance="350" swimtime="00:05:25.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Rożek" birthdate="1984-05-09" gender="M" nation="POL" athleteid="3057">
              <RESULTS>
                <RESULT comment="Przekroczony limit czasu" eventid="1182" status="OTL" swimtime="00:13:38.40" resultid="3058" heatid="4634" lane="1" entrytime="00:13:37.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:31.51" />
                    <SPLIT distance="150" swimtime="00:02:21.63" />
                    <SPLIT distance="200" swimtime="00:03:12.92" />
                    <SPLIT distance="250" swimtime="00:04:05.19" />
                    <SPLIT distance="300" swimtime="00:04:57.52" />
                    <SPLIT distance="350" swimtime="00:05:49.51" />
                    <SPLIT distance="400" swimtime="00:06:42.57" />
                    <SPLIT distance="450" swimtime="00:07:35.36" />
                    <SPLIT distance="500" swimtime="00:08:28.74" />
                    <SPLIT distance="550" swimtime="00:09:21.64" />
                    <SPLIT distance="600" swimtime="00:10:13.97" />
                    <SPLIT distance="650" swimtime="00:11:05.81" />
                    <SPLIT distance="700" swimtime="00:11:58.89" />
                    <SPLIT distance="750" swimtime="00:12:50.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="322" swimtime="00:01:14.07" resultid="3059" heatid="4669" lane="6" entrytime="00:01:14.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="222" swimtime="00:00:39.85" resultid="3060" heatid="4700" lane="0" entrytime="00:00:37.71" />
                <RESULT eventid="1524" points="244" swimtime="00:03:00.40" resultid="3061" heatid="4721" lane="1" entrytime="00:02:55.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                    <SPLIT distance="100" swimtime="00:01:25.00" />
                    <SPLIT distance="150" swimtime="00:02:13.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="3062" heatid="4757" lane="5" entrytime="00:00:48.28" />
                <RESULT eventid="1766" points="238" reactiontime="+170" swimtime="00:06:36.29" resultid="3063" heatid="4800" lane="4" entrytime="00:06:31.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:26.33" />
                    <SPLIT distance="150" swimtime="00:02:14.62" />
                    <SPLIT distance="200" swimtime="00:03:05.36" />
                    <SPLIT distance="250" swimtime="00:03:58.17" />
                    <SPLIT distance="300" swimtime="00:04:51.76" />
                    <SPLIT distance="350" swimtime="00:05:45.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="535" swimtime="00:01:54.30" resultid="3115" heatid="4728" lane="8" entrytime="00:01:57.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.29" />
                    <SPLIT distance="100" swimtime="00:00:56.89" />
                    <SPLIT distance="150" swimtime="00:01:28.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3041" number="1" />
                    <RELAYPOSITION athleteid="3057" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="3049" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3045" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="431" swimtime="00:02:19.62" resultid="3118" heatid="4683" lane="4" entrytime="00:02:29.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:48.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3064" number="1" />
                    <RELAYPOSITION athleteid="3053" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="3049" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3057" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1371" points="386" swimtime="00:02:56.93" resultid="3113" heatid="4682" lane="1" entrytime="00:02:44.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.50" />
                    <SPLIT distance="100" swimtime="00:01:41.94" />
                    <SPLIT distance="150" swimtime="00:02:22.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3102" number="1" />
                    <RELAYPOSITION athleteid="3072" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="3076" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3067" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1541" points="337" swimtime="00:02:44.69" resultid="3114" heatid="4726" lane="1" entrytime="00:02:37.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:25.81" />
                    <SPLIT distance="150" swimtime="00:02:04.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3067" number="1" />
                    <RELAYPOSITION athleteid="3072" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="3076" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3102" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1718" points="419" swimtime="00:02:40.27" resultid="3116" heatid="4764" lane="5" entrytime="00:02:35.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                    <SPLIT distance="100" swimtime="00:01:33.75" />
                    <SPLIT distance="150" swimtime="00:02:08.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3102" number="1" />
                    <RELAYPOSITION athleteid="3076" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3049" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3057" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1141" points="541" swimtime="00:02:02.85" resultid="3117" heatid="4630" lane="1" entrytime="00:02:02.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                    <SPLIT distance="100" swimtime="00:01:00.43" />
                    <SPLIT distance="150" swimtime="00:01:37.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3045" number="1" />
                    <RELAYPOSITION athleteid="3067" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3076" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3041" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1718" points="407" swimtime="00:02:29.40" resultid="3111" heatid="4765" lane="0" entrytime="00:02:19.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                    <SPLIT distance="150" swimtime="00:01:55.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3045" number="1" />
                    <RELAYPOSITION athleteid="3072" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="3041" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3067" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1141" points="322" swimtime="00:02:33.10" resultid="3112" heatid="4629" lane="5" entrytime="00:02:33.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:23.44" />
                    <SPLIT distance="150" swimtime="00:02:01.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3057" number="1" />
                    <RELAYPOSITION athleteid="3072" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3102" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3049" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="7PBOT" nation="POL" clubid="4045" name="7 Pomorska Brygada Obrony Terytorialnej" shortname="7PBOT">
          <ATHLETES>
            <ATHLETE firstname="Rafał" lastname="Stasiukiewicz" birthdate="1980-01-01" gender="M" nation="POL" athleteid="2002">
              <RESULTS>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="2004" heatid="4655" lane="5" entrytime="00:04:30.00" />
                <RESULT eventid="1422" points="156" swimtime="00:01:58.05" resultid="2006" heatid="4690" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="195" swimtime="00:00:49.71" resultid="2008" heatid="4757" lane="7" entrytime="00:00:59.00" />
                <RESULT eventid="1766" points="136" swimtime="00:07:59.35" resultid="2009" heatid="4800" lane="2" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                    <SPLIT distance="100" swimtime="00:01:44.78" />
                    <SPLIT distance="150" swimtime="00:02:45.71" />
                    <SPLIT distance="200" swimtime="00:03:49.43" />
                    <SPLIT distance="250" swimtime="00:04:50.57" />
                    <SPLIT distance="300" swimtime="00:05:56.20" />
                    <SPLIT distance="350" swimtime="00:06:58.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="4013" heatid="4646" lane="1" entrytime="00:00:55.00" />
                <RESULT eventid="1490" points="110" swimtime="00:02:01.70" resultid="4026" heatid="4710" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MSB" nation="POL" region="06" clubid="2612" name="UKS JASIEŃ Sucha Beskidzka" shortname="JASIEŃ Sucha Beskidzka">
          <ATHLETES>
            <ATHLETE firstname="Aneta" lastname="Pytel" birthdate="1979-01-01" gender="F" nation="POL" athleteid="2619">
              <RESULTS>
                <RESULT eventid="1234" points="199" swimtime="00:00:50.67" resultid="2620" heatid="4641" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1269" points="244" swimtime="00:04:13.36" resultid="2621" heatid="4652" lane="4" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.12" />
                    <SPLIT distance="100" swimtime="00:02:02.37" />
                    <SPLIT distance="150" swimtime="00:03:08.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" status="DNS" swimtime="00:00:00.00" resultid="2622" heatid="4660" lane="1" entrytime="00:01:32.00" />
                <RESULT eventid="1473" points="195" swimtime="00:01:51.48" resultid="2623" heatid="4707" lane="8" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="100" swimtime="00:02:16.31" resultid="2624" heatid="4735" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="246" swimtime="00:00:51.71" resultid="4595" heatid="4753" lane="8" entrytime="00:00:48.06" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sabina" lastname="Sikora" birthdate="1984-01-01" gender="F" nation="POL" athleteid="2611">
              <RESULTS>
                <RESULT eventid="1269" points="433" swimtime="00:03:25.37" resultid="2613" heatid="4653" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:39.14" />
                    <SPLIT distance="150" swimtime="00:02:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="599" swimtime="00:01:08.89" resultid="2614" heatid="4661" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="530" swimtime="00:01:27.07" resultid="2615" heatid="4688" lane="0" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="565" swimtime="00:00:33.20" resultid="2616" heatid="4695" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1684" points="606" swimtime="00:00:37.03" resultid="2617" heatid="4755" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1742" points="429" swimtime="00:05:52.90" resultid="2618" heatid="4791" lane="0" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:01:23.21" />
                    <SPLIT distance="150" swimtime="00:02:08.41" />
                    <SPLIT distance="200" swimtime="00:02:53.69" />
                    <SPLIT distance="250" swimtime="00:03:39.96" />
                    <SPLIT distance="300" swimtime="00:04:25.73" />
                    <SPLIT distance="350" swimtime="00:05:11.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KSPIE" nation="POL" clubid="2153" name="Klub Sportowy Pietraszyn" shortname="KS Pietraszyn">
          <ATHLETES>
            <ATHLETE firstname="Adolf" lastname="Piechula" birthdate="1957-04-11" gender="M" nation="POL" athleteid="2154">
              <RESULTS>
                <RESULT eventid="1090" points="430" swimtime="00:00:34.70" resultid="2155" heatid="4607" lane="9" entrytime="00:00:36.34" entrycourse="SCM" />
                <RESULT eventid="1124" points="383" swimtime="00:03:19.95" resultid="2156" heatid="4625" lane="2" entrytime="00:03:10.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:01:37.32" />
                    <SPLIT distance="150" swimtime="00:02:34.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="406" swimtime="00:03:38.01" resultid="2157" heatid="4656" lane="5" entrytime="00:03:34.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                    <SPLIT distance="100" swimtime="00:01:42.91" />
                    <SPLIT distance="150" swimtime="00:02:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="325" swimtime="00:03:42.97" resultid="2158" heatid="4680" lane="1" entrytime="00:03:35.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                    <SPLIT distance="100" swimtime="00:01:45.19" />
                    <SPLIT distance="150" swimtime="00:02:44.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="448" swimtime="00:01:37.65" resultid="2159" heatid="4691" lane="1" entrytime="00:01:36.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="348" swimtime="00:07:25.37" resultid="2160" heatid="4788" lane="2" entrytime="00:07:24.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.09" />
                    <SPLIT distance="100" swimtime="00:01:48.72" />
                    <SPLIT distance="150" swimtime="00:02:45.57" />
                    <SPLIT distance="200" swimtime="00:03:42.55" />
                    <SPLIT distance="250" swimtime="00:04:44.62" />
                    <SPLIT distance="300" swimtime="00:05:44.43" />
                    <SPLIT distance="350" swimtime="00:06:35.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="263" swimtime="00:01:42.62" resultid="2161" heatid="4739" lane="0" entrytime="00:01:33.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="474" swimtime="00:00:42.68" resultid="2162" heatid="4758" lane="8" entrytime="00:00:44.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02805" nation="POL" region="05" clubid="2375" name="MUKS Zgierz">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Bednarek" birthdate="1951-03-24" gender="M" nation="POL" license="502805700052" athleteid="2455">
              <RESULTS>
                <RESULT eventid="1090" points="462" swimtime="00:00:35.82" resultid="2456" heatid="4607" lane="3" entrytime="00:00:34.50" entrycourse="LCM" />
                <RESULT eventid="1124" points="323" swimtime="00:03:57.39" resultid="2457" heatid="4624" lane="4" entrytime="00:03:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.17" />
                    <SPLIT distance="100" swimtime="00:01:55.27" />
                    <SPLIT distance="150" swimtime="00:03:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="458" swimtime="00:01:22.13" resultid="2458" heatid="4668" lane="0" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="403" swimtime="00:03:13.91" resultid="2459" heatid="4720" lane="8" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.87" />
                    <SPLIT distance="100" swimtime="00:01:32.49" />
                    <SPLIT distance="150" swimtime="00:02:24.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" status="DNS" swimtime="00:00:00.00" resultid="2460" heatid="4789" lane="3" entrytime="00:08:02.00" />
                <RESULT eventid="1766" points="364" swimtime="00:07:04.99" resultid="2461" heatid="4799" lane="0" entrytime="00:06:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.87" />
                    <SPLIT distance="100" swimtime="00:01:34.29" />
                    <SPLIT distance="150" swimtime="00:02:27.48" />
                    <SPLIT distance="200" swimtime="00:03:23.29" />
                    <SPLIT distance="250" swimtime="00:04:18.53" />
                    <SPLIT distance="300" swimtime="00:05:14.43" />
                    <SPLIT distance="350" swimtime="00:06:10.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Kajdos" birthdate="1976-06-25" gender="F" nation="POL" license="502805600148" athleteid="2497">
              <RESULTS>
                <RESULT eventid="1059" points="239" swimtime="00:00:42.79" resultid="2498" heatid="4598" lane="9" entrytime="00:00:42.87" entrycourse="LCM" />
                <RESULT eventid="1234" points="254" swimtime="00:00:48.95" resultid="2499" heatid="4641" lane="7" entrytime="00:00:48.44" entrycourse="LCM" />
                <RESULT eventid="1303" points="194" swimtime="00:01:39.12" resultid="2500" heatid="4659" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="238" swimtime="00:01:48.07" resultid="2501" heatid="4706" lane="5" entrytime="00:01:56.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="232" swimtime="00:03:54.34" resultid="2502" heatid="4744" lane="2" entrytime="00:03:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.88" />
                    <SPLIT distance="100" swimtime="00:01:54.23" />
                    <SPLIT distance="150" swimtime="00:02:56.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Łatecki" birthdate="1957-05-25" gender="M" nation="POL" license="502805700022" athleteid="2382">
              <RESULTS>
                <RESULT comment="Przekroczony limit czasu" eventid="1216" status="OTL" swimtime="00:35:49.47" resultid="2383" heatid="4638" lane="7" entrytime="00:29:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.67" />
                    <SPLIT distance="100" swimtime="00:02:08.59" />
                    <SPLIT distance="150" swimtime="00:03:18.57" />
                    <SPLIT distance="200" swimtime="00:04:30.05" />
                    <SPLIT distance="250" swimtime="00:05:41.00" />
                    <SPLIT distance="300" swimtime="00:06:52.58" />
                    <SPLIT distance="350" swimtime="00:08:03.07" />
                    <SPLIT distance="400" swimtime="00:09:14.50" />
                    <SPLIT distance="450" swimtime="00:10:25.76" />
                    <SPLIT distance="500" swimtime="00:11:37.79" />
                    <SPLIT distance="550" swimtime="00:12:50.45" />
                    <SPLIT distance="600" swimtime="00:14:02.98" />
                    <SPLIT distance="650" swimtime="00:15:13.69" />
                    <SPLIT distance="700" swimtime="00:16:25.78" />
                    <SPLIT distance="750" swimtime="00:17:36.82" />
                    <SPLIT distance="800" swimtime="00:18:49.00" />
                    <SPLIT distance="850" swimtime="00:20:01.56" />
                    <SPLIT distance="900" swimtime="00:21:14.48" />
                    <SPLIT distance="950" swimtime="00:22:26.14" />
                    <SPLIT distance="1000" swimtime="00:23:39.01" />
                    <SPLIT distance="1050" swimtime="00:24:51.59" />
                    <SPLIT distance="1100" swimtime="00:26:04.85" />
                    <SPLIT distance="1150" swimtime="00:27:18.44" />
                    <SPLIT distance="1200" swimtime="00:28:30.81" />
                    <SPLIT distance="1250" swimtime="00:29:42.92" />
                    <SPLIT distance="1300" swimtime="00:30:57.99" />
                    <SPLIT distance="1350" swimtime="00:32:12.61" />
                    <SPLIT distance="1400" swimtime="00:33:25.95" />
                    <SPLIT distance="1450" swimtime="00:34:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1354" status="DSQ" swimtime="00:00:00.00" resultid="2384" heatid="4679" lane="1" entrytime="00:05:00.00" entrycourse="LCM" />
                <RESULT eventid="1524" status="DNS" swimtime="00:00:00.00" resultid="2385" heatid="4719" lane="0" entrytime="00:04:00.00" entrycourse="LCM" />
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="2386" heatid="4801" lane="7" entrytime="00:08:00.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Kuśmider" birthdate="1989-03-07" gender="M" nation="POL" license="502805700" athleteid="2548">
              <RESULTS>
                <RESULT eventid="1090" points="397" swimtime="00:00:30.10" resultid="2549" heatid="4612" lane="5" entrytime="00:00:28.70" entrycourse="LCM" />
                <RESULT eventid="1216" points="431" swimtime="00:20:25.32" resultid="2550" heatid="4639" lane="3" entrytime="00:20:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:15.73" />
                    <SPLIT distance="150" swimtime="00:01:56.37" />
                    <SPLIT distance="200" swimtime="00:02:37.77" />
                    <SPLIT distance="250" swimtime="00:03:19.43" />
                    <SPLIT distance="300" swimtime="00:04:00.68" />
                    <SPLIT distance="350" swimtime="00:04:42.11" />
                    <SPLIT distance="400" swimtime="00:05:23.10" />
                    <SPLIT distance="450" swimtime="00:06:03.92" />
                    <SPLIT distance="500" swimtime="00:06:44.97" />
                    <SPLIT distance="550" swimtime="00:07:25.94" />
                    <SPLIT distance="600" swimtime="00:08:06.76" />
                    <SPLIT distance="650" swimtime="00:08:47.85" />
                    <SPLIT distance="700" swimtime="00:09:28.61" />
                    <SPLIT distance="750" swimtime="00:10:09.56" />
                    <SPLIT distance="800" swimtime="00:10:50.60" />
                    <SPLIT distance="850" swimtime="00:11:31.38" />
                    <SPLIT distance="900" swimtime="00:12:12.94" />
                    <SPLIT distance="950" swimtime="00:12:54.19" />
                    <SPLIT distance="1000" swimtime="00:13:35.19" />
                    <SPLIT distance="1050" swimtime="00:14:15.78" />
                    <SPLIT distance="1100" swimtime="00:14:57.00" />
                    <SPLIT distance="1150" swimtime="00:15:38.46" />
                    <SPLIT distance="1200" swimtime="00:16:19.86" />
                    <SPLIT distance="1250" swimtime="00:17:01.25" />
                    <SPLIT distance="1300" swimtime="00:17:42.65" />
                    <SPLIT distance="1350" swimtime="00:18:23.96" />
                    <SPLIT distance="1400" swimtime="00:19:05.53" />
                    <SPLIT distance="1450" swimtime="00:19:46.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" athleteid="2421">
              <RESULTS>
                <RESULT eventid="1059" points="666" swimtime="00:00:31.02" resultid="2422" heatid="4600" lane="2" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1107" points="677" swimtime="00:02:51.96" resultid="2423" heatid="4621" lane="1" entrytime="00:02:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                    <SPLIT distance="150" swimtime="00:02:11.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="575" swimtime="00:00:37.98" resultid="2424" heatid="4643" lane="1" entrytime="00:00:35.50" entrycourse="LCM" />
                <RESULT eventid="1439" points="693" swimtime="00:00:33.30" resultid="2425" heatid="4697" lane="9" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1473" points="556" swimtime="00:01:22.85" resultid="2426" heatid="4708" lane="6" entrytime="00:01:14.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="675" swimtime="00:01:17.26" resultid="2427" heatid="4736" lane="6" entrytime="00:01:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Wiczel" birthdate="1948-01-22" gender="M" nation="POL" license="502805700021" athleteid="2376">
              <RESULTS>
                <RESULT eventid="1286" points="672" swimtime="00:03:41.40" resultid="2377" heatid="4656" lane="6" entrytime="00:03:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.98" />
                    <SPLIT distance="100" swimtime="00:01:47.69" />
                    <SPLIT distance="150" swimtime="00:02:46.28" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1422" points="671" swimtime="00:01:40.22" resultid="2378" heatid="4691" lane="8" entrytime="00:01:39.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1490" points="448" swimtime="00:01:40.79" resultid="2379" heatid="4710" lane="5" entrytime="00:01:39.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.87" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1667" points="451" swimtime="00:03:41.99" resultid="2380" heatid="4747" lane="3" entrytime="00:03:38.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                    <SPLIT distance="100" swimtime="00:01:52.00" />
                    <SPLIT distance="150" swimtime="00:02:50.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="626" swimtime="00:00:44.55" resultid="2381" heatid="4758" lane="2" entrytime="00:00:43.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Morozowski" birthdate="1973-05-09" gender="M" nation="POL" license="102805700051" athleteid="2433">
              <RESULTS>
                <RESULT eventid="1216" points="311" swimtime="00:25:16.21" resultid="2434" heatid="4639" lane="8" entrytime="00:25:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:26.07" />
                    <SPLIT distance="150" swimtime="00:02:15.53" />
                    <SPLIT distance="200" swimtime="00:03:05.24" />
                    <SPLIT distance="250" swimtime="00:03:55.84" />
                    <SPLIT distance="300" swimtime="00:04:45.97" />
                    <SPLIT distance="350" swimtime="00:05:37.27" />
                    <SPLIT distance="400" swimtime="00:06:28.38" />
                    <SPLIT distance="450" swimtime="00:07:20.04" />
                    <SPLIT distance="500" swimtime="00:08:10.42" />
                    <SPLIT distance="550" swimtime="00:09:02.80" />
                    <SPLIT distance="600" swimtime="00:09:54.10" />
                    <SPLIT distance="650" swimtime="00:10:45.06" />
                    <SPLIT distance="700" swimtime="00:11:35.86" />
                    <SPLIT distance="750" swimtime="00:12:27.40" />
                    <SPLIT distance="800" swimtime="00:13:18.88" />
                    <SPLIT distance="850" swimtime="00:14:09.98" />
                    <SPLIT distance="900" swimtime="00:15:01.42" />
                    <SPLIT distance="950" swimtime="00:15:52.69" />
                    <SPLIT distance="1000" swimtime="00:16:43.93" />
                    <SPLIT distance="1050" swimtime="00:17:35.35" />
                    <SPLIT distance="1100" swimtime="00:18:25.47" />
                    <SPLIT distance="1150" swimtime="00:19:17.74" />
                    <SPLIT distance="1200" swimtime="00:20:08.74" />
                    <SPLIT distance="1250" swimtime="00:20:59.88" />
                    <SPLIT distance="1300" swimtime="00:21:51.53" />
                    <SPLIT distance="1350" swimtime="00:22:43.46" />
                    <SPLIT distance="1400" swimtime="00:23:35.51" />
                    <SPLIT distance="1450" swimtime="00:24:26.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="280" swimtime="00:03:40.72" resultid="2435" heatid="4657" lane="0" entrytime="00:03:26.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:42.19" />
                    <SPLIT distance="150" swimtime="00:02:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" status="DNS" swimtime="00:00:00.00" resultid="2436" heatid="4680" lane="7" entrytime="00:03:30.00" entrycourse="LCM" />
                <RESULT eventid="1422" points="321" swimtime="00:01:36.56" resultid="2437" heatid="4691" lane="7" entrytime="00:01:35.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="248" swimtime="00:07:34.33" resultid="2438" heatid="4789" lane="5" entrytime="00:08:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.27" />
                    <SPLIT distance="100" swimtime="00:01:50.14" />
                    <SPLIT distance="150" swimtime="00:02:51.71" />
                    <SPLIT distance="200" swimtime="00:03:55.61" />
                    <SPLIT distance="250" swimtime="00:04:55.19" />
                    <SPLIT distance="300" swimtime="00:05:55.75" />
                    <SPLIT distance="350" swimtime="00:06:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="355" swimtime="00:00:42.21" resultid="2439" heatid="4759" lane="9" entrytime="00:00:40.33" entrycourse="LCM" />
                <RESULT eventid="1766" points="304" swimtime="00:06:20.38" resultid="2440" heatid="4799" lane="1" entrytime="00:06:24.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:23.52" />
                    <SPLIT distance="150" swimtime="00:02:12.20" />
                    <SPLIT distance="200" swimtime="00:03:02.27" />
                    <SPLIT distance="250" swimtime="00:03:52.65" />
                    <SPLIT distance="300" swimtime="00:04:43.60" />
                    <SPLIT distance="350" swimtime="00:05:31.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-26" gender="F" nation="POL" license="502805600123" athleteid="2396">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="2397" heatid="4597" lane="5" entrytime="00:00:44.00" entrycourse="LCM" />
                <RESULT eventid="1107" points="142" swimtime="00:04:37.36" resultid="2398" heatid="4618" lane="4" entrytime="00:04:56.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.36" />
                    <SPLIT distance="100" swimtime="00:02:23.40" />
                    <SPLIT distance="150" swimtime="00:03:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="187" swimtime="00:04:36.72" resultid="2399" heatid="4652" lane="6" entrytime="00:04:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.05" />
                    <SPLIT distance="100" swimtime="00:02:14.60" />
                    <SPLIT distance="150" swimtime="00:03:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" status="DNS" swimtime="00:00:00.00" resultid="2400" heatid="4659" lane="3" entrytime="00:02:01.00" entrycourse="LCM" />
                <RESULT eventid="1404" points="189" swimtime="00:02:05.87" resultid="2401" heatid="4686" lane="0" entrytime="00:02:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="135" swimtime="00:00:55.26" resultid="2402" heatid="4694" lane="3" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1684" points="182" swimtime="00:00:57.16" resultid="2403" heatid="4752" lane="4" entrytime="00:00:50.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Przytulski" birthdate="1957-01-09" gender="M" nation="POL" license="502805700049" athleteid="2387">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="2388" heatid="4625" lane="3" entrytime="00:03:05.00" entrycourse="LCM" />
                <RESULT eventid="1182" points="483" swimtime="00:12:47.09" resultid="2389" heatid="4634" lane="4" entrytime="00:12:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                    <SPLIT distance="150" swimtime="00:02:13.70" />
                    <SPLIT distance="200" swimtime="00:03:01.80" />
                    <SPLIT distance="250" swimtime="00:03:50.79" />
                    <SPLIT distance="300" swimtime="00:04:39.88" />
                    <SPLIT distance="350" swimtime="00:05:29.34" />
                    <SPLIT distance="400" swimtime="00:06:18.63" />
                    <SPLIT distance="450" swimtime="00:07:08.18" />
                    <SPLIT distance="500" swimtime="00:07:57.62" />
                    <SPLIT distance="550" swimtime="00:08:46.79" />
                    <SPLIT distance="600" swimtime="00:09:36.81" />
                    <SPLIT distance="650" swimtime="00:10:25.90" />
                    <SPLIT distance="700" swimtime="00:11:14.48" />
                    <SPLIT distance="750" swimtime="00:12:02.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="2390" heatid="4648" lane="2" entrytime="00:00:39.00" entrycourse="LCM" />
                <RESULT eventid="1354" points="400" swimtime="00:03:28.07" resultid="2391" heatid="4680" lane="2" entrytime="00:03:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                    <SPLIT distance="100" swimtime="00:01:37.45" />
                    <SPLIT distance="150" swimtime="00:02:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" status="DNS" swimtime="00:00:00.00" resultid="2392" heatid="4701" lane="9" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1597" points="408" swimtime="00:07:02.47" resultid="2393" heatid="4788" lane="6" entrytime="00:07:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                    <SPLIT distance="100" swimtime="00:01:38.58" />
                    <SPLIT distance="150" swimtime="00:02:33.63" />
                    <SPLIT distance="200" swimtime="00:03:29.10" />
                    <SPLIT distance="250" swimtime="00:04:33.38" />
                    <SPLIT distance="300" swimtime="00:05:36.74" />
                    <SPLIT distance="350" swimtime="00:06:20.26" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1633" points="469" swimtime="00:01:24.71" resultid="2394" heatid="4739" lane="7" entrytime="00:01:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="2395" heatid="4799" lane="3" entrytime="00:06:05.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Rembowska-Świeboda" birthdate="1968-06-27" gender="F" nation="POL" license="102805600031" athleteid="2428">
              <RESULTS>
                <RESULT eventid="1059" points="588" swimtime="00:00:33.72" resultid="2429" heatid="4599" lane="5" entrytime="00:00:33.74" entrycourse="LCM" />
                <RESULT eventid="1234" points="561" swimtime="00:00:38.77" resultid="2430" heatid="4642" lane="2" entrytime="00:00:38.80" entrycourse="LCM" />
                <RESULT eventid="1303" points="530" swimtime="00:01:16.62" resultid="2431" heatid="4661" lane="0" entrytime="00:01:18.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="555" swimtime="00:01:24.79" resultid="2432" heatid="4708" lane="9" entrytime="00:01:25.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Ścibiorek" birthdate="1997-02-19" gender="M" nation="POL" license="502805700" athleteid="2534">
              <RESULTS>
                <RESULT eventid="1490" points="519" swimtime="00:01:08.52" resultid="2535" heatid="4713" lane="1" entrytime="00:01:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="526" swimtime="00:02:32.05" resultid="2536" heatid="4750" lane="2" entrytime="00:02:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:01:53.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Rudziński" birthdate="1966-05-10" gender="M" nation="POL" license="502805700162" athleteid="2503">
              <RESULTS>
                <RESULT eventid="1286" points="345" swimtime="00:03:34.59" resultid="2504" heatid="4656" lane="3" entrytime="00:03:35.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:41.43" />
                    <SPLIT distance="150" swimtime="00:02:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="213" swimtime="00:03:48.81" resultid="2505" heatid="4680" lane="9" entrytime="00:03:47.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.86" />
                    <SPLIT distance="100" swimtime="00:01:45.49" />
                    <SPLIT distance="150" swimtime="00:02:47.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="254" swimtime="00:00:41.90" resultid="2506" heatid="4699" lane="8" entrytime="00:00:40.98" entrycourse="LCM" />
                <RESULT eventid="1597" points="227" swimtime="00:08:07.21" resultid="2507" heatid="4788" lane="8" entrytime="00:07:51.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                    <SPLIT distance="100" swimtime="00:01:48.82" />
                    <SPLIT distance="150" swimtime="00:03:03.37" />
                    <SPLIT distance="200" swimtime="00:04:19.83" />
                    <SPLIT distance="250" swimtime="00:05:21.71" />
                    <SPLIT distance="300" swimtime="00:06:23.30" />
                    <SPLIT distance="350" swimtime="00:07:17.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="229" swimtime="00:01:38.94" resultid="2508" heatid="4738" lane="4" entrytime="00:01:40.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="327" swimtime="00:00:43.53" resultid="2509" heatid="4756" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Klusek" birthdate="1975-01-12" gender="F" nation="POL" license="502805600030" athleteid="2528">
              <RESULTS>
                <RESULT eventid="1107" points="416" swimtime="00:03:09.37" resultid="2529" heatid="4620" lane="7" entrytime="00:03:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:27.78" />
                    <SPLIT distance="150" swimtime="00:02:23.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1337" points="364" swimtime="00:03:22.11" resultid="2530" heatid="4677" lane="1" entrytime="00:03:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:32.47" />
                    <SPLIT distance="150" swimtime="00:02:25.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="460" swimtime="00:01:33.70" resultid="2531" heatid="4687" lane="2" entrytime="00:01:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="462" swimtime="00:06:45.80" resultid="2532" heatid="4785" lane="1" entrytime="00:06:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:31.75" />
                    <SPLIT distance="150" swimtime="00:02:27.49" />
                    <SPLIT distance="200" swimtime="00:03:22.49" />
                    <SPLIT distance="250" swimtime="00:04:17.51" />
                    <SPLIT distance="300" swimtime="00:05:13.89" />
                    <SPLIT distance="350" swimtime="00:05:58.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="385" swimtime="00:06:13.68" resultid="2533" heatid="4792" lane="8" entrytime="00:05:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:25.03" />
                    <SPLIT distance="150" swimtime="00:02:12.29" />
                    <SPLIT distance="200" swimtime="00:03:01.05" />
                    <SPLIT distance="250" swimtime="00:03:50.57" />
                    <SPLIT distance="300" swimtime="00:04:39.32" />
                    <SPLIT distance="350" swimtime="00:05:27.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Dziarek" birthdate="1959-02-19" gender="M" nation="POL" license="502805700029" athleteid="2450">
              <RESULTS>
                <RESULT eventid="1216" points="391" swimtime="00:24:31.08" resultid="2451" heatid="4639" lane="0" entrytime="00:26:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:26.81" />
                    <SPLIT distance="150" swimtime="00:02:14.50" />
                    <SPLIT distance="200" swimtime="00:03:02.62" />
                    <SPLIT distance="250" swimtime="00:03:51.90" />
                    <SPLIT distance="300" swimtime="00:04:41.02" />
                    <SPLIT distance="350" swimtime="00:05:30.59" />
                    <SPLIT distance="400" swimtime="00:06:19.42" />
                    <SPLIT distance="450" swimtime="00:07:08.93" />
                    <SPLIT distance="500" swimtime="00:07:57.93" />
                    <SPLIT distance="550" swimtime="00:08:47.23" />
                    <SPLIT distance="600" swimtime="00:09:36.28" />
                    <SPLIT distance="650" swimtime="00:10:25.80" />
                    <SPLIT distance="700" swimtime="00:11:14.00" />
                    <SPLIT distance="750" swimtime="00:12:03.48" />
                    <SPLIT distance="800" swimtime="00:12:52.38" />
                    <SPLIT distance="850" swimtime="00:13:42.35" />
                    <SPLIT distance="900" swimtime="00:14:31.40" />
                    <SPLIT distance="950" swimtime="00:15:21.83" />
                    <SPLIT distance="1000" swimtime="00:16:10.84" />
                    <SPLIT distance="1050" swimtime="00:17:01.28" />
                    <SPLIT distance="1100" swimtime="00:17:50.69" />
                    <SPLIT distance="1150" swimtime="00:18:41.13" />
                    <SPLIT distance="1200" swimtime="00:19:29.73" />
                    <SPLIT distance="1250" swimtime="00:20:20.07" />
                    <SPLIT distance="1300" swimtime="00:21:09.95" />
                    <SPLIT distance="1350" swimtime="00:22:01.04" />
                    <SPLIT distance="1400" swimtime="00:22:51.46" />
                    <SPLIT distance="1450" swimtime="00:23:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="468" swimtime="00:01:14.24" resultid="2452" heatid="4667" lane="2" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="413" swimtime="00:02:51.40" resultid="2453" heatid="4720" lane="3" entrytime="00:03:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:19.01" />
                    <SPLIT distance="150" swimtime="00:02:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="413" swimtime="00:06:08.87" resultid="2454" heatid="4799" lane="9" entrytime="00:06:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:01:24.38" />
                    <SPLIT distance="150" swimtime="00:02:11.68" />
                    <SPLIT distance="200" swimtime="00:02:59.77" />
                    <SPLIT distance="250" swimtime="00:03:47.09" />
                    <SPLIT distance="300" swimtime="00:04:35.55" />
                    <SPLIT distance="350" swimtime="00:05:22.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="502805600152" athleteid="2479">
              <RESULTS>
                <RESULT eventid="1107" points="258" swimtime="00:03:41.94" resultid="2480" heatid="4619" lane="1" entrytime="00:03:49.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.45" />
                    <SPLIT distance="100" swimtime="00:01:54.19" />
                    <SPLIT distance="150" swimtime="00:02:55.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="267" swimtime="00:27:10.00" resultid="2481" heatid="4637" lane="3" entrytime="00:27:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                    <SPLIT distance="100" swimtime="00:01:40.51" />
                    <SPLIT distance="150" swimtime="00:02:34.59" />
                    <SPLIT distance="200" swimtime="00:03:28.63" />
                    <SPLIT distance="250" swimtime="00:04:23.34" />
                    <SPLIT distance="300" swimtime="00:05:17.81" />
                    <SPLIT distance="350" swimtime="00:06:12.31" />
                    <SPLIT distance="400" swimtime="00:07:06.12" />
                    <SPLIT distance="450" swimtime="00:08:00.77" />
                    <SPLIT distance="500" swimtime="00:08:55.47" />
                    <SPLIT distance="550" swimtime="00:09:50.09" />
                    <SPLIT distance="600" swimtime="00:10:44.87" />
                    <SPLIT distance="650" swimtime="00:11:41.15" />
                    <SPLIT distance="700" swimtime="00:12:35.18" />
                    <SPLIT distance="750" swimtime="00:13:30.23" />
                    <SPLIT distance="800" swimtime="00:14:24.12" />
                    <SPLIT distance="850" swimtime="00:15:19.94" />
                    <SPLIT distance="900" swimtime="00:16:14.63" />
                    <SPLIT distance="950" swimtime="00:17:10.70" />
                    <SPLIT distance="1000" swimtime="00:18:05.62" />
                    <SPLIT distance="1050" swimtime="00:19:01.67" />
                    <SPLIT distance="1100" swimtime="00:19:56.03" />
                    <SPLIT distance="1150" swimtime="00:20:50.93" />
                    <SPLIT distance="1200" swimtime="00:21:44.81" />
                    <SPLIT distance="1250" swimtime="00:22:40.24" />
                    <SPLIT distance="1300" swimtime="00:23:35.25" />
                    <SPLIT distance="1350" swimtime="00:24:30.57" />
                    <SPLIT distance="1400" swimtime="00:25:25.63" />
                    <SPLIT distance="1450" swimtime="00:26:19.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="315" swimtime="00:04:00.51" resultid="2482" heatid="4653" lane="0" entrytime="00:03:58.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.20" />
                    <SPLIT distance="100" swimtime="00:01:56.57" />
                    <SPLIT distance="150" swimtime="00:02:59.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1337" points="215" swimtime="00:04:00.92" resultid="2483" heatid="4676" lane="5" entrytime="00:03:57.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.18" />
                    <SPLIT distance="100" swimtime="00:01:56.31" />
                    <SPLIT distance="150" swimtime="00:02:59.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="275" swimtime="00:03:19.97" resultid="2484" heatid="4715" lane="7" entrytime="00:03:19.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                    <SPLIT distance="100" swimtime="00:01:38.36" />
                    <SPLIT distance="150" swimtime="00:02:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="261" swimtime="00:08:10.54" resultid="2485" heatid="4785" lane="9" entrytime="00:08:12.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.68" />
                    <SPLIT distance="100" swimtime="00:02:01.11" />
                    <SPLIT distance="150" swimtime="00:03:07.93" />
                    <SPLIT distance="200" swimtime="00:04:15.46" />
                    <SPLIT distance="250" swimtime="00:05:19.53" />
                    <SPLIT distance="300" swimtime="00:06:23.80" />
                    <SPLIT distance="350" swimtime="00:07:18.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="177" swimtime="00:04:16.18" resultid="2486" heatid="4743" lane="4" entrytime="00:04:21.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.62" />
                    <SPLIT distance="100" swimtime="00:02:10.77" />
                    <SPLIT distance="150" swimtime="00:03:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="264" swimtime="00:07:03.85" resultid="2487" heatid="4793" lane="8" entrytime="00:06:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.18" />
                    <SPLIT distance="100" swimtime="00:01:40.80" />
                    <SPLIT distance="150" swimtime="00:02:36.69" />
                    <SPLIT distance="200" swimtime="00:03:30.82" />
                    <SPLIT distance="250" swimtime="00:04:25.41" />
                    <SPLIT distance="300" swimtime="00:05:20.19" />
                    <SPLIT distance="350" swimtime="00:06:13.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-01-05" gender="F" nation="POL" license="502805600055" athleteid="2462">
              <RESULTS>
                <RESULT eventid="1059" points="300" swimtime="00:00:39.72" resultid="2463" heatid="4598" lane="7" entrytime="00:00:39.02" entrycourse="LCM" />
                <RESULT eventid="1107" points="258" swimtime="00:03:41.97" resultid="2464" heatid="4619" lane="2" entrytime="00:03:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.52" />
                    <SPLIT distance="100" swimtime="00:01:54.89" />
                    <SPLIT distance="150" swimtime="00:02:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="281" swimtime="00:00:47.33" resultid="2465" heatid="4640" lane="2" />
                <RESULT eventid="1269" points="373" swimtime="00:03:47.45" resultid="2466" heatid="4653" lane="6" entrytime="00:03:40.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.63" />
                    <SPLIT distance="100" swimtime="00:01:51.16" />
                    <SPLIT distance="150" swimtime="00:02:49.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="343" swimtime="00:01:43.27" resultid="2467" heatid="4687" lane="8" entrytime="00:01:43.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="240" swimtime="00:01:47.83" resultid="2468" heatid="4707" lane="0" entrytime="00:01:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="256" swimtime="00:03:46.64" resultid="2469" heatid="4744" lane="7" entrytime="00:03:50.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.55" />
                    <SPLIT distance="100" swimtime="00:01:54.73" />
                    <SPLIT distance="150" swimtime="00:02:54.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="346" swimtime="00:00:47.79" resultid="2470" heatid="4753" lane="4" entrytime="00:00:46.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Dziedziczak" birthdate="1977-02-04" gender="M" nation="POL" license="502805700153" athleteid="2471">
              <RESULTS>
                <RESULT eventid="1090" points="425" swimtime="00:00:31.31" resultid="2472" heatid="4609" lane="7" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1124" points="312" swimtime="00:03:11.62" resultid="2473" heatid="4625" lane="4" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:27.87" />
                    <SPLIT distance="150" swimtime="00:02:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="277" swimtime="00:00:42.36" resultid="2474" heatid="4648" lane="8" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1320" points="385" swimtime="00:01:11.78" resultid="2475" heatid="4670" lane="6" entrytime="00:01:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="407" swimtime="00:00:34.05" resultid="2476" heatid="4700" lane="3" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1524" points="323" swimtime="00:02:51.47" resultid="2477" heatid="4722" lane="0" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                    <SPLIT distance="100" swimtime="00:01:20.92" />
                    <SPLIT distance="150" swimtime="00:02:07.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="293" swimtime="00:03:17.99" resultid="2478" heatid="4748" lane="6" entrytime="00:03:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                    <SPLIT distance="100" swimtime="00:01:36.70" />
                    <SPLIT distance="150" swimtime="00:02:29.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dagmara" lastname="Luźniakowska" birthdate="1980-04-29" gender="F" nation="POL" license="502805600154" athleteid="2405">
              <RESULTS>
                <RESULT eventid="1059" points="304" swimtime="00:00:39.32" resultid="2406" heatid="4599" lane="0" entrytime="00:00:36.52" entrycourse="LCM" />
                <RESULT eventid="1303" points="331" swimtime="00:01:23.88" resultid="2407" heatid="4661" lane="9" entrytime="00:01:18.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="280" swimtime="00:00:43.33" resultid="2408" heatid="4695" lane="9" entrytime="00:00:42.87" entrycourse="LCM" />
                <RESULT eventid="1507" points="376" swimtime="00:02:59.07" resultid="2409" heatid="4715" lane="5" entrytime="00:02:53.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:28.26" />
                    <SPLIT distance="150" swimtime="00:02:14.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" status="DNS" swimtime="00:00:00.00" resultid="2410" heatid="4751" lane="3" />
                <RESULT eventid="1742" points="334" swimtime="00:06:18.56" resultid="2411" heatid="4793" lane="7" entrytime="00:06:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:01:29.93" />
                    <SPLIT distance="150" swimtime="00:02:18.60" />
                    <SPLIT distance="200" swimtime="00:03:07.32" />
                    <SPLIT distance="250" swimtime="00:03:56.74" />
                    <SPLIT distance="300" swimtime="00:04:45.03" />
                    <SPLIT distance="350" swimtime="00:05:34.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Sypniewski" birthdate="1957-02-01" gender="M" nation="POL" license="102805700035" athleteid="2488">
              <RESULTS>
                <RESULT eventid="1090" points="457" swimtime="00:00:34.02" resultid="2489" heatid="4608" lane="2" entrytime="00:00:33.45" entrycourse="LCM" />
                <RESULT eventid="1124" points="306" swimtime="00:03:35.41" resultid="2490" heatid="4625" lane="1" entrytime="00:03:26.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                    <SPLIT distance="100" swimtime="00:01:43.81" />
                    <SPLIT distance="150" swimtime="00:02:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="409" swimtime="00:00:41.69" resultid="2491" heatid="4647" lane="4" entrytime="00:00:40.93" entrycourse="LCM" />
                <RESULT eventid="1286" points="345" swimtime="00:03:50.18" resultid="2492" heatid="4656" lane="7" entrytime="00:03:43.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.56" />
                    <SPLIT distance="100" swimtime="00:01:49.44" />
                    <SPLIT distance="150" swimtime="00:02:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" status="DNS" swimtime="00:00:00.00" resultid="2493" heatid="4699" lane="3" entrytime="00:00:38.08" entrycourse="LCM" />
                <RESULT eventid="1490" points="409" swimtime="00:01:31.80" resultid="2494" heatid="4711" lane="9" entrytime="00:01:36.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" status="DNS" swimtime="00:00:00.00" resultid="2495" heatid="4738" lane="2" entrytime="00:01:48.95" entrycourse="LCM" />
                <RESULT eventid="1701" points="458" swimtime="00:00:43.17" resultid="2496" heatid="4758" lane="1" entrytime="00:00:44.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sergiusz" lastname="Olejniczak" birthdate="1978-12-01" gender="M" nation="POL" license="502805700058" athleteid="2537">
              <RESULTS>
                <RESULT eventid="1252" points="497" swimtime="00:00:34.86" resultid="2538" heatid="4651" lane="0" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1286" points="458" swimtime="00:03:00.88" resultid="2539" heatid="4658" lane="7" entrytime="00:02:38.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:25.68" />
                    <SPLIT distance="150" swimtime="00:02:12.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="468" swimtime="00:01:23.42" resultid="2540" heatid="4693" lane="7" entrytime="00:01:11.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="455" swimtime="00:01:18.16" resultid="2541" heatid="4713" lane="0" entrytime="00:01:09.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="507" swimtime="00:02:44.91" resultid="2542" heatid="4750" lane="7" entrytime="00:02:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                    <SPLIT distance="100" swimtime="00:01:19.10" />
                    <SPLIT distance="150" swimtime="00:02:02.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="487" swimtime="00:00:37.12" resultid="2543" heatid="4761" lane="2" entrytime="00:00:34.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" athleteid="2412">
              <RESULTS>
                <RESULT eventid="1059" points="576" swimtime="00:00:34.72" resultid="2413" heatid="4599" lane="1" entrytime="00:00:34.76" entrycourse="LCM" />
                <RESULT eventid="1107" points="551" swimtime="00:03:20.70" resultid="2414" heatid="4619" lane="5" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.32" />
                    <SPLIT distance="100" swimtime="00:01:38.08" />
                    <SPLIT distance="150" swimtime="00:02:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="534" swimtime="00:00:41.68" resultid="2415" heatid="4641" lane="5" entrytime="00:00:42.55" entrycourse="LCM" />
                <RESULT eventid="1303" points="529" swimtime="00:01:18.89" resultid="2416" heatid="4661" lane="7" entrytime="00:01:17.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1439" points="664" swimtime="00:00:35.65" resultid="2417" heatid="4695" lane="5" entrytime="00:00:36.34" entrycourse="LCM" />
                <RESULT eventid="1473" points="470" swimtime="00:01:35.50" resultid="2418" heatid="4707" lane="7" entrytime="00:01:37.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="487" swimtime="00:01:31.53" resultid="2419" heatid="4736" lane="0" entrytime="00:01:30.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="576" swimtime="00:00:44.98" resultid="2420" heatid="4754" lane="9" entrytime="00:00:45.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Jasiński" birthdate="1960-07-23" gender="M" nation="POL" license="502805700027" athleteid="2441">
              <RESULTS>
                <RESULT eventid="1090" points="410" swimtime="00:00:33.95" resultid="2442" heatid="4608" lane="8" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT comment="Z2 - Pływak pokonał jednym stylem więcej niż 1 dystansu." eventid="1124" status="DSQ" swimtime="00:03:41.53" resultid="2443" heatid="4625" lane="9" entrytime="00:03:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:50.39" />
                    <SPLIT distance="150" swimtime="00:02:53.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="365" swimtime="00:03:43.12" resultid="2444" heatid="4656" lane="2" entrytime="00:03:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.86" />
                    <SPLIT distance="100" swimtime="00:01:47.23" />
                    <SPLIT distance="150" swimtime="00:02:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2445" heatid="4669" lane="1" entrytime="00:01:15.00" entrycourse="LCM" />
                <RESULT eventid="1422" points="354" swimtime="00:01:41.18" resultid="2446" heatid="4691" lane="5" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="340" swimtime="00:00:39.58" resultid="2447" heatid="4699" lane="5" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1701" points="386" swimtime="00:00:43.86" resultid="2448" heatid="4758" lane="3" entrytime="00:00:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Wypych-Staszewska" birthdate="1970-08-16" gender="F" nation="POL" license="502805600164" athleteid="2510">
              <RESULTS>
                <RESULT eventid="1107" points="392" swimtime="00:03:26.27" resultid="2511" heatid="4619" lane="3" entrytime="00:03:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:01:37.05" />
                    <SPLIT distance="150" swimtime="00:02:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="328" swimtime="00:13:52.27" resultid="2512" heatid="4631" lane="6" entrytime="00:13:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                    <SPLIT distance="100" swimtime="00:01:37.68" />
                    <SPLIT distance="150" swimtime="00:02:26.29" />
                    <SPLIT distance="200" swimtime="00:03:24.63" />
                    <SPLIT distance="250" swimtime="00:04:17.03" />
                    <SPLIT distance="300" swimtime="00:05:10.07" />
                    <SPLIT distance="350" swimtime="00:06:02.32" />
                    <SPLIT distance="400" swimtime="00:06:54.85" />
                    <SPLIT distance="450" swimtime="00:07:47.30" />
                    <SPLIT distance="500" swimtime="00:08:40.39" />
                    <SPLIT distance="550" swimtime="00:09:33.34" />
                    <SPLIT distance="600" swimtime="00:10:26.53" />
                    <SPLIT distance="650" swimtime="00:11:19.57" />
                    <SPLIT distance="700" swimtime="00:12:12.47" />
                    <SPLIT distance="750" swimtime="00:13:04.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="373" swimtime="00:00:43.88" resultid="2513" heatid="4640" lane="1" />
                <RESULT eventid="1337" points="348" swimtime="00:03:35.33" resultid="2514" heatid="4676" lane="4" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.04" />
                    <SPLIT distance="100" swimtime="00:01:46.31" />
                    <SPLIT distance="150" swimtime="00:02:43.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="406" swimtime="00:00:39.77" resultid="2515" heatid="4695" lane="7" entrytime="00:00:39.00" entrycourse="LCM" />
                <RESULT eventid="1573" points="385" swimtime="00:07:20.77" resultid="2516" heatid="4786" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.88" />
                    <SPLIT distance="100" swimtime="00:01:46.77" />
                    <SPLIT distance="150" swimtime="00:02:43.05" />
                    <SPLIT distance="200" swimtime="00:03:41.02" />
                    <SPLIT distance="250" swimtime="00:04:42.75" />
                    <SPLIT distance="300" swimtime="00:05:45.79" />
                    <SPLIT distance="350" swimtime="00:06:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="325" swimtime="00:01:38.60" resultid="2517" heatid="4736" lane="9" entrytime="00:01:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="338" swimtime="00:03:30.49" resultid="2518" heatid="4744" lane="3" entrytime="00:03:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.34" />
                    <SPLIT distance="100" swimtime="00:01:43.92" />
                    <SPLIT distance="150" swimtime="00:02:40.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Lis-Piwowarski" birthdate="1984-05-29" gender="M" nation="POL" license="502805700146" athleteid="2519">
              <RESULTS>
                <RESULT eventid="1090" points="223" swimtime="00:00:37.51" resultid="2520" heatid="4606" lane="2" entrytime="00:00:37.34" entrycourse="LCM" />
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu." eventid="1124" status="DSQ" swimtime="00:04:44.44" resultid="2521" heatid="4623" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.47" />
                    <SPLIT distance="100" swimtime="00:02:10.12" />
                    <SPLIT distance="150" swimtime="00:03:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="101" swimtime="00:00:56.07" resultid="2522" heatid="4645" lane="8" />
                <RESULT eventid="1320" points="152" swimtime="00:01:35.01" resultid="2523" heatid="4666" lane="2" entrytime="00:01:33.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="111" swimtime="00:00:50.21" resultid="2524" heatid="4698" lane="7" entrytime="00:00:48.20" entrycourse="LCM" />
                <RESULT eventid="1524" points="120" swimtime="00:03:48.70" resultid="2525" heatid="4719" lane="8" entrytime="00:03:57.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.51" />
                    <SPLIT distance="100" swimtime="00:01:43.85" />
                    <SPLIT distance="150" swimtime="00:02:47.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="94" swimtime="00:01:57.72" resultid="2526" heatid="4737" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="117" swimtime="00:00:57.89" resultid="2527" heatid="4756" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kotulski" birthdate="1981-07-03" gender="M" nation="POL" license="502805700" athleteid="2544">
              <RESULTS>
                <RESULT eventid="1090" points="406" swimtime="00:00:31.33" resultid="2545" heatid="4608" lane="6" entrytime="00:00:33.04" entrycourse="LCM" />
                <RESULT eventid="1320" points="332" swimtime="00:01:13.90" resultid="2546" heatid="4668" lane="4" entrytime="00:01:15.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="366" swimtime="00:00:33.97" resultid="2547" heatid="4701" lane="1" entrytime="00:00:33.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="456" swimtime="00:02:32.54" resultid="2558" heatid="4683" lane="5" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:24.82" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2387" number="1" />
                    <RELAYPOSITION athleteid="2488" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="2537" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="2450" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="445" swimtime="00:02:14.09" resultid="2559" heatid="4727" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:10.27" />
                    <SPLIT distance="150" swimtime="00:01:44.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2455" number="1" />
                    <RELAYPOSITION athleteid="2488" number="2" reactiontime="+21" />
                    <RELAYPOSITION athleteid="2450" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2537" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1395" points="358" swimtime="00:02:35.96" resultid="2560" heatid="4683" lane="3" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.84" />
                    <SPLIT distance="100" swimtime="00:01:30.38" />
                    <SPLIT distance="150" swimtime="00:02:06.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2441" number="1" />
                    <RELAYPOSITION athleteid="2433" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="2471" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="2544" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1565" points="436" swimtime="00:02:09.47" resultid="2564" heatid="4727" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:07.88" />
                    <SPLIT distance="150" swimtime="00:01:38.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2441" number="1" />
                    <RELAYPOSITION athleteid="2433" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="2544" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2471" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1541" points="640" swimtime="00:02:13.08" resultid="2551" heatid="4726" lane="2" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:08.63" />
                    <SPLIT distance="150" swimtime="00:01:41.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2412" number="1" />
                    <RELAYPOSITION athleteid="2528" number="2" reactiontime="+17" />
                    <RELAYPOSITION athleteid="2428" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="2421" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1371" points="632" swimtime="00:02:30.11" resultid="2552" heatid="4682" lane="2" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:21.43" />
                    <SPLIT distance="150" swimtime="00:01:55.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2428" number="1" />
                    <RELAYPOSITION athleteid="2528" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="2421" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2412" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1371" points="377" swimtime="00:02:52.63" resultid="2556" heatid="4682" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.88" />
                    <SPLIT distance="100" swimtime="00:01:34.66" />
                    <SPLIT distance="150" swimtime="00:02:14.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2497" number="1" />
                    <RELAYPOSITION athleteid="2462" number="2" reactiontime="-4" />
                    <RELAYPOSITION athleteid="2510" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="2405" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1541" points="337" swimtime="00:02:35.68" resultid="2557" heatid="4726" lane="7" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="150" swimtime="00:01:54.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2462" number="1" />
                    <RELAYPOSITION athleteid="2405" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2510" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="2479" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1141" points="495" swimtime="00:02:12.67" resultid="2553" heatid="4630" lane="9" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:07.66" />
                    <SPLIT distance="150" swimtime="00:01:40.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2428" number="1" />
                    <RELAYPOSITION athleteid="2441" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2528" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2471" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1718" points="605" swimtime="00:02:31.39" resultid="2561" heatid="4764" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:22.00" />
                    <SPLIT distance="150" swimtime="00:01:58.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2387" number="1" />
                    <RELAYPOSITION athleteid="2421" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2412" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2450" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1141" points="297" swimtime="00:02:33.18" resultid="2555" heatid="4630" lane="0" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2497" number="1" />
                    <RELAYPOSITION athleteid="2433" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2510" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2519" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1718" points="416" swimtime="00:02:40.73" resultid="2562" heatid="4764" lane="2" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:29.49" />
                    <SPLIT distance="150" swimtime="00:02:03.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2488" number="1" />
                    <RELAYPOSITION athleteid="2462" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="2471" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2405" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1718" points="453" swimtime="00:02:36.18" resultid="2554" heatid="4764" lane="6" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                    <SPLIT distance="100" swimtime="00:01:31.03" />
                    <SPLIT distance="150" swimtime="00:02:03.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2497" number="1" />
                    <RELAYPOSITION athleteid="2528" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2537" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2441" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1718" points="365" swimtime="00:02:38.37" resultid="2563" heatid="4764" lane="7" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:53.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2534" number="1" />
                    <RELAYPOSITION athleteid="2433" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2510" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2396" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="10414" nation="POL" region="14" clubid="2953" name="KS MAKO Warszawa" shortname="MAKO Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Rurak" birthdate="1988-05-09" gender="M" nation="POL" athleteid="2954">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="2955" heatid="4616" lane="0" entrytime="00:00:25.66" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Safrończyk" birthdate="1988-05-30" gender="M" nation="POL" athleteid="2973">
              <RESULTS>
                <RESULT eventid="1090" points="737" swimtime="00:00:25.19" resultid="2974" heatid="4616" lane="8" entrytime="00:00:25.66" />
                <RESULT eventid="1422" points="734" swimtime="00:01:09.16" resultid="2975" heatid="4693" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1701" points="826" swimtime="00:00:30.21" resultid="2976" heatid="4762" lane="5" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Butkiewicz" birthdate="1980-03-19" gender="F" nation="POL" athleteid="2956">
              <RESULTS>
                <RESULT eventid="1059" points="510" swimtime="00:00:33.08" resultid="2957" heatid="4600" lane="0" entrytime="00:00:33.00" />
                <RESULT comment="Przekroczony limit czasu" eventid="1158" status="OTL" swimtime="00:13:53.90" resultid="2958" heatid="4631" lane="3" entrytime="00:13:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:01:31.32" />
                    <SPLIT distance="150" swimtime="00:02:22.38" />
                    <SPLIT distance="200" swimtime="00:03:15.37" />
                    <SPLIT distance="250" swimtime="00:04:09.30" />
                    <SPLIT distance="300" swimtime="00:05:03.31" />
                    <SPLIT distance="350" swimtime="00:05:56.76" />
                    <SPLIT distance="400" swimtime="00:06:51.20" />
                    <SPLIT distance="450" swimtime="00:07:45.64" />
                    <SPLIT distance="500" swimtime="00:08:39.93" />
                    <SPLIT distance="550" swimtime="00:09:34.80" />
                    <SPLIT distance="600" swimtime="00:10:28.77" />
                    <SPLIT distance="650" swimtime="00:11:23.08" />
                    <SPLIT distance="700" swimtime="00:12:16.38" />
                    <SPLIT distance="750" swimtime="00:13:07.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" status="DNS" swimtime="00:00:00.00" resultid="2959" heatid="4660" lane="8" entrytime="00:01:35.00" />
                <RESULT eventid="1439" points="438" swimtime="00:00:37.32" resultid="2960" heatid="4695" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1507" points="394" swimtime="00:02:56.29" resultid="2961" heatid="4715" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:23.27" />
                    <SPLIT distance="150" swimtime="00:02:11.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Suda" birthdate="1978-02-20" gender="M" nation="POL" athleteid="2987">
              <RESULTS>
                <RESULT eventid="1320" points="332" swimtime="00:01:15.44" resultid="2988" heatid="4667" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kosiela" birthdate="1985-02-03" gender="M" nation="POL" athleteid="2980">
              <RESULTS>
                <RESULT eventid="1090" points="244" swimtime="00:00:36.38" resultid="2981" heatid="4606" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1124" points="204" swimtime="00:03:33.27" resultid="2982" heatid="4624" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                    <SPLIT distance="100" swimtime="00:01:42.32" />
                    <SPLIT distance="150" swimtime="00:02:44.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="227" swimtime="00:00:39.56" resultid="2983" heatid="4699" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Wiatr" birthdate="1984-05-21" gender="F" nation="POL" athleteid="2977">
              <RESULTS>
                <RESULT eventid="1059" points="306" swimtime="00:00:38.55" resultid="2978" heatid="4598" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1303" points="265" swimtime="00:01:30.40" resultid="2979" heatid="4660" lane="6" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Solecka" birthdate="1974-07-13" gender="F" nation="POL" athleteid="2962">
              <RESULTS>
                <RESULT eventid="1059" points="338" swimtime="00:00:38.17" resultid="2963" heatid="4598" lane="3" entrytime="00:00:38.23" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Siergiej" lastname="Kulinicz" birthdate="1984-01-01" gender="M" nation="POL" athleteid="2989" />
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" athleteid="2967">
              <RESULTS>
                <RESULT eventid="1090" points="266" swimtime="00:00:37.98" resultid="2968" heatid="4606" lane="0" entrytime="00:00:38.38" />
                <RESULT eventid="1252" points="252" swimtime="00:00:45.96" resultid="2969" heatid="4646" lane="6" entrytime="00:00:50.28" />
                <RESULT eventid="1320" points="287" swimtime="00:01:24.80" resultid="2970" heatid="4666" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="230" swimtime="00:03:22.13" resultid="2971" heatid="4719" lane="2" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:36.93" />
                    <SPLIT distance="150" swimtime="00:02:30.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="212" swimtime="00:03:55.92" resultid="2972" heatid="4747" lane="7" entrytime="00:03:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.96" />
                    <SPLIT distance="100" swimtime="00:01:56.51" />
                    <SPLIT distance="150" swimtime="00:02:58.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Pacławska" birthdate="1981-11-03" gender="F" nation="POL" athleteid="2984">
              <RESULTS>
                <RESULT eventid="1234" points="153" swimtime="00:00:55.37" resultid="2985" heatid="4641" lane="8" entrytime="00:00:52.00" />
                <RESULT eventid="1473" points="131" swimtime="00:02:07.17" resultid="2986" heatid="4706" lane="4" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Bystry" birthdate="1977-03-14" gender="M" nation="POL" athleteid="2964">
              <RESULTS>
                <RESULT eventid="1090" points="521" swimtime="00:00:29.25" resultid="2965" heatid="4613" lane="9" entrytime="00:00:28.50" />
                <RESULT eventid="1456" status="DNS" swimtime="00:00:00.00" resultid="2966" heatid="4702" lane="9" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="403" swimtime="00:02:22.75" resultid="2993" heatid="4683" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                    <SPLIT distance="100" swimtime="00:01:15.62" />
                    <SPLIT distance="150" swimtime="00:01:54.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2967" number="1" />
                    <RELAYPOSITION athleteid="2973" number="2" reactiontime="-20" />
                    <RELAYPOSITION athleteid="2980" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="2989" number="4" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="1565" status="DSQ" swimtime="00:02:00.24" resultid="2994" heatid="4728" lane="0" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.17" />
                    <SPLIT distance="100" swimtime="00:00:59.25" />
                    <SPLIT distance="150" swimtime="00:01:31.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2973" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2980" number="2" reactiontime="+62" status="DSQ" />
                    <RELAYPOSITION athleteid="2987" number="3" reactiontime="+54" status="DSQ" />
                    <RELAYPOSITION athleteid="2989" number="4" reactiontime="+42" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="1141" status="DSQ" swimtime="00:02:01.62" resultid="2990" heatid="4630" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.13" />
                    <SPLIT distance="100" swimtime="00:00:53.25" />
                    <SPLIT distance="150" swimtime="00:01:25.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2973" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2964" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="2956" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="2977" number="4" reactiontime="+22" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZ" nation="POL" clubid="1925" name="Niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Tobiasz" lastname="Jankowski" birthdate="1983-01-01" gender="M" nation="POL" athleteid="3642">
              <RESULTS>
                <RESULT eventid="1456" points="396" swimtime="00:00:33.10" resultid="3643" heatid="4701" lane="8" entrytime="00:00:33.70" />
                <RESULT eventid="1701" points="511" swimtime="00:00:36.07" resultid="3644" heatid="4760" lane="3" entrytime="00:00:36.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Karnaszewski" birthdate="1994-01-01" gender="M" nation="POL" athleteid="2625">
              <RESULTS>
                <RESULT eventid="1090" points="690" swimtime="00:00:25.23" resultid="2626" heatid="4617" lane="6" entrytime="00:00:24.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Grzybowski" birthdate="2000-01-01" gender="M" nation="POL" athleteid="2656">
              <RESULTS>
                <RESULT eventid="1090" swimtime="00:00:25.35" resultid="2657" heatid="4617" lane="7" entrytime="00:00:24.33" />
                <RESULT eventid="1124" swimtime="00:02:28.27" resultid="2658" heatid="4627" lane="7" entrytime="00:02:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                    <SPLIT distance="150" swimtime="00:01:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" swimtime="00:00:28.01" resultid="2659" heatid="4651" lane="5" entrytime="00:00:27.20" />
                <RESULT eventid="1320" swimtime="00:00:56.49" resultid="2660" heatid="4675" lane="2" entrytime="00:00:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" swimtime="00:00:26.34" resultid="2661" heatid="4705" lane="2" entrytime="00:00:25.90" />
                <RESULT eventid="1490" swimtime="00:01:03.15" resultid="2662" heatid="4713" lane="2" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M1 - Pływak nie złamał powierzchni wody głową przed lub na linii 15 m po starcie lub nawrocie." eventid="1633" status="DSQ" swimtime="00:00:59.75" resultid="2663" heatid="4741" lane="2" entrytime="00:01:05.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" swimtime="00:00:35.83" resultid="2664" heatid="4760" lane="4" entrytime="00:00:35.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Bryła" birthdate="1992-01-01" gender="M" nation="POL" athleteid="3600">
              <RESULTS>
                <RESULT eventid="1090" points="233" swimtime="00:00:35.93" resultid="3601" heatid="4610" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1124" points="180" swimtime="00:03:36.37" resultid="3602" heatid="4626" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                    <SPLIT distance="100" swimtime="00:01:46.24" />
                    <SPLIT distance="150" swimtime="00:02:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="313" swimtime="00:03:23.17" resultid="3603" heatid="4657" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                    <SPLIT distance="100" swimtime="00:01:34.02" />
                    <SPLIT distance="150" swimtime="00:02:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="189" swimtime="00:01:26.63" resultid="3604" heatid="4670" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="325" swimtime="00:01:29.01" resultid="3605" heatid="4692" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="196" swimtime="00:03:08.35" resultid="3606" heatid="4722" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:24.93" />
                    <SPLIT distance="150" swimtime="00:02:16.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="319" swimtime="00:00:40.58" resultid="3607" heatid="4759" lane="5" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tadeusz" lastname="Vorbrodt" birthdate="1953-01-01" gender="M" nation="POL" athleteid="4803">
              <RESULTS>
                <RESULT eventid="1252" points="223" swimtime="00:00:55.34" resultid="4805" heatid="4644" lane="6" late="yes" />
                <RESULT eventid="1490" points="207" swimtime="00:02:04.15" resultid="4806" heatid="4709" lane="9" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" status="DNS" swimtime="00:00:00.00" resultid="4807" heatid="4746" lane="8" late="yes" />
                <RESULT eventid="1766" points="272" swimtime="00:07:48.38" resultid="5399" heatid="4801" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.56" />
                    <SPLIT distance="100" swimtime="00:01:51.35" />
                    <SPLIT distance="150" swimtime="00:02:49.57" />
                    <SPLIT distance="200" swimtime="00:03:48.59" />
                    <SPLIT distance="250" swimtime="00:04:48.95" />
                    <SPLIT distance="300" swimtime="00:05:50.33" />
                    <SPLIT distance="350" swimtime="00:06:51.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Teodorczyk" birthdate="1985-01-01" gender="M" nation="POL" athleteid="1932">
              <RESULTS>
                <RESULT eventid="1124" points="486" swimtime="00:02:39.76" resultid="1933" heatid="4626" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:02:02.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="585" swimtime="00:01:00.70" resultid="1934" heatid="4672" lane="3" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="527" swimtime="00:00:29.87" resultid="1935" heatid="4702" lane="5" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Gruca" birthdate="2000-01-01" gender="F" nation="POL" athleteid="3634">
              <RESULTS>
                <RESULT eventid="1107" swimtime="00:03:00.95" resultid="3635" heatid="4618" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:24.30" />
                    <SPLIT distance="150" swimtime="00:02:15.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" swimtime="00:03:20.20" resultid="3636" heatid="4654" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                    <SPLIT distance="100" swimtime="00:01:34.44" />
                    <SPLIT distance="150" swimtime="00:02:28.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" swimtime="00:01:35.16" resultid="3637" heatid="4688" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" swimtime="00:00:36.46" resultid="3638" heatid="4695" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1684" status="DNS" swimtime="00:00:00.00" resultid="3639" heatid="4754" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1303" swimtime="00:01:15.19" resultid="3640" heatid="4660" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1059" swimtime="00:00:31.93" resultid="3641" heatid="4598" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Bistron" birthdate="1989-01-01" gender="M" nation="POL" athleteid="4040">
              <RESULTS>
                <RESULT eventid="1354" points="171" swimtime="00:03:42.16" resultid="4041" heatid="4679" lane="5" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.74" />
                    <SPLIT distance="100" swimtime="00:01:43.80" />
                    <SPLIT distance="150" swimtime="00:02:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="174" swimtime="00:01:40.12" resultid="4042" heatid="4710" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" status="DNS" swimtime="00:00:00.00" resultid="4043" heatid="4746" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Szymański" birthdate="1978-01-01" gender="M" nation="POL" athleteid="2010">
              <RESULTS>
                <RESULT eventid="1090" points="493" swimtime="00:00:29.80" resultid="2011" heatid="4610" lane="3" entrytime="00:00:30.60" />
                <RESULT eventid="1252" points="468" swimtime="00:00:35.57" resultid="2012" heatid="4648" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1320" points="472" swimtime="00:01:07.09" resultid="2013" heatid="4671" lane="0" entrytime="00:01:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="430" swimtime="00:01:19.63" resultid="2014" heatid="4711" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernard" lastname="Poloczek" birthdate="1947-02-25" gender="M" nation="POL" athleteid="2015">
              <RESULTS>
                <RESULT eventid="1090" points="400" swimtime="00:00:39.59" resultid="2016" heatid="4605" lane="4" entrytime="00:00:39.30" />
                <RESULT eventid="1252" points="405" swimtime="00:00:46.53" resultid="2017" heatid="4647" lane="9" entrytime="00:00:45.70" />
                <RESULT eventid="1320" points="313" swimtime="00:01:37.72" resultid="2018" heatid="4666" lane="0" entrytime="00:01:36.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="324" swimtime="00:00:46.20" resultid="2019" heatid="4698" lane="3" entrytime="00:00:45.70" />
                <RESULT eventid="1490" points="392" swimtime="00:01:45.36" resultid="2020" heatid="4710" lane="6" entrytime="00:01:43.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="343" swimtime="00:04:02.99" resultid="2021" heatid="4747" lane="2" entrytime="00:03:53.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.20" />
                    <SPLIT distance="100" swimtime="00:01:56.61" />
                    <SPLIT distance="150" swimtime="00:03:00.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Źródlak" birthdate="1997-01-01" gender="M" nation="POL" athleteid="2637">
              <RESULTS>
                <RESULT eventid="1090" points="421" swimtime="00:00:29.74" resultid="2638" heatid="4611" lane="9" entrytime="00:00:30.02" />
                <RESULT eventid="1252" points="326" swimtime="00:00:36.95" resultid="2639" heatid="4648" lane="4" entrytime="00:00:36.80" />
                <RESULT eventid="1320" points="389" swimtime="00:01:09.07" resultid="2640" heatid="4667" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="297" swimtime="00:01:22.54" resultid="2641" heatid="4711" lane="6" entrytime="00:01:29.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="307" swimtime="00:00:40.33" resultid="2642" heatid="4758" lane="5" entrytime="00:00:41.71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anton" lastname="Bortnik" birthdate="1987-01-01" gender="M" nation="POL" athleteid="2670">
              <RESULTS>
                <RESULT eventid="1090" points="432" swimtime="00:00:30.09" resultid="2671" heatid="4609" lane="6" entrytime="00:00:31.89" />
                <RESULT eventid="1320" points="406" swimtime="00:01:08.56" resultid="2672" heatid="4670" lane="8" entrytime="00:01:11.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Pomierny" birthdate="1978-01-01" gender="M" nation="POL" athleteid="2668">
              <RESULTS>
                <RESULT eventid="1182" points="440" swimtime="00:11:24.32" resultid="2669" heatid="4635" lane="2" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="100" swimtime="00:01:21.81" />
                    <SPLIT distance="150" swimtime="00:02:04.83" />
                    <SPLIT distance="200" swimtime="00:02:48.25" />
                    <SPLIT distance="250" swimtime="00:03:31.80" />
                    <SPLIT distance="300" swimtime="00:04:15.02" />
                    <SPLIT distance="350" swimtime="00:04:58.13" />
                    <SPLIT distance="400" swimtime="00:05:41.48" />
                    <SPLIT distance="450" swimtime="00:06:24.83" />
                    <SPLIT distance="500" swimtime="00:07:08.17" />
                    <SPLIT distance="550" swimtime="00:07:51.38" />
                    <SPLIT distance="600" swimtime="00:08:34.88" />
                    <SPLIT distance="650" swimtime="00:09:18.29" />
                    <SPLIT distance="700" swimtime="00:10:01.62" />
                    <SPLIT distance="750" swimtime="00:10:44.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Wiśniewski" birthdate="2002-01-01" gender="M" nation="POL" athleteid="2680">
              <RESULTS>
                <RESULT eventid="1090" swimtime="00:00:26.17" resultid="2681" heatid="4616" lane="3" entrytime="00:00:25.01" />
                <RESULT eventid="1252" swimtime="00:00:33.35" resultid="2682" heatid="4651" lane="9" entrytime="00:00:30.12" />
                <RESULT eventid="1320" swimtime="00:00:59.55" resultid="2683" heatid="4675" lane="0" entrytime="00:00:56.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" swimtime="00:00:29.16" resultid="2684" heatid="4703" lane="6" entrytime="00:00:29.32" />
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="2685" heatid="4761" lane="3" entrytime="00:00:33.34" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Szydłowski" birthdate="1998-01-01" gender="M" nation="POL" athleteid="1953">
              <RESULTS>
                <RESULT eventid="1320" points="338" swimtime="00:01:12.42" resultid="1954" heatid="4666" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Lubiński" birthdate="1992-01-01" gender="M" nation="POL" athleteid="1993">
              <RESULTS>
                <RESULT eventid="1124" points="430" swimtime="00:02:41.84" resultid="1994" heatid="4626" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:17.24" />
                    <SPLIT distance="150" swimtime="00:02:03.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="361" swimtime="00:11:25.78" resultid="1995" heatid="4635" lane="7" entrytime="00:11:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:01.83" />
                    <SPLIT distance="200" swimtime="00:02:44.21" />
                    <SPLIT distance="250" swimtime="00:03:26.42" />
                    <SPLIT distance="300" swimtime="00:04:09.43" />
                    <SPLIT distance="350" swimtime="00:04:52.50" />
                    <SPLIT distance="400" swimtime="00:05:35.74" />
                    <SPLIT distance="450" swimtime="00:06:19.33" />
                    <SPLIT distance="500" swimtime="00:07:03.72" />
                    <SPLIT distance="550" swimtime="00:07:47.53" />
                    <SPLIT distance="600" swimtime="00:08:31.75" />
                    <SPLIT distance="650" swimtime="00:09:16.22" />
                    <SPLIT distance="700" swimtime="00:10:00.73" />
                    <SPLIT distance="750" swimtime="00:10:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="1996" heatid="4649" lane="7" entrytime="00:00:34.83" />
                <RESULT eventid="1354" points="244" swimtime="00:03:17.38" resultid="1997" heatid="4680" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="100" swimtime="00:01:35.37" />
                    <SPLIT distance="150" swimtime="00:02:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="403" swimtime="00:00:31.47" resultid="1998" heatid="4701" lane="7" entrytime="00:00:33.50" />
                <RESULT eventid="1597" points="349" swimtime="00:06:10.34" resultid="1999" heatid="4787" lane="0" entrytime="00:05:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:28.14" />
                    <SPLIT distance="150" swimtime="00:02:16.73" />
                    <SPLIT distance="200" swimtime="00:03:04.73" />
                    <SPLIT distance="250" swimtime="00:03:54.98" />
                    <SPLIT distance="300" swimtime="00:04:46.66" />
                    <SPLIT distance="350" swimtime="00:05:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="339" swimtime="00:02:56.04" resultid="2000" heatid="4749" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                    <SPLIT distance="100" swimtime="00:01:26.15" />
                    <SPLIT distance="150" swimtime="00:02:11.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="397" swimtime="00:05:23.91" resultid="2001" heatid="4797" lane="2" entrytime="00:05:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:16.67" />
                    <SPLIT distance="150" swimtime="00:01:57.07" />
                    <SPLIT distance="200" swimtime="00:02:37.48" />
                    <SPLIT distance="250" swimtime="00:03:18.59" />
                    <SPLIT distance="300" swimtime="00:04:00.17" />
                    <SPLIT distance="350" swimtime="00:04:42.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Grochowski" birthdate="1991-01-01" gender="M" nation="POL" athleteid="1939">
              <RESULTS>
                <RESULT eventid="1182" points="382" swimtime="00:11:12.98" resultid="1940" heatid="4635" lane="3" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:19.05" />
                    <SPLIT distance="150" swimtime="00:02:00.59" />
                    <SPLIT distance="200" swimtime="00:02:42.96" />
                    <SPLIT distance="250" swimtime="00:03:25.19" />
                    <SPLIT distance="300" swimtime="00:04:07.51" />
                    <SPLIT distance="350" swimtime="00:04:50.09" />
                    <SPLIT distance="400" swimtime="00:05:32.80" />
                    <SPLIT distance="450" swimtime="00:06:15.50" />
                    <SPLIT distance="500" swimtime="00:06:57.60" />
                    <SPLIT distance="550" swimtime="00:07:39.93" />
                    <SPLIT distance="600" swimtime="00:08:22.24" />
                    <SPLIT distance="650" swimtime="00:09:05.02" />
                    <SPLIT distance="700" swimtime="00:09:47.85" />
                    <SPLIT distance="750" swimtime="00:10:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="320" swimtime="00:00:37.96" resultid="1941" heatid="4648" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1422" points="368" swimtime="00:01:25.44" resultid="1942" heatid="4689" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="409" swimtime="00:05:20.68" resultid="1943" heatid="4797" lane="0" entrytime="00:05:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                    <SPLIT distance="100" swimtime="00:01:18.53" />
                    <SPLIT distance="150" swimtime="00:01:59.63" />
                    <SPLIT distance="200" swimtime="00:02:40.78" />
                    <SPLIT distance="250" swimtime="00:03:21.70" />
                    <SPLIT distance="300" swimtime="00:04:02.32" />
                    <SPLIT distance="350" swimtime="00:04:42.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Gleb" birthdate="1967-01-01" gender="M" nation="POL" athleteid="1936">
              <RESULTS>
                <RESULT eventid="1090" points="426" swimtime="00:00:32.49" resultid="1937" heatid="4610" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1216" points="428" swimtime="00:23:03.24" resultid="1938" heatid="4639" lane="1" entrytime="00:22:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:01:23.17" />
                    <SPLIT distance="150" swimtime="00:02:09.07" />
                    <SPLIT distance="200" swimtime="00:02:55.34" />
                    <SPLIT distance="250" swimtime="00:03:42.35" />
                    <SPLIT distance="300" swimtime="00:04:29.41" />
                    <SPLIT distance="350" swimtime="00:05:15.24" />
                    <SPLIT distance="400" swimtime="00:06:01.03" />
                    <SPLIT distance="450" swimtime="00:06:47.33" />
                    <SPLIT distance="500" swimtime="00:07:33.87" />
                    <SPLIT distance="550" swimtime="00:08:20.24" />
                    <SPLIT distance="600" swimtime="00:09:07.26" />
                    <SPLIT distance="650" swimtime="00:09:54.76" />
                    <SPLIT distance="700" swimtime="00:10:42.38" />
                    <SPLIT distance="750" swimtime="00:11:29.82" />
                    <SPLIT distance="800" swimtime="00:12:17.25" />
                    <SPLIT distance="850" swimtime="00:13:04.52" />
                    <SPLIT distance="900" swimtime="00:13:52.12" />
                    <SPLIT distance="950" swimtime="00:14:38.82" />
                    <SPLIT distance="1000" swimtime="00:15:25.15" />
                    <SPLIT distance="1050" swimtime="00:16:11.44" />
                    <SPLIT distance="1100" swimtime="00:16:57.52" />
                    <SPLIT distance="1150" swimtime="00:17:43.01" />
                    <SPLIT distance="1200" swimtime="00:18:29.56" />
                    <SPLIT distance="1250" swimtime="00:19:15.80" />
                    <SPLIT distance="1300" swimtime="00:20:02.62" />
                    <SPLIT distance="1350" swimtime="00:20:49.04" />
                    <SPLIT distance="1400" swimtime="00:21:35.21" />
                    <SPLIT distance="1450" swimtime="00:22:20.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Opałko" birthdate="1999-01-01" gender="F" nation="POL" athleteid="2643">
              <RESULTS>
                <RESULT eventid="1059" swimtime="00:00:30.97" resultid="2644" heatid="4601" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1107" swimtime="00:02:55.03" resultid="2645" heatid="4620" lane="5" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                    <SPLIT distance="150" swimtime="00:02:11.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" swimtime="00:00:37.18" resultid="2646" heatid="4643" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1303" swimtime="00:01:09.70" resultid="2647" heatid="4662" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" swimtime="00:00:34.41" resultid="2648" heatid="4696" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1473" swimtime="00:01:23.18" resultid="2649" heatid="4708" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" swimtime="00:01:27.34" resultid="2650" heatid="4736" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" swimtime="00:00:40.53" resultid="2651" heatid="4754" lane="5" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ciecior" birthdate="1953-11-24" gender="M" nation="POL" athleteid="2022">
              <RESULTS>
                <RESULT comment="K13 - Pływak nie zwrócił stóp na zewnątrz w trakcie napędzającej części ruchu nóg." eventid="1124" status="DSQ" swimtime="00:03:47.63" resultid="2023" heatid="4624" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.00" />
                    <SPLIT distance="100" swimtime="00:01:50.17" />
                    <SPLIT distance="150" swimtime="00:02:58.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="376" swimtime="00:28:18.69" resultid="2024" heatid="4638" lane="5" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:42.28" />
                    <SPLIT distance="150" swimtime="00:02:38.29" />
                    <SPLIT distance="200" swimtime="00:03:35.15" />
                    <SPLIT distance="250" swimtime="00:04:31.67" />
                    <SPLIT distance="300" swimtime="00:05:28.06" />
                    <SPLIT distance="350" swimtime="00:06:24.87" />
                    <SPLIT distance="400" swimtime="00:07:21.71" />
                    <SPLIT distance="450" swimtime="00:08:18.21" />
                    <SPLIT distance="500" swimtime="00:09:15.54" />
                    <SPLIT distance="550" swimtime="00:10:11.64" />
                    <SPLIT distance="600" swimtime="00:11:08.80" />
                    <SPLIT distance="650" swimtime="00:12:05.07" />
                    <SPLIT distance="700" swimtime="00:13:02.61" />
                    <SPLIT distance="750" swimtime="00:13:58.78" />
                    <SPLIT distance="800" swimtime="00:14:56.48" />
                    <SPLIT distance="850" swimtime="00:15:52.91" />
                    <SPLIT distance="900" swimtime="00:16:50.40" />
                    <SPLIT distance="950" swimtime="00:17:47.77" />
                    <SPLIT distance="1000" swimtime="00:18:46.40" />
                    <SPLIT distance="1050" swimtime="00:19:43.93" />
                    <SPLIT distance="1100" swimtime="00:20:41.32" />
                    <SPLIT distance="1150" swimtime="00:21:38.01" />
                    <SPLIT distance="1200" swimtime="00:22:35.68" />
                    <SPLIT distance="1250" swimtime="00:23:33.63" />
                    <SPLIT distance="1300" swimtime="00:24:31.78" />
                    <SPLIT distance="1350" swimtime="00:25:29.06" />
                    <SPLIT distance="1400" swimtime="00:26:27.37" />
                    <SPLIT distance="1450" swimtime="00:27:24.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="459" swimtime="00:00:43.53" resultid="2025" heatid="4647" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1354" points="247" swimtime="00:04:26.31" resultid="2026" heatid="4679" lane="2" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.71" />
                    <SPLIT distance="100" swimtime="00:02:04.25" />
                    <SPLIT distance="150" swimtime="00:03:16.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="359" swimtime="00:01:43.34" resultid="2027" heatid="4710" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="344" swimtime="00:08:27.86" resultid="2028" heatid="4788" lane="0" entrytime="00:07:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.03" />
                    <SPLIT distance="100" swimtime="00:02:05.64" />
                    <SPLIT distance="150" swimtime="00:03:10.48" />
                    <SPLIT distance="200" swimtime="00:04:15.85" />
                    <SPLIT distance="250" swimtime="00:05:28.29" />
                    <SPLIT distance="300" swimtime="00:06:40.79" />
                    <SPLIT distance="350" swimtime="00:07:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="211" swimtime="00:01:53.16" resultid="2029" heatid="4738" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="332" swimtime="00:03:51.20" resultid="2030" heatid="4748" lane="9" entrytime="00:03:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.75" />
                    <SPLIT distance="100" swimtime="00:01:54.08" />
                    <SPLIT distance="150" swimtime="00:02:54.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Konieczny" birthdate="1998-01-01" gender="M" nation="POL" athleteid="3645">
              <RESULTS>
                <RESULT eventid="1124" points="228" swimtime="00:03:22.16" resultid="3646" heatid="4624" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:35.56" />
                    <SPLIT distance="150" swimtime="00:02:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="281" swimtime="00:01:16.94" resultid="3647" heatid="4667" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="233" swimtime="00:00:38.53" resultid="3648" heatid="4700" lane="1" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Łopuszyński" birthdate="1969-01-01" gender="M" nation="POL" athleteid="1926">
              <RESULTS>
                <RESULT eventid="1124" points="152" swimtime="00:04:05.67" resultid="1927" heatid="4623" lane="4" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                    <SPLIT distance="100" swimtime="00:01:59.51" />
                    <SPLIT distance="150" swimtime="00:03:09.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="136" swimtime="00:04:18.72" resultid="1928" heatid="4679" lane="6" entrytime="00:04:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.12" />
                    <SPLIT distance="100" swimtime="00:01:59.44" />
                    <SPLIT distance="150" swimtime="00:03:07.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="131" swimtime="00:00:50.86" resultid="1929" heatid="4698" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1597" points="145" swimtime="00:09:03.03" resultid="1930" heatid="4789" lane="7" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.98" />
                    <SPLIT distance="100" swimtime="00:02:00.32" />
                    <SPLIT distance="150" swimtime="00:03:18.75" />
                    <SPLIT distance="200" swimtime="00:04:32.38" />
                    <SPLIT distance="250" swimtime="00:05:44.87" />
                    <SPLIT distance="300" swimtime="00:06:59.15" />
                    <SPLIT distance="350" swimtime="00:08:01.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="124" swimtime="00:01:54.61" resultid="1931" heatid="4738" lane="7" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Kamiński" birthdate="1965-01-01" gender="M" nation="POL" athleteid="1965">
              <RESULTS>
                <RESULT eventid="1090" points="355" swimtime="00:00:34.50" resultid="1966" heatid="4606" lane="4" entrytime="00:00:36.82" />
                <RESULT eventid="1182" points="344" swimtime="00:12:50.53" resultid="1967" heatid="4633" lane="4" entrytime="00:14:19.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:12.60" />
                    <SPLIT distance="200" swimtime="00:02:59.67" />
                    <SPLIT distance="250" swimtime="00:03:47.91" />
                    <SPLIT distance="300" swimtime="00:04:36.26" />
                    <SPLIT distance="350" swimtime="00:05:25.33" />
                    <SPLIT distance="400" swimtime="00:06:14.37" />
                    <SPLIT distance="450" swimtime="00:07:03.06" />
                    <SPLIT distance="500" swimtime="00:07:51.77" />
                    <SPLIT distance="550" swimtime="00:08:41.59" />
                    <SPLIT distance="600" swimtime="00:09:30.61" />
                    <SPLIT distance="650" swimtime="00:10:19.96" />
                    <SPLIT distance="700" swimtime="00:11:09.79" />
                    <SPLIT distance="750" swimtime="00:12:00.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="359" swimtime="00:00:40.83" resultid="1968" heatid="4647" lane="1" entrytime="00:00:44.45" />
                <RESULT eventid="1320" points="407" swimtime="00:01:15.56" resultid="1969" heatid="4668" lane="7" entrytime="00:01:17.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="366" swimtime="00:01:28.77" resultid="1970" heatid="4711" lane="8" entrytime="00:01:35.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="387" swimtime="00:03:13.23" resultid="1971" heatid="4748" lane="1" entrytime="00:03:24.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.48" />
                    <SPLIT distance="100" swimtime="00:01:34.01" />
                    <SPLIT distance="150" swimtime="00:02:23.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Chłąd" birthdate="2001-01-01" gender="M" nation="POL" athleteid="3627">
              <RESULTS>
                <RESULT eventid="1124" swimtime="00:02:44.92" resultid="3628" heatid="4626" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:17.01" />
                    <SPLIT distance="150" swimtime="00:02:06.74" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Przekroczony limit czasu" eventid="1182" status="OTL" swimtime="00:11:15.17" resultid="3629" heatid="4633" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                    <SPLIT distance="150" swimtime="00:01:56.88" />
                    <SPLIT distance="200" swimtime="00:02:39.40" />
                    <SPLIT distance="250" swimtime="00:03:22.36" />
                    <SPLIT distance="300" swimtime="00:04:05.54" />
                    <SPLIT distance="350" swimtime="00:04:48.73" />
                    <SPLIT distance="400" swimtime="00:05:32.41" />
                    <SPLIT distance="450" swimtime="00:06:15.34" />
                    <SPLIT distance="500" swimtime="00:06:58.86" />
                    <SPLIT distance="550" swimtime="00:07:42.38" />
                    <SPLIT distance="600" swimtime="00:08:26.48" />
                    <SPLIT distance="650" swimtime="00:09:10.09" />
                    <SPLIT distance="700" swimtime="00:09:53.80" />
                    <SPLIT distance="750" swimtime="00:10:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" swimtime="00:00:34.10" resultid="3630" heatid="4649" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1286" swimtime="00:03:15.69" resultid="3631" heatid="4655" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                    <SPLIT distance="100" swimtime="00:01:33.47" />
                    <SPLIT distance="150" swimtime="00:02:25.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" swimtime="00:01:15.61" resultid="3632" heatid="4712" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" swimtime="00:06:06.12" resultid="3633" heatid="4790" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:20.70" />
                    <SPLIT distance="150" swimtime="00:02:08.67" />
                    <SPLIT distance="200" swimtime="00:02:55.47" />
                    <SPLIT distance="250" swimtime="00:03:47.89" />
                    <SPLIT distance="300" swimtime="00:04:41.11" />
                    <SPLIT distance="350" swimtime="00:05:24.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Wilmowicz" birthdate="1979-01-01" gender="M" nation="POL" athleteid="4019">
              <RESULTS>
                <RESULT eventid="1090" points="501" swimtime="00:00:29.21" resultid="4020" heatid="4612" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1216" points="477" swimtime="00:21:00.28" resultid="4021" heatid="4639" lane="2" entrytime="00:20:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:01:54.36" />
                    <SPLIT distance="200" swimtime="00:02:35.58" />
                    <SPLIT distance="250" swimtime="00:03:17.28" />
                    <SPLIT distance="300" swimtime="00:03:59.10" />
                    <SPLIT distance="350" swimtime="00:04:40.62" />
                    <SPLIT distance="400" swimtime="00:05:23.01" />
                    <SPLIT distance="450" swimtime="00:06:05.23" />
                    <SPLIT distance="500" swimtime="00:06:47.36" />
                    <SPLIT distance="550" swimtime="00:07:29.59" />
                    <SPLIT distance="600" swimtime="00:08:11.90" />
                    <SPLIT distance="650" swimtime="00:08:54.42" />
                    <SPLIT distance="700" swimtime="00:09:36.93" />
                    <SPLIT distance="750" swimtime="00:10:19.15" />
                    <SPLIT distance="800" swimtime="00:11:01.72" />
                    <SPLIT distance="850" swimtime="00:11:44.67" />
                    <SPLIT distance="900" swimtime="00:12:27.57" />
                    <SPLIT distance="950" swimtime="00:13:10.29" />
                    <SPLIT distance="1000" swimtime="00:13:53.21" />
                    <SPLIT distance="1050" swimtime="00:14:35.96" />
                    <SPLIT distance="1100" swimtime="00:15:18.98" />
                    <SPLIT distance="1150" swimtime="00:16:02.20" />
                    <SPLIT distance="1200" swimtime="00:16:45.24" />
                    <SPLIT distance="1250" swimtime="00:17:29.45" />
                    <SPLIT distance="1300" swimtime="00:18:12.59" />
                    <SPLIT distance="1350" swimtime="00:18:55.37" />
                    <SPLIT distance="1400" swimtime="00:19:38.07" />
                    <SPLIT distance="1450" swimtime="00:20:20.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="510" swimtime="00:01:04.07" resultid="4022" heatid="4672" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="487" swimtime="00:02:24.37" resultid="4023" heatid="4724" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:08.65" />
                    <SPLIT distance="150" swimtime="00:01:46.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="488" swimtime="00:05:13.24" resultid="4024" heatid="4796" lane="1" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:13.23" />
                    <SPLIT distance="150" swimtime="00:01:53.42" />
                    <SPLIT distance="200" swimtime="00:02:33.88" />
                    <SPLIT distance="250" swimtime="00:03:14.80" />
                    <SPLIT distance="300" swimtime="00:03:55.34" />
                    <SPLIT distance="350" swimtime="00:04:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)." eventid="1422" status="DSQ" swimtime="00:01:22.33" resultid="4025" heatid="4692" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Krzekotowski" birthdate="1966-01-01" gender="M" nation="POL" athleteid="1944">
              <RESULTS>
                <RESULT eventid="1090" points="237" swimtime="00:00:39.46" resultid="1945" heatid="4605" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1124" points="196" swimtime="00:04:02.01" resultid="1946" heatid="4624" lane="0" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.95" />
                    <SPLIT distance="100" swimtime="00:02:04.24" />
                    <SPLIT distance="150" swimtime="00:03:07.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="228" swimtime="00:04:06.50" resultid="1947" heatid="4656" lane="8" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.98" />
                    <SPLIT distance="100" swimtime="00:01:58.52" />
                    <SPLIT distance="150" swimtime="00:03:01.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="127" swimtime="00:04:31.90" resultid="1948" heatid="4679" lane="7" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.86" />
                    <SPLIT distance="100" swimtime="00:02:07.13" />
                    <SPLIT distance="150" swimtime="00:03:19.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="224" swimtime="00:03:23.95" resultid="1949" heatid="4719" lane="5" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                    <SPLIT distance="100" swimtime="00:01:40.58" />
                    <SPLIT distance="150" swimtime="00:02:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="199" swimtime="00:08:28.96" resultid="1950" heatid="4789" lane="2" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.34" />
                    <SPLIT distance="100" swimtime="00:02:10.17" />
                    <SPLIT distance="150" swimtime="00:03:25.19" />
                    <SPLIT distance="200" swimtime="00:04:37.66" />
                    <SPLIT distance="250" swimtime="00:05:42.21" />
                    <SPLIT distance="300" swimtime="00:06:45.07" />
                    <SPLIT distance="350" swimtime="00:07:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="118" swimtime="00:02:03.40" resultid="1951" heatid="4738" lane="1" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="183" swimtime="00:07:41.78" resultid="1952" heatid="4801" lane="3" entrytime="00:07:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                    <SPLIT distance="100" swimtime="00:01:48.86" />
                    <SPLIT distance="150" swimtime="00:02:47.22" />
                    <SPLIT distance="200" swimtime="00:03:46.97" />
                    <SPLIT distance="250" swimtime="00:04:46.87" />
                    <SPLIT distance="300" swimtime="00:05:46.33" />
                    <SPLIT distance="350" swimtime="00:06:45.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Gorczyca" birthdate="1990-01-01" gender="M" nation="POL" athleteid="2652">
              <RESULTS>
                <RESULT eventid="1286" points="740" swimtime="00:02:32.58" resultid="2653" heatid="4658" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="817" swimtime="00:01:05.51" resultid="2654" heatid="4693" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1701" points="896" swimtime="00:00:28.77" resultid="2655" heatid="4762" lane="3" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Irena" lastname="Skowron" birthdate="1960-01-01" gender="F" nation="POL" athleteid="2031">
              <RESULTS>
                <RESULT comment="Przekroczony limit czasu" eventid="1199" status="OTL" swimtime="00:36:32.62" resultid="2032" heatid="4637" lane="2" entrytime="00:33:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.30" />
                    <SPLIT distance="100" swimtime="00:02:08.07" />
                    <SPLIT distance="150" swimtime="00:03:17.71" />
                    <SPLIT distance="200" swimtime="00:04:28.14" />
                    <SPLIT distance="250" swimtime="00:05:36.90" />
                    <SPLIT distance="300" swimtime="00:06:48.02" />
                    <SPLIT distance="350" swimtime="00:07:59.01" />
                    <SPLIT distance="400" swimtime="00:09:09.25" />
                    <SPLIT distance="450" swimtime="00:10:20.23" />
                    <SPLIT distance="500" swimtime="00:11:33.35" />
                    <SPLIT distance="550" swimtime="00:12:44.22" />
                    <SPLIT distance="600" swimtime="00:13:58.36" />
                    <SPLIT distance="650" swimtime="00:15:09.82" />
                    <SPLIT distance="700" swimtime="00:16:23.34" />
                    <SPLIT distance="750" swimtime="00:17:35.11" />
                    <SPLIT distance="800" swimtime="00:18:50.90" />
                    <SPLIT distance="850" swimtime="00:20:04.53" />
                    <SPLIT distance="900" swimtime="00:21:20.03" />
                    <SPLIT distance="950" swimtime="00:22:33.77" />
                    <SPLIT distance="1000" swimtime="00:23:49.13" />
                    <SPLIT distance="1050" swimtime="00:25:06.53" />
                    <SPLIT distance="1100" swimtime="00:26:23.36" />
                    <SPLIT distance="1150" swimtime="00:27:37.24" />
                    <SPLIT distance="1200" swimtime="00:28:54.81" />
                    <SPLIT distance="1250" swimtime="00:30:10.43" />
                    <SPLIT distance="1300" swimtime="00:31:28.95" />
                    <SPLIT distance="1350" swimtime="00:32:35.48" />
                    <SPLIT distance="1400" swimtime="00:34:03.87" />
                    <SPLIT distance="1450" swimtime="00:35:20.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="198" swimtime="00:02:22.43" resultid="2033" heatid="4685" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Płonka" birthdate="1948-01-01" gender="M" nation="POL" athleteid="1980">
              <RESULTS>
                <RESULT eventid="1124" points="156" swimtime="00:05:29.53" resultid="1981" heatid="4623" lane="1" entrytime="00:05:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.11" />
                    <SPLIT distance="100" swimtime="00:02:48.56" />
                    <SPLIT distance="150" swimtime="00:04:25.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="123" swimtime="00:06:29.03" resultid="1982" heatid="4655" lane="2" entrytime="00:05:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.31" />
                    <SPLIT distance="100" swimtime="00:03:11.99" />
                    <SPLIT distance="150" swimtime="00:04:53.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="105" swimtime="00:06:44.86" resultid="1983" heatid="4678" lane="4" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.41" />
                    <SPLIT distance="100" swimtime="00:03:19.23" />
                    <SPLIT distance="150" swimtime="00:05:10.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="158" swimtime="00:00:58.66" resultid="1984" heatid="4698" lane="8" entrytime="00:00:59.00" />
                <RESULT eventid="1524" points="96" swimtime="00:05:17.26" resultid="1985" heatid="4718" lane="5" entrytime="00:04:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.58" />
                    <SPLIT distance="100" swimtime="00:02:37.26" />
                    <SPLIT distance="150" swimtime="00:04:01.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="117" swimtime="00:02:44.53" resultid="1986" heatid="4738" lane="9" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="126" swimtime="00:10:33.11" resultid="1987" heatid="4802" lane="3" entrytime="00:11:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.87" />
                    <SPLIT distance="100" swimtime="00:02:31.17" />
                    <SPLIT distance="150" swimtime="00:03:53.37" />
                    <SPLIT distance="200" swimtime="00:05:15.65" />
                    <SPLIT distance="250" swimtime="00:06:37.21" />
                    <SPLIT distance="300" swimtime="00:07:59.29" />
                    <SPLIT distance="350" swimtime="00:09:19.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Poloch" birthdate="1983-01-01" gender="M" nation="POL" athleteid="4002">
              <RESULTS>
                <RESULT eventid="1090" points="372" swimtime="00:00:32.24" resultid="4003" heatid="4608" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1320" points="317" swimtime="00:01:15.10" resultid="4004" heatid="4666" lane="8" entrytime="00:01:35.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="219" swimtime="00:03:08.29" resultid="4005" heatid="4720" lane="9" entrytime="00:03:20.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:01:25.62" />
                    <SPLIT distance="150" swimtime="00:02:20.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="4006" heatid="4758" lane="0" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Gawkowski" birthdate="1958-01-01" gender="M" nation="POL" athleteid="2608">
              <RESULTS>
                <RESULT eventid="1090" points="309" swimtime="00:00:38.75" resultid="2609" heatid="4606" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1216" points="344" swimtime="00:27:54.25" resultid="2610" heatid="4638" lane="6" entrytime="00:27:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.68" />
                    <SPLIT distance="100" swimtime="00:01:44.71" />
                    <SPLIT distance="150" swimtime="00:02:40.04" />
                    <SPLIT distance="200" swimtime="00:03:36.54" />
                    <SPLIT distance="250" swimtime="00:04:33.70" />
                    <SPLIT distance="300" swimtime="00:05:30.88" />
                    <SPLIT distance="350" swimtime="00:06:26.74" />
                    <SPLIT distance="400" swimtime="00:07:23.42" />
                    <SPLIT distance="450" swimtime="00:08:19.79" />
                    <SPLIT distance="500" swimtime="00:09:16.11" />
                    <SPLIT distance="550" swimtime="00:10:13.25" />
                    <SPLIT distance="600" swimtime="00:11:09.35" />
                    <SPLIT distance="650" swimtime="00:12:06.21" />
                    <SPLIT distance="700" swimtime="00:13:02.58" />
                    <SPLIT distance="750" swimtime="00:13:59.42" />
                    <SPLIT distance="800" swimtime="00:14:55.30" />
                    <SPLIT distance="850" swimtime="00:15:51.52" />
                    <SPLIT distance="900" swimtime="00:16:47.54" />
                    <SPLIT distance="950" swimtime="00:17:43.53" />
                    <SPLIT distance="1000" swimtime="00:18:38.67" />
                    <SPLIT distance="1050" swimtime="00:19:33.79" />
                    <SPLIT distance="1100" swimtime="00:20:28.83" />
                    <SPLIT distance="1150" swimtime="00:21:25.31" />
                    <SPLIT distance="1200" swimtime="00:22:21.45" />
                    <SPLIT distance="1250" swimtime="00:23:17.57" />
                    <SPLIT distance="1300" swimtime="00:24:13.62" />
                    <SPLIT distance="1350" swimtime="00:25:10.08" />
                    <SPLIT distance="1400" swimtime="00:26:05.78" />
                    <SPLIT distance="1450" swimtime="00:27:01.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Woźniak" birthdate="1986-01-01" gender="M" nation="POL" athleteid="2665">
              <RESULTS>
                <RESULT eventid="1090" points="204" swimtime="00:00:38.62" resultid="2666" heatid="4606" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1320" points="172" swimtime="00:01:31.21" resultid="2667" heatid="4665" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kraśniewski" birthdate="1990-01-01" gender="M" nation="POL" athleteid="1988">
              <RESULTS>
                <RESULT eventid="1090" points="407" swimtime="00:00:29.84" resultid="1989" heatid="4612" lane="8" entrytime="00:00:29.53" />
                <RESULT eventid="1456" status="DNS" swimtime="00:00:00.00" resultid="1990" heatid="4701" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1524" points="362" swimtime="00:02:33.61" resultid="1991" heatid="4722" lane="7" entrytime="00:02:36.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:53.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="328" swimtime="00:05:45.18" resultid="1992" heatid="4798" lane="6" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                    <SPLIT distance="100" swimtime="00:01:20.58" />
                    <SPLIT distance="150" swimtime="00:02:03.95" />
                    <SPLIT distance="200" swimtime="00:02:48.04" />
                    <SPLIT distance="250" swimtime="00:03:32.14" />
                    <SPLIT distance="300" swimtime="00:04:17.07" />
                    <SPLIT distance="350" swimtime="00:05:02.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dagmara" lastname="Jankiewicz" birthdate="1984-01-01" gender="F" nation="POL" athleteid="3609">
              <RESULTS>
                <RESULT eventid="1303" points="187" swimtime="00:01:41.44" resultid="3610" heatid="4660" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K15 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="1684" status="DSQ" swimtime="00:00:51.68" resultid="3611" heatid="4752" lane="7" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Apolonia" lastname="Popławska" birthdate="2002-01-01" gender="F" nation="POL" athleteid="4007">
              <RESULTS>
                <RESULT eventid="1059" swimtime="00:00:29.73" resultid="4008" heatid="4601" lane="3" entrytime="00:00:29.17" />
                <RESULT eventid="1234" swimtime="00:00:35.47" resultid="4009" heatid="4643" lane="3" entrytime="00:00:33.50" />
                <RESULT eventid="1303" swimtime="00:01:06.23" resultid="4010" heatid="4663" lane="1" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" swimtime="00:00:32.08" resultid="4011" heatid="4697" lane="0" entrytime="00:00:31.67" />
                <RESULT eventid="1684" status="DNS" swimtime="00:00:00.00" resultid="4012" heatid="4755" lane="2" entrytime="00:00:36.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Lara" birthdate="1985-01-01" gender="F" nation="POL" athleteid="3992">
              <RESULTS>
                <RESULT eventid="1107" points="278" swimtime="00:03:36.03" resultid="3993" heatid="4619" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.42" />
                    <SPLIT distance="100" swimtime="00:01:52.56" />
                    <SPLIT distance="150" swimtime="00:02:50.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="362" swimtime="00:12:49.53" resultid="3994" heatid="4632" lane="9" entrytime="00:12:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="150" swimtime="00:02:10.60" />
                    <SPLIT distance="200" swimtime="00:02:58.30" />
                    <SPLIT distance="250" swimtime="00:03:46.64" />
                    <SPLIT distance="300" swimtime="00:04:35.84" />
                    <SPLIT distance="350" swimtime="00:05:24.92" />
                    <SPLIT distance="400" swimtime="00:06:14.22" />
                    <SPLIT distance="450" swimtime="00:07:03.38" />
                    <SPLIT distance="500" swimtime="00:07:53.06" />
                    <SPLIT distance="550" swimtime="00:08:42.42" />
                    <SPLIT distance="600" swimtime="00:09:32.34" />
                    <SPLIT distance="650" swimtime="00:10:22.11" />
                    <SPLIT distance="700" swimtime="00:11:12.26" />
                    <SPLIT distance="750" swimtime="00:12:01.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G7 - Pływak znajdował się w pozycji na piersiach po opuszczaniu ściany nawrotowej." eventid="1573" status="DSQ" swimtime="00:07:34.49" resultid="3995" heatid="4785" lane="8" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                    <SPLIT distance="100" swimtime="00:01:48.71" />
                    <SPLIT distance="150" swimtime="00:02:55.02" />
                    <SPLIT distance="200" swimtime="00:04:03.50" />
                    <SPLIT distance="250" swimtime="00:05:01.40" />
                    <SPLIT distance="300" swimtime="00:06:00.79" />
                    <SPLIT distance="350" swimtime="00:06:46.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="185" swimtime="00:01:48.83" resultid="3996" heatid="4735" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Rybicki" birthdate="1963-01-01" gender="M" nation="POL" athleteid="1962">
              <RESULTS>
                <RESULT eventid="1090" points="522" swimtime="00:00:31.33" resultid="1963" heatid="4609" lane="5" entrytime="00:00:31.30" />
                <RESULT eventid="1320" points="469" swimtime="00:01:14.20" resultid="1964" heatid="4669" lane="5" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Lipka" birthdate="1958-01-01" gender="M" nation="POL" athleteid="3997">
              <RESULTS>
                <RESULT eventid="1124" points="200" swimtime="00:04:07.92" resultid="3998" heatid="4624" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.71" />
                    <SPLIT distance="100" swimtime="00:02:01.74" />
                    <SPLIT distance="150" swimtime="00:03:13.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="304" swimtime="00:14:54.65" resultid="3999" heatid="4634" lane="0" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="100" swimtime="00:01:36.24" />
                    <SPLIT distance="150" swimtime="00:02:29.54" />
                    <SPLIT distance="200" swimtime="00:03:25.50" />
                    <SPLIT distance="250" swimtime="00:04:20.37" />
                    <SPLIT distance="300" swimtime="00:05:16.38" />
                    <SPLIT distance="350" swimtime="00:06:12.04" />
                    <SPLIT distance="400" swimtime="00:07:09.04" />
                    <SPLIT distance="450" swimtime="00:08:05.16" />
                    <SPLIT distance="500" swimtime="00:09:02.61" />
                    <SPLIT distance="550" swimtime="00:09:59.53" />
                    <SPLIT distance="600" swimtime="00:10:58.12" />
                    <SPLIT distance="650" swimtime="00:11:56.59" />
                    <SPLIT distance="700" swimtime="00:12:57.47" />
                    <SPLIT distance="750" swimtime="00:13:56.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="232" swimtime="00:08:29.57" resultid="4000" heatid="4789" lane="4" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.14" />
                    <SPLIT distance="100" swimtime="00:01:51.28" />
                    <SPLIT distance="150" swimtime="00:03:08.06" />
                    <SPLIT distance="200" swimtime="00:04:20.85" />
                    <SPLIT distance="250" swimtime="00:05:31.68" />
                    <SPLIT distance="300" swimtime="00:06:41.52" />
                    <SPLIT distance="350" swimtime="00:07:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="264" swimtime="00:01:42.55" resultid="4001" heatid="4739" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Miler" birthdate="2002-01-01" gender="M" nation="POL" athleteid="1955">
              <RESULTS>
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="1956" heatid="4647" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="1286" swimtime="00:03:33.37" resultid="1957" heatid="4655" lane="4" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="100" swimtime="00:01:40.94" />
                    <SPLIT distance="150" swimtime="00:02:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" swimtime="00:01:36.63" resultid="1958" heatid="4690" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" swimtime="00:00:34.22" resultid="1959" heatid="4700" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1667" status="DNS" swimtime="00:00:00.00" resultid="1960" heatid="4747" lane="8" entrytime="00:04:00.00" />
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="1961" heatid="4758" lane="9" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Walerzak" birthdate="1978-01-01" gender="F" nation="POL" athleteid="2627">
              <RESULTS>
                <RESULT eventid="1684" points="261" swimtime="00:00:52.50" resultid="2628" heatid="4753" lane="7" entrytime="00:00:47.08" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kędzior" birthdate="1973-01-01" gender="M" nation="POL" athleteid="2599">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="2600" heatid="4625" lane="0" entrytime="00:03:30.00" />
                <RESULT eventid="1182" points="305" swimtime="00:13:14.35" resultid="2601" heatid="4634" lane="3" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:26.07" />
                    <SPLIT distance="150" swimtime="00:02:14.53" />
                    <SPLIT distance="200" swimtime="00:03:05.43" />
                    <SPLIT distance="250" swimtime="00:03:56.67" />
                    <SPLIT distance="300" swimtime="00:04:48.44" />
                    <SPLIT distance="350" swimtime="00:05:39.16" />
                    <SPLIT distance="400" swimtime="00:06:30.34" />
                    <SPLIT distance="450" swimtime="00:07:22.33" />
                    <SPLIT distance="500" swimtime="00:08:14.97" />
                    <SPLIT distance="550" swimtime="00:09:06.61" />
                    <SPLIT distance="600" swimtime="00:09:56.92" />
                    <SPLIT distance="650" swimtime="00:10:46.47" />
                    <SPLIT distance="700" swimtime="00:11:36.96" />
                    <SPLIT distance="750" swimtime="00:12:26.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="379" swimtime="00:00:39.48" resultid="2602" heatid="4647" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1320" points="367" swimtime="00:01:15.61" resultid="2603" heatid="4669" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="275" swimtime="00:01:34.62" resultid="2604" heatid="4711" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="219" swimtime="00:07:53.69" resultid="2605" heatid="4788" lane="1" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.52" />
                    <SPLIT distance="100" swimtime="00:01:51.22" />
                    <SPLIT distance="150" swimtime="00:02:52.34" />
                    <SPLIT distance="200" swimtime="00:03:51.29" />
                    <SPLIT distance="250" swimtime="00:05:05.36" />
                    <SPLIT distance="300" swimtime="00:06:19.12" />
                    <SPLIT distance="350" swimtime="00:07:03.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="263" swimtime="00:03:29.85" resultid="2606" heatid="4748" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.53" />
                    <SPLIT distance="100" swimtime="00:01:43.10" />
                    <SPLIT distance="150" swimtime="00:02:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="321" swimtime="00:06:13.43" resultid="2607" heatid="4799" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="150" swimtime="00:02:08.91" />
                    <SPLIT distance="200" swimtime="00:02:57.20" />
                    <SPLIT distance="250" swimtime="00:03:45.66" />
                    <SPLIT distance="300" swimtime="00:04:35.29" />
                    <SPLIT distance="350" swimtime="00:05:24.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Szwolgin" birthdate="1943-01-01" gender="M" nation="POL" athleteid="4014">
              <RESULTS>
                <RESULT eventid="1124" points="233" swimtime="00:05:23.12" resultid="4015" heatid="4623" lane="5" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.12" />
                    <SPLIT distance="100" swimtime="00:02:43.24" />
                    <SPLIT distance="150" swimtime="00:04:12.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="377" swimtime="00:00:52.80" resultid="4016" heatid="4646" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1490" points="364" swimtime="00:02:00.96" resultid="4017" heatid="4710" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="348" swimtime="00:04:33.96" resultid="4018" heatid="4748" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.34" />
                    <SPLIT distance="100" swimtime="00:02:21.88" />
                    <SPLIT distance="150" swimtime="00:03:32.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Marszałek" birthdate="1954-01-01" gender="M" nation="POL" athleteid="1977">
              <RESULTS>
                <RESULT eventid="1124" points="178" swimtime="00:04:17.86" resultid="1978" heatid="4623" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.36" />
                    <SPLIT distance="100" swimtime="00:02:07.45" />
                    <SPLIT distance="150" swimtime="00:03:22.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="247" swimtime="00:15:58.08" resultid="1979" heatid="4633" lane="5" entrytime="00:15:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.59" />
                    <SPLIT distance="100" swimtime="00:01:55.57" />
                    <SPLIT distance="150" swimtime="00:02:56.15" />
                    <SPLIT distance="200" swimtime="00:03:57.31" />
                    <SPLIT distance="250" swimtime="00:04:57.61" />
                    <SPLIT distance="300" swimtime="00:05:58.95" />
                    <SPLIT distance="350" swimtime="00:06:58.25" />
                    <SPLIT distance="400" swimtime="00:07:59.82" />
                    <SPLIT distance="450" swimtime="00:08:59.35" />
                    <SPLIT distance="500" swimtime="00:10:00.92" />
                    <SPLIT distance="550" swimtime="00:11:00.48" />
                    <SPLIT distance="600" swimtime="00:12:02.54" />
                    <SPLIT distance="650" swimtime="00:13:02.19" />
                    <SPLIT distance="700" swimtime="00:14:03.75" />
                    <SPLIT distance="750" swimtime="00:15:01.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01713" nation="POL" region="13" clubid="2259" name="St. Pływackie MASTERS Olsztyn" shortname="MASTERS Olsztyn">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Konopacki" birthdate="1978-04-01" gender="M" nation="POL" license="501713700019" athleteid="3663">
              <RESULTS>
                <RESULT eventid="1090" points="593" swimtime="00:00:28.02" resultid="3664" heatid="4613" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1216" points="561" swimtime="00:20:10.55" resultid="3665" heatid="4639" lane="4" entrytime="00:19:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:14.88" />
                    <SPLIT distance="150" swimtime="00:01:55.22" />
                    <SPLIT distance="200" swimtime="00:02:35.15" />
                    <SPLIT distance="250" swimtime="00:03:15.54" />
                    <SPLIT distance="300" swimtime="00:03:56.41" />
                    <SPLIT distance="350" swimtime="00:04:36.98" />
                    <SPLIT distance="400" swimtime="00:05:17.20" />
                    <SPLIT distance="450" swimtime="00:05:58.23" />
                    <SPLIT distance="500" swimtime="00:06:38.57" />
                    <SPLIT distance="550" swimtime="00:07:18.93" />
                    <SPLIT distance="600" swimtime="00:07:59.73" />
                    <SPLIT distance="650" swimtime="00:08:40.26" />
                    <SPLIT distance="700" swimtime="00:09:20.89" />
                    <SPLIT distance="750" swimtime="00:10:01.45" />
                    <SPLIT distance="800" swimtime="00:10:41.90" />
                    <SPLIT distance="850" swimtime="00:11:22.66" />
                    <SPLIT distance="900" swimtime="00:12:03.18" />
                    <SPLIT distance="950" swimtime="00:12:43.71" />
                    <SPLIT distance="1000" swimtime="00:13:24.00" />
                    <SPLIT distance="1050" swimtime="00:14:04.70" />
                    <SPLIT distance="1100" swimtime="00:14:45.35" />
                    <SPLIT distance="1150" swimtime="00:15:25.60" />
                    <SPLIT distance="1200" swimtime="00:16:06.16" />
                    <SPLIT distance="1250" swimtime="00:16:46.91" />
                    <SPLIT distance="1300" swimtime="00:17:27.49" />
                    <SPLIT distance="1350" swimtime="00:18:08.37" />
                    <SPLIT distance="1400" swimtime="00:18:49.25" />
                    <SPLIT distance="1450" swimtime="00:19:29.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="538" swimtime="00:00:33.94" resultid="3666" heatid="4649" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1320" points="586" swimtime="00:01:02.40" resultid="3667" heatid="4673" lane="8" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="613" swimtime="00:02:18.61" resultid="3668" heatid="4724" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:43.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="533" swimtime="00:05:50.01" resultid="3669" heatid="4787" lane="7" entrytime="00:05:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:22.79" />
                    <SPLIT distance="150" swimtime="00:02:08.72" />
                    <SPLIT distance="200" swimtime="00:02:54.20" />
                    <SPLIT distance="250" swimtime="00:03:45.36" />
                    <SPLIT distance="300" swimtime="00:04:34.47" />
                    <SPLIT distance="350" swimtime="00:05:12.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="463" swimtime="00:02:50.01" resultid="3670" heatid="4749" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:23.28" />
                    <SPLIT distance="150" swimtime="00:02:07.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="592" swimtime="00:04:58.93" resultid="3671" heatid="4796" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="150" swimtime="00:01:47.98" />
                    <SPLIT distance="200" swimtime="00:02:27.04" />
                    <SPLIT distance="250" swimtime="00:03:06.25" />
                    <SPLIT distance="300" swimtime="00:03:45.83" />
                    <SPLIT distance="350" swimtime="00:04:24.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Gregorowicz" birthdate="1974-10-30" gender="M" nation="POL" license="101713700002" athleteid="3655">
              <RESULTS>
                <RESULT eventid="1090" points="690" swimtime="00:00:26.65" resultid="3656" heatid="4614" lane="6" entrytime="00:00:27.47" />
                <RESULT eventid="1182" points="687" swimtime="00:09:50.13" resultid="3657" heatid="4636" lane="2" entrytime="00:09:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:47.05" />
                    <SPLIT distance="200" swimtime="00:02:24.57" />
                    <SPLIT distance="250" swimtime="00:03:01.98" />
                    <SPLIT distance="300" swimtime="00:03:39.54" />
                    <SPLIT distance="350" swimtime="00:04:17.04" />
                    <SPLIT distance="400" swimtime="00:04:54.42" />
                    <SPLIT distance="450" swimtime="00:05:31.71" />
                    <SPLIT distance="500" swimtime="00:06:09.11" />
                    <SPLIT distance="550" swimtime="00:06:46.63" />
                    <SPLIT distance="600" swimtime="00:07:24.15" />
                    <SPLIT distance="650" swimtime="00:08:01.67" />
                    <SPLIT distance="700" swimtime="00:08:38.96" />
                    <SPLIT distance="750" swimtime="00:09:16.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="642" swimtime="00:02:27.13" resultid="3658" heatid="4681" lane="2" entrytime="00:02:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="719" swimtime="00:00:28.17" resultid="3659" heatid="4703" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="1597" points="666" swimtime="00:05:24.96" resultid="3660" heatid="4787" lane="2" entrytime="00:05:20.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:55.57" />
                    <SPLIT distance="200" swimtime="00:02:38.38" />
                    <SPLIT distance="250" swimtime="00:03:25.39" />
                    <SPLIT distance="300" swimtime="00:04:12.62" />
                    <SPLIT distance="350" swimtime="00:04:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="747" swimtime="00:01:02.65" resultid="3661" heatid="4741" lane="5" entrytime="00:01:04.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="700" swimtime="00:04:42.64" resultid="3662" heatid="4795" lane="2" entrytime="00:04:40.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:07.23" />
                    <SPLIT distance="150" swimtime="00:01:42.93" />
                    <SPLIT distance="200" swimtime="00:02:18.93" />
                    <SPLIT distance="250" swimtime="00:02:55.16" />
                    <SPLIT distance="300" swimtime="00:03:31.30" />
                    <SPLIT distance="350" swimtime="00:04:07.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kieres" birthdate="1984-06-13" gender="M" nation="POL" license="101713700001" athleteid="3686">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="3687" heatid="4626" lane="6" entrytime="00:02:50.00" />
                <RESULT eventid="1286" points="378" swimtime="00:03:13.97" resultid="3688" heatid="4657" lane="3" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="100" swimtime="00:01:30.12" />
                    <SPLIT distance="150" swimtime="00:02:21.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="317" swimtime="00:02:59.70" resultid="3689" heatid="4681" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:19.03" />
                    <SPLIT distance="150" swimtime="00:02:08.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="335" swimtime="00:01:29.78" resultid="3690" heatid="4692" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="369" swimtime="00:06:25.56" resultid="3691" heatid="4787" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:23.94" />
                    <SPLIT distance="150" swimtime="00:02:15.79" />
                    <SPLIT distance="200" swimtime="00:03:07.65" />
                    <SPLIT distance="250" swimtime="00:04:02.46" />
                    <SPLIT distance="300" swimtime="00:04:57.59" />
                    <SPLIT distance="350" swimtime="00:05:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" status="DNS" swimtime="00:00:00.00" resultid="3692" heatid="4740" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="3693" heatid="4759" lane="4" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Matusiak vel Matuszewski" birthdate="1974-06-25" gender="M" nation="POL" license="501713700004" athleteid="3677">
              <RESULTS>
                <RESULT eventid="1090" points="324" swimtime="00:00:34.27" resultid="3678" heatid="4608" lane="9" entrytime="00:00:34.13" />
                <RESULT eventid="1182" status="DNS" swimtime="00:00:00.00" resultid="3679" heatid="4635" lane="8" entrytime="00:11:47.93" />
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="3680" heatid="4647" lane="2" entrytime="00:00:42.13" />
                <RESULT eventid="1320" points="306" swimtime="00:01:17.49" resultid="3681" heatid="4669" lane="3" entrytime="00:01:14.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" status="DNS" swimtime="00:00:00.00" resultid="3682" heatid="4699" lane="1" entrytime="00:00:40.45" />
                <RESULT eventid="1524" points="355" swimtime="00:02:46.29" resultid="3683" heatid="4722" lane="9" entrytime="00:02:41.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:20.19" />
                    <SPLIT distance="150" swimtime="00:02:03.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" status="DNS" swimtime="00:00:00.00" resultid="3684" heatid="4748" lane="2" entrytime="00:03:16.90" />
                <RESULT eventid="1766" points="342" swimtime="00:05:58.88" resultid="3685" heatid="4798" lane="1" entrytime="00:05:46.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:01:24.82" />
                    <SPLIT distance="150" swimtime="00:02:10.28" />
                    <SPLIT distance="200" swimtime="00:02:56.20" />
                    <SPLIT distance="250" swimtime="00:03:42.70" />
                    <SPLIT distance="300" swimtime="00:04:29.03" />
                    <SPLIT distance="350" swimtime="00:05:14.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Mówiński" birthdate="1969-09-01" gender="M" nation="POL" license="501713700007" athleteid="3700">
              <RESULTS>
                <RESULT eventid="1182" points="412" swimtime="00:11:59.05" resultid="3701" heatid="4635" lane="9" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:01:24.63" />
                    <SPLIT distance="150" swimtime="00:02:09.60" />
                    <SPLIT distance="200" swimtime="00:02:54.29" />
                    <SPLIT distance="250" swimtime="00:03:39.66" />
                    <SPLIT distance="300" swimtime="00:04:25.65" />
                    <SPLIT distance="350" swimtime="00:05:11.29" />
                    <SPLIT distance="400" swimtime="00:05:56.92" />
                    <SPLIT distance="450" swimtime="00:06:42.65" />
                    <SPLIT distance="500" swimtime="00:07:28.60" />
                    <SPLIT distance="550" swimtime="00:08:13.56" />
                    <SPLIT distance="600" swimtime="00:08:59.25" />
                    <SPLIT distance="650" swimtime="00:09:44.59" />
                    <SPLIT distance="700" swimtime="00:10:30.65" />
                    <SPLIT distance="750" swimtime="00:11:16.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="340" swimtime="00:03:10.89" resultid="3702" heatid="4680" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:02:22.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="399" swimtime="00:02:41.09" resultid="3703" heatid="4721" lane="5" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:01.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="305" swimtime="00:01:24.99" resultid="3704" heatid="4739" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="400" swimtime="00:05:47.10" resultid="3705" heatid="4798" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:22.41" />
                    <SPLIT distance="150" swimtime="00:02:06.48" />
                    <SPLIT distance="200" swimtime="00:02:51.48" />
                    <SPLIT distance="250" swimtime="00:03:36.33" />
                    <SPLIT distance="300" swimtime="00:04:21.02" />
                    <SPLIT distance="350" swimtime="00:05:05.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jowita" lastname="Kucharska" birthdate="1980-02-15" gender="F" nation="POL" license="501713600018" athleteid="3649">
              <RESULTS>
                <RESULT eventid="1059" points="445" swimtime="00:00:34.63" resultid="3650" heatid="4599" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1234" points="350" swimtime="00:00:42.00" resultid="3651" heatid="4642" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1303" status="DNS" swimtime="00:00:00.00" resultid="3652" heatid="4661" lane="2" entrytime="00:01:18.00" />
                <RESULT eventid="1473" points="320" swimtime="00:01:34.50" resultid="3653" heatid="4707" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="312" swimtime="00:03:30.98" resultid="3654" heatid="4744" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                    <SPLIT distance="100" swimtime="00:01:43.10" />
                    <SPLIT distance="150" swimtime="00:02:38.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Łuczak" birthdate="1978-03-18" gender="M" nation="POL" license="501713700016" athleteid="3672">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="3673" heatid="4611" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1286" points="363" swimtime="00:03:15.31" resultid="3674" heatid="4657" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                    <SPLIT distance="100" swimtime="00:01:36.63" />
                    <SPLIT distance="150" swimtime="00:02:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="457" swimtime="00:01:24.05" resultid="3675" heatid="4692" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="499" swimtime="00:00:36.83" resultid="3676" heatid="4760" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oriana" lastname="Kowalińska" birthdate="1993-03-19" gender="F" nation="POL" license="101713600052" athleteid="3694">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1158" points="576" swimtime="00:10:32.62" resultid="3695" heatid="4632" lane="4" entrytime="00:10:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:01:15.85" />
                    <SPLIT distance="150" swimtime="00:01:55.05" />
                    <SPLIT distance="200" swimtime="00:02:34.88" />
                    <SPLIT distance="250" swimtime="00:03:11.57" />
                    <SPLIT distance="300" swimtime="00:03:53.89" />
                    <SPLIT distance="350" swimtime="00:04:33.56" />
                    <SPLIT distance="400" swimtime="00:05:13.05" />
                    <SPLIT distance="450" swimtime="00:05:50.20" />
                    <SPLIT distance="500" swimtime="00:06:33.11" />
                    <SPLIT distance="550" swimtime="00:07:13.20" />
                    <SPLIT distance="600" swimtime="00:07:53.35" />
                    <SPLIT distance="650" swimtime="00:08:33.89" />
                    <SPLIT distance="700" swimtime="00:09:14.18" />
                    <SPLIT distance="750" swimtime="00:09:54.55" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1337" points="608" swimtime="00:02:37.64" resultid="3696" heatid="4677" lane="4" entrytime="00:02:35.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                    <SPLIT distance="150" swimtime="00:01:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="651" swimtime="00:05:41.61" resultid="3697" heatid="4785" lane="3" entrytime="00:05:40.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:02:00.40" />
                    <SPLIT distance="200" swimtime="00:02:44.97" />
                    <SPLIT distance="250" swimtime="00:03:35.36" />
                    <SPLIT distance="300" swimtime="00:04:24.78" />
                    <SPLIT distance="350" swimtime="00:05:04.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="557" swimtime="00:01:11.44" resultid="3698" heatid="4736" lane="5" entrytime="00:01:10.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="575" swimtime="00:05:10.92" resultid="3699" heatid="4791" lane="3" entrytime="00:05:05.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:16.49" />
                    <SPLIT distance="150" swimtime="00:01:55.79" />
                    <SPLIT distance="200" swimtime="00:02:35.23" />
                    <SPLIT distance="250" swimtime="00:03:14.67" />
                    <SPLIT distance="300" swimtime="00:03:53.95" />
                    <SPLIT distance="350" swimtime="00:04:33.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Lach" birthdate="1978-04-09" gender="F" nation="POL" athleteid="2260">
              <RESULTS>
                <RESULT eventid="1059" points="174" swimtime="00:00:47.54" resultid="2261" heatid="4597" lane="8" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" status="DNS" swimtime="00:00:00.00" resultid="3707" heatid="4683" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" status="DNS" swimtime="00:00:00.00" resultid="3708" heatid="4727" lane="8">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1141" status="DNS" swimtime="00:00:00.00" resultid="3706" heatid="4629" lane="7">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1718" status="DNS" swimtime="00:00:00.00" resultid="3709" heatid="4763" lane="4" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00908" nation="POL" region="08" clubid="3009" name="MOTYL MASTERS Stalowa Wola">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Petecka" birthdate="1967-04-17" gender="F" nation="POL" athleteid="3010">
              <RESULTS>
                <RESULT eventid="1059" points="441" swimtime="00:00:37.09" resultid="3011" heatid="4599" lane="9" entrytime="00:00:36.80" />
                <RESULT eventid="1107" points="434" swimtime="00:03:20.03" resultid="3012" heatid="4619" lane="4" entrytime="00:03:19.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:38.52" />
                    <SPLIT distance="150" swimtime="00:02:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="523" swimtime="00:03:41.88" resultid="3013" heatid="4653" lane="2" entrytime="00:03:43.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.51" />
                    <SPLIT distance="100" swimtime="00:01:48.65" />
                    <SPLIT distance="150" swimtime="00:02:45.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="422" swimtime="00:01:46.51" resultid="3014" heatid="4686" lane="4" entrytime="00:01:47.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="420" swimtime="00:00:40.74" resultid="3015" heatid="4695" lane="8" entrytime="00:00:41.89" />
                <RESULT eventid="1615" points="283" swimtime="00:01:44.69" resultid="3016" heatid="4735" lane="4" entrytime="00:01:39.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="406" swimtime="00:00:48.51" resultid="3017" heatid="4753" lane="0" entrytime="00:00:48.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arkadiusz" lastname="Berwecki" birthdate="1973-01-14" gender="M" nation="POL" athleteid="3024">
              <RESULTS>
                <RESULT eventid="1124" points="712" swimtime="00:02:26.86" resultid="3025" heatid="4628" lane="1" entrytime="00:02:25.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="100" swimtime="00:01:09.38" />
                    <SPLIT distance="150" swimtime="00:01:51.22" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1354" points="702" swimtime="00:02:29.90" resultid="3026" heatid="4681" lane="3" entrytime="00:02:26.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                    <SPLIT distance="150" swimtime="00:01:50.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="755" swimtime="00:00:28.42" resultid="3027" heatid="4704" lane="8" entrytime="00:00:28.19" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1524" points="757" swimtime="00:02:10.12" resultid="3028" heatid="4725" lane="0" entrytime="00:02:09.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:04.91" />
                    <SPLIT distance="150" swimtime="00:01:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1633" points="772" swimtime="00:01:02.37" resultid="3029" heatid="4742" lane="7" entrytime="00:01:02.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1766" points="745" swimtime="00:04:42.29" resultid="3030" heatid="4795" lane="6" entrytime="00:04:39.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:07.01" />
                    <SPLIT distance="150" swimtime="00:01:43.26" />
                    <SPLIT distance="200" swimtime="00:02:19.99" />
                    <SPLIT distance="250" swimtime="00:02:56.35" />
                    <SPLIT distance="300" swimtime="00:03:33.14" />
                    <SPLIT distance="350" swimtime="00:04:09.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Lorkowski" birthdate="1960-02-27" gender="M" nation="POL" athleteid="3031">
              <RESULTS>
                <RESULT eventid="1090" points="456" swimtime="00:00:32.76" resultid="3032" heatid="4609" lane="2" entrytime="00:00:31.89" />
                <RESULT eventid="1124" points="452" swimtime="00:03:04.91" resultid="3033" heatid="4625" lane="6" entrytime="00:03:05.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:27.85" />
                    <SPLIT distance="150" swimtime="00:02:24.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3034" heatid="4669" lane="2" entrytime="00:01:14.97" />
                <RESULT comment="M11 - Pływak dotknął ścianę nierównocześnie dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="1354" status="DSQ" swimtime="00:03:31.58" resultid="3035" heatid="4680" lane="8" entrytime="00:03:38.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                    <SPLIT distance="100" swimtime="00:01:36.97" />
                    <SPLIT distance="150" swimtime="00:02:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" status="DNS" swimtime="00:00:00.00" resultid="3036" heatid="4721" lane="3" entrytime="00:02:48.12" />
                <RESULT eventid="1597" points="453" swimtime="00:06:41.06" resultid="3037" heatid="4788" lane="3" entrytime="00:06:47.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:01:33.15" />
                    <SPLIT distance="150" swimtime="00:02:24.23" />
                    <SPLIT distance="200" swimtime="00:03:14.79" />
                    <SPLIT distance="250" swimtime="00:04:13.97" />
                    <SPLIT distance="300" swimtime="00:05:11.98" />
                    <SPLIT distance="350" swimtime="00:05:58.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="466" swimtime="00:03:08.40" resultid="3038" heatid="4748" lane="5" entrytime="00:03:07.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.57" />
                    <SPLIT distance="100" swimtime="00:01:30.69" />
                    <SPLIT distance="150" swimtime="00:02:20.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="3039" heatid="4798" lane="9" entrytime="00:05:54.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Baran" birthdate="1975-03-19" gender="M" nation="POL" athleteid="3018">
              <RESULTS>
                <RESULT eventid="1090" points="579" swimtime="00:00:28.24" resultid="3019" heatid="4614" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1252" points="665" swimtime="00:00:31.64" resultid="3020" heatid="4650" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="1354" points="420" swimtime="00:02:49.48" resultid="3021" heatid="4680" lane="3" entrytime="00:03:02.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:24.12" />
                    <SPLIT distance="150" swimtime="00:02:10.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="651" swimtime="00:01:09.37" resultid="3022" heatid="4713" lane="8" entrytime="00:01:08.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="555" swimtime="00:02:40.02" resultid="3023" heatid="4749" lane="4" entrytime="00:02:38.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:16.96" />
                    <SPLIT distance="150" swimtime="00:01:59.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02207" nation="POL" region="07" clubid="1903" name="MASTERS Zdzieszowice">
          <ATHLETES>
            <ATHLETE firstname="Dorota" lastname="Woźniak" birthdate="1973-09-18" gender="F" nation="POL" athleteid="1904">
              <RESULTS>
                <RESULT eventid="1234" points="451" swimtime="00:00:41.17" resultid="1905" heatid="4642" lane="3" entrytime="00:00:37.11" />
                <RESULT eventid="1337" points="390" swimtime="00:03:27.28" resultid="1906" heatid="4677" lane="7" entrytime="00:03:13.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                    <SPLIT distance="100" swimtime="00:01:38.44" />
                    <SPLIT distance="150" swimtime="00:02:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="444" swimtime="00:01:29.31" resultid="1907" heatid="4708" lane="0" entrytime="00:01:24.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="437" swimtime="00:07:02.39" resultid="1908" heatid="4785" lane="2" entrytime="00:06:12.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:38.47" />
                    <SPLIT distance="150" swimtime="00:02:32.26" />
                    <SPLIT distance="200" swimtime="00:03:25.13" />
                    <SPLIT distance="250" swimtime="00:04:25.99" />
                    <SPLIT distance="300" swimtime="00:05:26.80" />
                    <SPLIT distance="350" swimtime="00:06:15.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="422" swimtime="00:03:15.35" resultid="1909" heatid="4745" lane="9" entrytime="00:03:15.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:34.80" />
                    <SPLIT distance="150" swimtime="00:02:26.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sasha" lastname="Broshevan" birthdate="1986-10-15" gender="M" nation="POL" athleteid="3004">
              <RESULTS>
                <RESULT eventid="1090" points="509" swimtime="00:00:28.50" resultid="3005" heatid="4613" lane="1" entrytime="00:00:28.20" />
                <RESULT eventid="1252" points="415" swimtime="00:00:35.09" resultid="3006" heatid="4649" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1456" points="493" swimtime="00:00:30.55" resultid="3007" heatid="4703" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1701" points="387" swimtime="00:00:38.87" resultid="3008" heatid="4760" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01610" nation="POL" region="10" clubid="2190" name="MASTERS Gdynia">
          <ATHLETES>
            <ATHLETE firstname="Grażyna" lastname="Heisler" birthdate="1951-01-01" gender="F" nation="POL" athleteid="2198">
              <RESULTS>
                <RESULT eventid="1059" points="317" swimtime="00:00:45.03" resultid="2199" heatid="4597" lane="3" entrytime="00:00:48.00" />
                <RESULT eventid="1404" points="304" swimtime="00:02:22.64" resultid="2200" heatid="4685" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="190" swimtime="00:02:14.26" resultid="2201" heatid="4706" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="179" swimtime="00:05:00.25" resultid="2202" heatid="4744" lane="8" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.71" />
                    <SPLIT distance="100" swimtime="00:02:25.69" />
                    <SPLIT distance="150" swimtime="00:03:46.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="297" swimtime="00:01:02.39" resultid="2203" heatid="4751" lane="4" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Gorbaczow" birthdate="1958-01-01" gender="M" nation="POL" athleteid="2209">
              <RESULTS>
                <RESULT eventid="1090" points="645" swimtime="00:00:30.32" resultid="2210" heatid="4607" lane="4" entrytime="00:00:34.20" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1124" points="528" swimtime="00:02:59.67" resultid="2211" heatid="4625" lane="5" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:29.19" />
                    <SPLIT distance="150" swimtime="00:02:21.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1252" points="633" swimtime="00:00:36.04" resultid="2212" heatid="4649" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1320" points="673" swimtime="00:01:07.88" resultid="2213" heatid="4671" lane="8" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1456" points="685" swimtime="00:00:32.18" resultid="2214" heatid="4702" lane="7" entrytime="00:00:31.10" />
                <RESULT eventid="1524" points="528" swimtime="00:02:40.02" resultid="2215" heatid="4722" lane="3" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                    <SPLIT distance="150" swimtime="00:02:00.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Boboli" birthdate="1948-01-01" gender="M" nation="POL" athleteid="2204">
              <RESULTS>
                <RESULT eventid="1090" points="393" swimtime="00:00:39.84" resultid="2205" heatid="4606" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1252" points="175" swimtime="00:01:01.54" resultid="2206" heatid="4646" lane="9" entrytime="00:01:00.00" />
                <RESULT eventid="1456" points="179" swimtime="00:00:56.29" resultid="2207" heatid="4699" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="1701" points="101" swimtime="00:01:21.72" resultid="2208" heatid="4757" lane="8" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Skwarło" birthdate="1939-01-01" gender="M" nation="POL" athleteid="2191">
              <RESULTS>
                <RESULT eventid="1090" points="158" swimtime="00:00:59.05" resultid="2192" heatid="4604" lane="5" entrytime="00:00:54.00" />
                <RESULT eventid="1252" points="215" swimtime="00:01:03.63" resultid="2193" heatid="4645" lane="5" entrytime="00:01:03.50" />
                <RESULT eventid="1286" points="244" swimtime="00:05:31.99" resultid="2194" heatid="4655" lane="6" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.81" />
                    <SPLIT distance="100" swimtime="00:02:38.25" />
                    <SPLIT distance="150" swimtime="00:04:08.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="222" swimtime="00:02:35.84" resultid="2195" heatid="4690" lane="7" entrytime="00:02:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="186" swimtime="00:02:31.35" resultid="2196" heatid="4709" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="281" swimtime="00:01:03.57" resultid="2197" heatid="4757" lane="2" entrytime="00:00:57.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Gorbaczow" birthdate="1987-01-01" gender="M" nation="POL" athleteid="2216">
              <RESULTS>
                <RESULT eventid="1090" points="382" swimtime="00:00:31.35" resultid="2217" heatid="4609" lane="4" entrytime="00:00:31.20" />
                <RESULT eventid="1320" points="315" swimtime="00:01:14.60" resultid="2218" heatid="4670" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="276" swimtime="00:00:37.04" resultid="2219" heatid="4700" lane="8" entrytime="00:00:37.10" />
                <RESULT eventid="1524" points="217" swimtime="00:03:07.68" resultid="2220" heatid="4720" lane="5" entrytime="00:03:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                    <SPLIT distance="150" swimtime="00:02:22.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="281" swimtime="00:02:59.21" resultid="2221" heatid="4683" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                    <SPLIT distance="150" swimtime="00:02:18.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2216" number="1" />
                    <RELAYPOSITION athleteid="2191" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2209" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2204" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="253" swimtime="00:02:41.74" resultid="2222" heatid="4727" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                    <SPLIT distance="150" swimtime="00:02:12.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2216" number="1" />
                    <RELAYPOSITION athleteid="2191" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2209" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="2204" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02602" nation="POL" region="02" clubid="2280" name="MULTISPORT TEAM Toruń">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Lietz" birthdate="1952-04-23" gender="M" nation="POL" athleteid="2281">
              <RESULTS>
                <RESULT eventid="1090" points="505" swimtime="00:00:34.78" resultid="2282" heatid="4607" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1182" points="392" swimtime="00:14:31.25" resultid="2283" heatid="4634" lane="9" entrytime="00:14:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.96" />
                    <SPLIT distance="100" swimtime="00:01:40.77" />
                    <SPLIT distance="150" swimtime="00:02:34.98" />
                    <SPLIT distance="200" swimtime="00:03:29.84" />
                    <SPLIT distance="250" swimtime="00:04:24.99" />
                    <SPLIT distance="300" swimtime="00:05:20.72" />
                    <SPLIT distance="350" swimtime="00:06:17.48" />
                    <SPLIT distance="400" swimtime="00:07:14.57" />
                    <SPLIT distance="450" swimtime="00:08:11.06" />
                    <SPLIT distance="500" swimtime="00:09:08.23" />
                    <SPLIT distance="550" swimtime="00:10:04.70" />
                    <SPLIT distance="600" swimtime="00:11:00.00" />
                    <SPLIT distance="650" swimtime="00:11:54.56" />
                    <SPLIT distance="700" swimtime="00:12:48.65" />
                    <SPLIT distance="750" swimtime="00:13:40.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="484" swimtime="00:01:20.60" resultid="2284" heatid="4668" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="437" swimtime="00:00:39.49" resultid="2285" heatid="4699" lane="6" entrytime="00:00:39.10" />
                <RESULT eventid="1524" points="454" swimtime="00:03:06.41" resultid="2286" heatid="4721" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                    <SPLIT distance="100" swimtime="00:01:32.06" />
                    <SPLIT distance="150" swimtime="00:02:21.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="411" swimtime="00:06:48.01" resultid="2287" heatid="4800" lane="5" entrytime="00:06:35.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:35.65" />
                    <SPLIT distance="150" swimtime="00:02:28.22" />
                    <SPLIT distance="200" swimtime="00:03:22.35" />
                    <SPLIT distance="250" swimtime="00:04:16.08" />
                    <SPLIT distance="300" swimtime="00:05:09.39" />
                    <SPLIT distance="350" swimtime="00:06:01.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12914" nation="POL" region="14" clubid="3314" name="WATER SQUAD Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Fluder" birthdate="1986-03-01" gender="M" nation="POL" license="512914700007" athleteid="3387">
              <RESULTS>
                <RESULT eventid="1090" points="650" swimtime="00:00:26.27" resultid="3388" heatid="4615" lane="7" entrytime="00:00:26.40" />
                <RESULT eventid="1320" points="687" swimtime="00:00:57.53" resultid="3389" heatid="4674" lane="3" entrytime="00:00:56.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="693" swimtime="00:02:07.47" resultid="3390" heatid="4725" lane="2" entrytime="00:02:07.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                    <SPLIT distance="100" swimtime="00:01:00.96" />
                    <SPLIT distance="150" swimtime="00:01:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="733" swimtime="00:04:32.73" resultid="3391" heatid="4795" lane="3" entrytime="00:04:32.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:40.12" />
                    <SPLIT distance="200" swimtime="00:02:15.09" />
                    <SPLIT distance="250" swimtime="00:02:49.69" />
                    <SPLIT distance="300" swimtime="00:03:24.68" />
                    <SPLIT distance="350" swimtime="00:03:59.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Markowski" birthdate="1976-01-04" gender="M" nation="POL" license="512914700011" athleteid="3392">
              <RESULTS>
                <RESULT eventid="1124" points="505" swimtime="00:02:43.30" resultid="3393" heatid="4627" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="150" swimtime="00:02:04.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="511" swimtime="00:01:15.21" resultid="3394" heatid="4712" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="487" swimtime="00:06:00.55" resultid="3395" heatid="4787" lane="1" entrytime="00:05:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:01:22.78" />
                    <SPLIT distance="150" swimtime="00:02:10.03" />
                    <SPLIT distance="200" swimtime="00:02:55.29" />
                    <SPLIT distance="250" swimtime="00:03:46.37" />
                    <SPLIT distance="300" swimtime="00:04:37.33" />
                    <SPLIT distance="350" swimtime="00:05:20.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="560" swimtime="00:01:08.96" resultid="3396" heatid="4741" lane="9" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="503" swimtime="00:02:45.41" resultid="3397" heatid="4749" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:21.56" />
                    <SPLIT distance="150" swimtime="00:02:04.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Mikicin" birthdate="1993-10-18" gender="M" nation="POL" license="112914700058" athleteid="3353">
              <RESULTS>
                <RESULT eventid="1090" points="684" swimtime="00:00:25.11" resultid="3354" heatid="4615" lane="5" entrytime="00:00:26.00" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1252" points="835" swimtime="00:00:27.57" resultid="3355" heatid="4651" lane="2" entrytime="00:00:28.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arkadiusz" lastname="Aptewicz" birthdate="1993-12-20" gender="M" nation="POL" license="112914700053" athleteid="3315">
              <RESULTS>
                <RESULT eventid="1124" points="715" swimtime="00:02:16.62" resultid="3316" heatid="4628" lane="5" entrytime="00:02:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="100" swimtime="00:01:04.47" />
                    <SPLIT distance="150" swimtime="00:01:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="788" swimtime="00:02:29.44" resultid="3317" heatid="4658" lane="4" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                    <SPLIT distance="150" swimtime="00:01:50.33" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1597" points="675" swimtime="00:04:57.21" resultid="3318" heatid="4787" lane="5" entrytime="00:04:51.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="150" swimtime="00:01:48.74" />
                    <SPLIT distance="200" swimtime="00:02:28.73" />
                    <SPLIT distance="250" swimtime="00:03:09.12" />
                    <SPLIT distance="300" swimtime="00:03:50.05" />
                    <SPLIT distance="350" swimtime="00:04:24.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="688" swimtime="00:00:31.41" resultid="3319" heatid="4762" lane="0" entrytime="00:00:31.50" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1766" points="713" swimtime="00:04:26.53" resultid="3320" heatid="4795" lane="4" entrytime="00:04:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                    <SPLIT distance="100" swimtime="00:01:02.81" />
                    <SPLIT distance="150" swimtime="00:01:37.20" />
                    <SPLIT distance="200" swimtime="00:02:11.51" />
                    <SPLIT distance="250" swimtime="00:02:45.73" />
                    <SPLIT distance="300" swimtime="00:03:20.22" />
                    <SPLIT distance="350" swimtime="00:03:54.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Dąbrowska" birthdate="1987-05-20" gender="F" nation="POL" license="512914600064" athleteid="3321">
              <RESULTS>
                <RESULT eventid="1059" points="265" swimtime="00:00:40.44" resultid="3322" heatid="4598" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="3323" heatid="4619" lane="0" entrytime="00:04:00.00" />
                <RESULT eventid="1234" points="148" swimtime="00:00:54.12" resultid="3324" heatid="4641" lane="9" entrytime="00:00:54.00" />
                <RESULT eventid="1303" points="221" swimtime="00:01:36.04" resultid="3325" heatid="4660" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="154" swimtime="00:00:51.20" resultid="3326" heatid="4694" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1507" points="187" swimtime="00:03:40.21" resultid="3327" heatid="4715" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.15" />
                    <SPLIT distance="100" swimtime="00:01:44.52" />
                    <SPLIT distance="150" swimtime="00:02:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="3328" heatid="4735" lane="5" entrytime="00:01:40.00" />
                <RESULT eventid="1742" status="DNS" swimtime="00:00:00.00" resultid="3329" heatid="4793" lane="0" entrytime="00:07:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Hebel" birthdate="1987-06-22" gender="F" nation="POL" license="512914600059" athleteid="3405">
              <RESULTS>
                <RESULT eventid="1059" points="424" swimtime="00:00:34.58" resultid="3406" heatid="4599" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1269" points="266" swimtime="00:04:01.54" resultid="3407" heatid="4652" lane="5" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.55" />
                    <SPLIT distance="100" swimtime="00:01:54.68" />
                    <SPLIT distance="150" swimtime="00:02:58.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="415" swimtime="00:01:17.83" resultid="3408" heatid="4661" lane="3" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="271" swimtime="00:01:35.33" resultid="3409" heatid="4707" lane="5" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="347" swimtime="00:02:59.18" resultid="3410" heatid="4716" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:01:24.96" />
                    <SPLIT distance="150" swimtime="00:02:12.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="343" swimtime="00:03:17.35" resultid="3411" heatid="4745" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:35.70" />
                    <SPLIT distance="150" swimtime="00:02:26.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Solis" birthdate="1970-07-15" gender="F" nation="POL" athleteid="3493">
              <RESULTS>
                <RESULT eventid="1059" points="460" swimtime="00:00:35.07" resultid="3494" heatid="4598" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1234" points="337" swimtime="00:00:45.36" resultid="3495" heatid="4641" lane="6" entrytime="00:00:46.00" />
                <RESULT eventid="1684" points="358" swimtime="00:00:48.13" resultid="3496" heatid="4752" lane="2" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Brożyna" birthdate="1980-04-28" gender="M" nation="POL" license="512914700006" athleteid="3398">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="3399" heatid="4627" lane="9" entrytime="00:02:45.00" />
                <RESULT eventid="1252" points="500" swimtime="00:00:34.16" resultid="3400" heatid="4649" lane="6" entrytime="00:00:34.40" />
                <RESULT eventid="1490" points="500" swimtime="00:01:13.60" resultid="3401" heatid="4712" lane="1" entrytime="00:01:16.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="449" swimtime="00:06:09.48" resultid="3402" heatid="4788" lane="4" entrytime="00:06:03.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:30.00" />
                    <SPLIT distance="150" swimtime="00:02:14.05" />
                    <SPLIT distance="200" swimtime="00:02:58.29" />
                    <SPLIT distance="250" swimtime="00:03:51.84" />
                    <SPLIT distance="300" swimtime="00:04:45.96" />
                    <SPLIT distance="350" swimtime="00:05:28.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="519" swimtime="00:02:39.32" resultid="3403" heatid="4749" lane="3" entrytime="00:02:41.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:02:00.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="418" swimtime="00:05:29.74" resultid="3404" heatid="4797" lane="8" entrytime="00:05:22.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:01:58.00" />
                    <SPLIT distance="200" swimtime="00:02:41.40" />
                    <SPLIT distance="250" swimtime="00:03:23.27" />
                    <SPLIT distance="300" swimtime="00:04:05.65" />
                    <SPLIT distance="350" swimtime="00:04:50.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kośmider" birthdate="1966-03-01" gender="M" nation="POL" license="512914700009" athleteid="3437">
              <RESULTS>
                <RESULT eventid="1090" points="454" swimtime="00:00:31.80" resultid="3438" heatid="4610" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="1182" points="487" swimtime="00:11:26.17" resultid="3439" heatid="4635" lane="6" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:23.30" />
                    <SPLIT distance="150" swimtime="00:02:07.28" />
                    <SPLIT distance="200" swimtime="00:02:51.82" />
                    <SPLIT distance="250" swimtime="00:03:36.23" />
                    <SPLIT distance="300" swimtime="00:04:20.49" />
                    <SPLIT distance="350" swimtime="00:05:04.00" />
                    <SPLIT distance="400" swimtime="00:05:47.18" />
                    <SPLIT distance="450" swimtime="00:06:25.94" />
                    <SPLIT distance="500" swimtime="00:07:11.54" />
                    <SPLIT distance="550" swimtime="00:07:54.07" />
                    <SPLIT distance="600" swimtime="00:08:36.30" />
                    <SPLIT distance="650" swimtime="00:09:18.55" />
                    <SPLIT distance="700" swimtime="00:10:01.95" />
                    <SPLIT distance="750" swimtime="00:10:45.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="457" swimtime="00:03:15.50" resultid="3440" heatid="4657" lane="6" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                    <SPLIT distance="100" swimtime="00:01:33.65" />
                    <SPLIT distance="150" swimtime="00:02:24.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="251" swimtime="00:03:36.79" resultid="3441" heatid="4680" lane="0" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                    <SPLIT distance="100" swimtime="00:01:44.20" />
                    <SPLIT distance="150" swimtime="00:02:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" status="DNS" swimtime="00:00:00.00" resultid="3442" heatid="4722" lane="6" entrytime="00:02:35.00" />
                <RESULT eventid="1597" points="507" swimtime="00:06:12.98" resultid="3443" heatid="4788" lane="5" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                    <SPLIT distance="100" swimtime="00:01:33.09" />
                    <SPLIT distance="150" swimtime="00:02:21.76" />
                    <SPLIT distance="200" swimtime="00:03:09.27" />
                    <SPLIT distance="250" swimtime="00:03:59.66" />
                    <SPLIT distance="300" swimtime="00:04:50.78" />
                    <SPLIT distance="350" swimtime="00:05:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="352" swimtime="00:01:25.72" resultid="3444" heatid="4739" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="536" swimtime="00:05:23.05" resultid="3445" heatid="4797" lane="7" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:17.65" />
                    <SPLIT distance="150" swimtime="00:01:58.98" />
                    <SPLIT distance="200" swimtime="00:02:41.02" />
                    <SPLIT distance="250" swimtime="00:03:22.44" />
                    <SPLIT distance="300" swimtime="00:04:03.84" />
                    <SPLIT distance="350" swimtime="00:04:44.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Matyszewski" birthdate="1971-10-11" gender="M" nation="POL" license="512914700065" athleteid="3468">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="3469" heatid="4608" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="3470" heatid="4625" lane="7" entrytime="00:03:20.00" />
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="3471" heatid="4647" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="3472" heatid="4657" lane="7" entrytime="00:03:20.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="3473" heatid="4691" lane="4" entrytime="00:01:30.00" />
                <RESULT eventid="1524" status="DNS" swimtime="00:00:00.00" resultid="3474" heatid="4718" lane="6" entrytime="00:03:10.00" />
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="3475" heatid="4759" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="3476" heatid="4800" lane="7" entrytime="00:07:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Kaczmarek" birthdate="1985-05-07" gender="F" nation="POL" license="512914600004" athleteid="3341">
              <RESULTS>
                <RESULT eventid="1107" points="580" swimtime="00:02:49.09" resultid="3342" heatid="4621" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:17.64" />
                    <SPLIT distance="150" swimtime="00:02:07.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="589" swimtime="00:00:34.14" resultid="3343" heatid="4643" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1303" points="628" swimtime="00:01:07.81" resultid="3344" heatid="4662" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="544" swimtime="00:01:15.63" resultid="3345" heatid="4708" lane="5" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" status="DNS" swimtime="00:00:00.00" resultid="3346" heatid="4785" lane="0" entrytime="00:08:00.00" />
                <RESULT eventid="1650" status="DNS" swimtime="00:00:00.00" resultid="3347" heatid="4745" lane="3" entrytime="00:02:40.00" />
                <RESULT eventid="1742" status="DNS" swimtime="00:00:00.00" resultid="3348" heatid="4794" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Rudzki" birthdate="1992-06-21" gender="M" nation="POL" athleteid="3429">
              <RESULTS>
                <RESULT eventid="1090" points="599" swimtime="00:00:26.24" resultid="3430" heatid="4614" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1124" points="569" swimtime="00:02:27.40" resultid="3431" heatid="4628" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                    <SPLIT distance="100" swimtime="00:01:05.50" />
                    <SPLIT distance="150" swimtime="00:01:49.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="616" swimtime="00:00:30.52" resultid="3432" heatid="4650" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3433" heatid="4672" lane="8" entrytime="00:01:03.00" />
                <RESULT eventid="1456" points="601" swimtime="00:00:27.56" resultid="3434" heatid="4703" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1633" points="591" swimtime="00:01:03.27" resultid="3435" heatid="4741" lane="7" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="590" swimtime="00:00:33.07" resultid="3436" heatid="4761" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Piaściński" birthdate="1976-09-19" gender="M" nation="POL" license="512914700066" athleteid="3334">
              <RESULTS>
                <RESULT eventid="1124" points="555" swimtime="00:02:38.23" resultid="3335" heatid="4627" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:02:00.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="615" swimtime="00:00:32.47" resultid="3336" heatid="4650" lane="9" entrytime="00:00:33.24" />
                <RESULT eventid="1490" points="660" swimtime="00:01:09.03" resultid="3337" heatid="4712" lane="5" entrytime="00:01:11.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="605" swimtime="00:02:35.50" resultid="3338" heatid="4749" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:15.53" />
                    <SPLIT distance="150" swimtime="00:01:55.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Korc" birthdate="1986-03-27" gender="F" nation="POL" license="512914600038" athleteid="3465">
              <RESULTS>
                <RESULT eventid="1059" points="844" swimtime="00:00:27.49" resultid="3466" heatid="4602" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="1439" points="791" swimtime="00:00:29.69" resultid="3467" heatid="4697" lane="3" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Gajdowska" birthdate="1995-07-17" gender="F" nation="POL" license="512914600068" athleteid="3422">
              <RESULTS>
                <RESULT eventid="1059" points="759" swimtime="00:00:27.86" resultid="3423" heatid="4602" lane="3" entrytime="00:00:27.61" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1303" points="847" swimtime="00:01:00.19" resultid="3424" heatid="4663" lane="4" entrytime="00:00:59.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="642" swimtime="00:00:30.50" resultid="3425" heatid="4697" lane="1" entrytime="00:00:30.03" />
                <RESULT eventid="1507" points="799" swimtime="00:02:14.23" resultid="3426" heatid="4717" lane="5" entrytime="00:02:15.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:04.66" />
                    <SPLIT distance="150" swimtime="00:01:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="566" swimtime="00:00:38.18" resultid="3427" heatid="4755" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1742" points="691" swimtime="00:04:52.43" resultid="3428" heatid="4794" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:06.54" />
                    <SPLIT distance="150" swimtime="00:01:44.50" />
                    <SPLIT distance="200" swimtime="00:02:23.07" />
                    <SPLIT distance="250" swimtime="00:03:01.69" />
                    <SPLIT distance="300" swimtime="00:03:40.53" />
                    <SPLIT distance="350" swimtime="00:04:18.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Dolińska" birthdate="1990-07-06" gender="F" nation="POL" license="512914600056" athleteid="3458">
              <RESULTS>
                <RESULT eventid="1059" points="511" swimtime="00:00:32.18" resultid="3459" heatid="4600" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="1234" points="293" swimtime="00:00:43.01" resultid="3460" heatid="4642" lane="1" entrytime="00:00:39.50" />
                <RESULT eventid="1303" points="428" swimtime="00:01:13.25" resultid="3461" heatid="4662" lane="7" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="300" swimtime="00:01:32.19" resultid="3462" heatid="4707" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="416" swimtime="00:02:43.78" resultid="3463" heatid="4716" lane="3" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="150" swimtime="00:02:01.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" status="DNS" swimtime="00:00:00.00" resultid="3464" heatid="4792" lane="2" entrytime="00:05:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" license="512914700063" athleteid="3497">
              <RESULTS>
                <RESULT eventid="1090" points="264" swimtime="00:00:38.11" resultid="3498" heatid="4606" lane="9" entrytime="00:00:38.78" />
                <RESULT eventid="1286" points="289" swimtime="00:03:47.81" resultid="3499" heatid="4656" lane="0" entrytime="00:03:59.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.40" />
                    <SPLIT distance="100" swimtime="00:01:51.22" />
                    <SPLIT distance="150" swimtime="00:02:51.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3500" heatid="4666" lane="6" entrytime="00:01:32.64" />
                <RESULT eventid="1422" points="291" swimtime="00:01:42.05" resultid="3501" heatid="4691" lane="0" entrytime="00:01:43.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="228" swimtime="00:03:22.90" resultid="3502" heatid="4719" lane="3" entrytime="00:03:33.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                    <SPLIT distance="100" swimtime="00:01:37.80" />
                    <SPLIT distance="150" swimtime="00:02:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="343" swimtime="00:00:42.87" resultid="3503" heatid="4758" lane="7" entrytime="00:00:44.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bożena" lastname="Ayomo" birthdate="1966-02-08" gender="F" nation="POL" license="512914600061" athleteid="3454">
              <RESULTS>
                <RESULT eventid="1059" points="372" swimtime="00:00:39.25" resultid="3455" heatid="4598" lane="0" entrytime="00:00:42.32" />
                <RESULT eventid="1234" points="338" swimtime="00:00:45.91" resultid="3456" heatid="4641" lane="2" entrytime="00:00:46.06" />
                <RESULT eventid="1684" points="324" swimtime="00:00:52.32" resultid="3457" heatid="4752" lane="0" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Lewandowski" birthdate="1986-05-29" gender="M" nation="POL" athleteid="3339">
              <RESULTS>
                <RESULT eventid="1456" points="714" swimtime="00:00:27.00" resultid="3340" heatid="4705" lane="7" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Szyszkowska" birthdate="1996-11-05" gender="F" nation="POL" license="512914600054" athleteid="3377">
              <RESULTS>
                <RESULT eventid="1059" points="703" swimtime="00:00:28.58" resultid="3378" heatid="4602" lane="7" entrytime="00:00:28.50" />
                <RESULT eventid="1107" points="732" swimtime="00:02:36.07" resultid="3379" heatid="4621" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:15.68" />
                    <SPLIT distance="150" swimtime="00:01:59.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="715" swimtime="00:02:52.68" resultid="3380" heatid="4654" lane="4" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:22.97" />
                    <SPLIT distance="150" swimtime="00:02:06.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="755" swimtime="00:01:17.46" resultid="3381" heatid="4688" lane="4" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="717" swimtime="00:00:35.30" resultid="3382" heatid="4755" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Sienicka" birthdate="1990-06-15" gender="F" nation="POL" athleteid="3330">
              <RESULTS>
                <RESULT eventid="1269" points="350" swimtime="00:03:31.22" resultid="3331" heatid="4653" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.86" />
                    <SPLIT distance="100" swimtime="00:01:41.91" />
                    <SPLIT distance="150" swimtime="00:02:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="383" swimtime="00:01:36.45" resultid="3332" heatid="4686" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="404" swimtime="00:00:43.57" resultid="3333" heatid="4752" lane="6" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kulisz" birthdate="1977-06-16" gender="M" nation="POL" license="512914700002" athleteid="3477">
              <RESULTS>
                <RESULT eventid="1090" points="480" swimtime="00:00:30.06" resultid="3478" heatid="4611" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1320" points="466" swimtime="00:01:07.35" resultid="3479" heatid="4671" lane="9" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="437" swimtime="00:00:33.24" resultid="3480" heatid="4699" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1524" status="DNS" swimtime="00:00:00.00" resultid="3481" heatid="4723" lane="1" entrytime="00:02:24.00" />
                <RESULT eventid="1633" points="355" swimtime="00:01:20.22" resultid="3482" heatid="4739" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Uladzislau" lastname="Kunkevich" birthdate="1998-07-15" gender="M" nation="POL" license="512914700069" athleteid="3364">
              <RESULTS>
                <RESULT eventid="1090" points="742" swimtime="00:00:24.63" resultid="3365" heatid="4617" lane="0" entrytime="00:00:24.50" />
                <RESULT eventid="1252" points="769" swimtime="00:00:27.76" resultid="3366" heatid="4651" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1456" status="DNS" swimtime="00:00:00.00" resultid="3367" heatid="4704" lane="2" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Koba-Gołaszewska" birthdate="1986-07-01" gender="F" nation="POL" athleteid="3413">
              <RESULTS>
                <RESULT eventid="1059" points="574" swimtime="00:00:31.26" resultid="3414" heatid="4600" lane="5" entrytime="00:00:31.30" />
                <RESULT eventid="1303" points="543" swimtime="00:01:11.18" resultid="3415" heatid="4662" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="505" swimtime="00:00:34.48" resultid="3416" heatid="4695" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1507" points="379" swimtime="00:02:53.93" resultid="3417" heatid="4716" lane="2" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:23.19" />
                    <SPLIT distance="150" swimtime="00:02:09.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="355" swimtime="00:06:15.86" resultid="3418" heatid="4793" lane="5" entrytime="00:06:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:24.53" />
                    <SPLIT distance="150" swimtime="00:02:12.12" />
                    <SPLIT distance="200" swimtime="00:03:00.48" />
                    <SPLIT distance="250" swimtime="00:03:49.64" />
                    <SPLIT distance="300" swimtime="00:04:40.11" />
                    <SPLIT distance="350" swimtime="00:05:29.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Romuald" lastname="Kozłowski" birthdate="1966-08-13" gender="M" nation="POL" license="512914700012" athleteid="3446">
              <RESULTS>
                <RESULT eventid="1090" points="625" swimtime="00:00:28.59" resultid="3447" heatid="4613" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1286" points="566" swimtime="00:03:02.01" resultid="3448" heatid="4657" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="100" swimtime="00:01:25.30" />
                    <SPLIT distance="150" swimtime="00:02:13.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="572" swimtime="00:01:21.46" resultid="3449" heatid="4693" lane="9" entrytime="00:01:16.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="610" swimtime="00:00:35.38" resultid="3450" heatid="4761" lane="7" entrytime="00:00:34.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Żemier" birthdate="1982-11-09" gender="M" nation="POL" license="512914700051" athleteid="3484">
              <RESULTS>
                <RESULT eventid="1090" points="748" swimtime="00:00:25.55" resultid="3485" heatid="4607" lane="0" entrytime="00:00:35.40" />
                <RESULT eventid="1124" points="743" swimtime="00:02:24.19" resultid="3486" heatid="4623" lane="7" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="100" swimtime="00:01:06.09" />
                    <SPLIT distance="150" swimtime="00:01:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="769" swimtime="00:00:29.60" resultid="3487" heatid="4651" lane="7" entrytime="00:00:28.30" />
                <RESULT eventid="1320" points="719" swimtime="00:00:57.14" resultid="3488" heatid="4674" lane="7" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="695" swimtime="00:00:27.45" resultid="3489" heatid="4698" lane="6" entrytime="00:00:47.20" />
                <RESULT eventid="1490" points="723" swimtime="00:01:05.11" resultid="3490" heatid="4713" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="742" swimtime="00:01:02.03" resultid="3491" heatid="4739" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="678" swimtime="00:02:25.76" resultid="3492" heatid="4750" lane="6" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:49.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Morawski" birthdate="1994-06-29" gender="M" nation="POL" athleteid="3383">
              <RESULTS>
                <RESULT eventid="1252" points="779" swimtime="00:00:27.64" resultid="3384" heatid="4651" lane="8" entrytime="00:00:29.21" />
                <RESULT eventid="1490" points="761" swimtime="00:01:00.33" resultid="3385" heatid="4713" lane="5" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G1 - Pływak nie złamał powierzchni wody głową przed lub na linii 15 m po starcie lub nawrocie." eventid="1667" status="DSQ" swimtime="00:02:20.71" resultid="3386" heatid="4750" lane="4" entrytime="00:02:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:06.42" />
                    <SPLIT distance="150" swimtime="00:01:44.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Matuzewicz" birthdate="1978-05-05" gender="M" nation="POL" license="512914700017" athleteid="3419">
              <RESULTS>
                <RESULT eventid="1320" points="558" swimtime="00:01:03.45" resultid="3420" heatid="4673" lane="9" entrytime="00:01:01.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="523" swimtime="00:02:26.06" resultid="3421" heatid="4722" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:48.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Timea" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" license="512914600062" athleteid="3368">
              <RESULTS>
                <RESULT eventid="1107" points="519" swimtime="00:03:07.84" resultid="3369" heatid="4620" lane="2" entrytime="00:03:03.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:01:34.38" />
                    <SPLIT distance="150" swimtime="00:02:25.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="462" swimtime="00:23:36.94" resultid="3370" heatid="4637" lane="5" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:01:27.61" />
                    <SPLIT distance="150" swimtime="00:02:15.41" />
                    <SPLIT distance="200" swimtime="00:03:03.42" />
                    <SPLIT distance="250" swimtime="00:03:51.24" />
                    <SPLIT distance="300" swimtime="00:04:39.33" />
                    <SPLIT distance="350" swimtime="00:05:27.18" />
                    <SPLIT distance="400" swimtime="00:06:15.03" />
                    <SPLIT distance="450" swimtime="00:07:02.94" />
                    <SPLIT distance="500" swimtime="00:07:50.88" />
                    <SPLIT distance="550" swimtime="00:08:38.29" />
                    <SPLIT distance="600" swimtime="00:09:25.82" />
                    <SPLIT distance="650" swimtime="00:10:13.40" />
                    <SPLIT distance="700" swimtime="00:11:00.72" />
                    <SPLIT distance="750" swimtime="00:11:48.54" />
                    <SPLIT distance="800" swimtime="00:12:36.34" />
                    <SPLIT distance="850" swimtime="00:13:23.95" />
                    <SPLIT distance="900" swimtime="00:14:11.98" />
                    <SPLIT distance="950" swimtime="00:15:00.13" />
                    <SPLIT distance="1000" swimtime="00:15:48.48" />
                    <SPLIT distance="1050" swimtime="00:16:35.15" />
                    <SPLIT distance="1100" swimtime="00:17:22.18" />
                    <SPLIT distance="1150" swimtime="00:18:09.54" />
                    <SPLIT distance="1200" swimtime="00:18:57.15" />
                    <SPLIT distance="1250" swimtime="00:19:44.34" />
                    <SPLIT distance="1300" swimtime="00:20:31.65" />
                    <SPLIT distance="1350" swimtime="00:21:18.44" />
                    <SPLIT distance="1400" swimtime="00:22:05.78" />
                    <SPLIT distance="1450" swimtime="00:22:52.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="571" swimtime="00:03:18.37" resultid="3371" heatid="4654" lane="7" entrytime="00:03:08.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                    <SPLIT distance="100" swimtime="00:01:36.52" />
                    <SPLIT distance="150" swimtime="00:02:27.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="461" swimtime="00:01:18.19" resultid="3372" heatid="4660" lane="5" entrytime="00:01:18.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="565" swimtime="00:01:31.22" resultid="3373" heatid="4688" lane="8" entrytime="00:01:25.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="491" swimtime="00:02:48.72" resultid="3374" heatid="4716" lane="7" entrytime="00:02:44.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:22.09" />
                    <SPLIT distance="150" swimtime="00:02:05.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="651" swimtime="00:00:39.43" resultid="3375" heatid="4755" lane="9" entrytime="00:00:38.71" />
                <RESULT eventid="1742" points="458" swimtime="00:06:03.87" resultid="3376" heatid="4792" lane="3" entrytime="00:05:49.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:24.78" />
                    <SPLIT distance="150" swimtime="00:02:11.72" />
                    <SPLIT distance="200" swimtime="00:02:59.36" />
                    <SPLIT distance="250" swimtime="00:03:46.00" />
                    <SPLIT distance="300" swimtime="00:04:33.28" />
                    <SPLIT distance="350" swimtime="00:05:19.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kaczmarek" birthdate="1977-06-25" gender="M" nation="POL" license="512914700003" athleteid="3349">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1090" points="787" swimtime="00:00:25.50" resultid="3350" heatid="4616" lane="9" entrytime="00:00:25.66" />
                <RESULT eventid="1252" points="971" swimtime="00:00:27.89" resultid="3351" heatid="4651" lane="3" entrytime="00:00:27.82" />
                <RESULT eventid="1456" points="892" swimtime="00:00:26.22" resultid="3352" heatid="4705" lane="6" entrytime="00:00:25.74" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Miński" birthdate="1956-01-14" gender="M" nation="POL" license="512914700021" athleteid="3451">
              <RESULTS>
                <RESULT eventid="1090" points="268" swimtime="00:00:40.65" resultid="3452" heatid="4605" lane="8" entrytime="00:00:46.00" />
                <RESULT eventid="1182" points="251" swimtime="00:15:53.91" resultid="3453" heatid="4633" lane="6" entrytime="00:16:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                    <SPLIT distance="100" swimtime="00:01:44.99" />
                    <SPLIT distance="150" swimtime="00:02:43.69" />
                    <SPLIT distance="200" swimtime="00:03:45.07" />
                    <SPLIT distance="250" swimtime="00:04:45.89" />
                    <SPLIT distance="300" swimtime="00:05:47.27" />
                    <SPLIT distance="350" swimtime="00:06:48.29" />
                    <SPLIT distance="400" swimtime="00:07:50.20" />
                    <SPLIT distance="450" swimtime="00:08:51.93" />
                    <SPLIT distance="500" swimtime="00:09:53.70" />
                    <SPLIT distance="550" swimtime="00:10:54.29" />
                    <SPLIT distance="600" swimtime="00:11:55.53" />
                    <SPLIT distance="650" swimtime="00:12:56.98" />
                    <SPLIT distance="700" swimtime="00:13:59.03" />
                    <SPLIT distance="750" swimtime="00:14:59.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Korpetta" birthdate="1959-12-27" gender="M" nation="POL" license="112914700013" athleteid="3356">
              <RESULTS>
                <RESULT eventid="1124" points="307" swimtime="00:03:30.48" resultid="3357" heatid="4623" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                    <SPLIT distance="100" swimtime="00:01:44.46" />
                    <SPLIT distance="150" swimtime="00:02:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="340" swimtime="00:13:23.87" resultid="3358" heatid="4634" lane="7" entrytime="00:13:13.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                    <SPLIT distance="100" swimtime="00:01:29.24" />
                    <SPLIT distance="150" swimtime="00:02:20.13" />
                    <SPLIT distance="200" swimtime="00:03:11.84" />
                    <SPLIT distance="250" swimtime="00:04:04.11" />
                    <SPLIT distance="300" swimtime="00:04:56.82" />
                    <SPLIT distance="350" swimtime="00:05:49.65" />
                    <SPLIT distance="400" swimtime="00:06:42.04" />
                    <SPLIT distance="450" swimtime="00:07:34.63" />
                    <SPLIT distance="500" swimtime="00:08:26.38" />
                    <SPLIT distance="550" swimtime="00:09:18.26" />
                    <SPLIT distance="600" swimtime="00:10:09.97" />
                    <SPLIT distance="650" swimtime="00:11:00.66" />
                    <SPLIT distance="700" swimtime="00:11:50.96" />
                    <SPLIT distance="750" swimtime="00:12:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="380" swimtime="00:01:19.57" resultid="3359" heatid="4668" lane="8" entrytime="00:01:19.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="332" swimtime="00:01:35.43" resultid="3360" heatid="4711" lane="7" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="373" swimtime="00:02:57.27" resultid="3361" heatid="4721" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:01:26.60" />
                    <SPLIT distance="150" swimtime="00:02:13.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="370" swimtime="00:03:23.41" resultid="3362" heatid="4748" lane="8" entrytime="00:03:26.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.17" />
                    <SPLIT distance="100" swimtime="00:01:39.26" />
                    <SPLIT distance="150" swimtime="00:02:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="367" swimtime="00:06:23.75" resultid="3363" heatid="4799" lane="7" entrytime="00:06:21.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:02:19.77" />
                    <SPLIT distance="200" swimtime="00:03:10.10" />
                    <SPLIT distance="250" swimtime="00:04:00.96" />
                    <SPLIT distance="300" swimtime="00:04:51.36" />
                    <SPLIT distance="350" swimtime="00:05:38.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1395" points="838" swimtime="00:01:47.94" resultid="3515" heatid="4684" lane="4" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                    <SPLIT distance="100" swimtime="00:00:57.87" />
                    <SPLIT distance="150" swimtime="00:01:23.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3353" number="1" />
                    <RELAYPOSITION athleteid="3315" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3383" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="3364" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" status="DNS" swimtime="00:00:00.00" resultid="3525" heatid="4728" lane="2" entrytime="00:01:48.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1395" points="655" swimtime="00:02:01.39" resultid="3516" heatid="4684" lane="7" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                    <SPLIT distance="150" swimtime="00:01:34.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3334" number="1" />
                    <RELAYPOSITION athleteid="3429" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="3387" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3419" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1565" points="789" swimtime="00:01:42.71" resultid="3517" heatid="4728" lane="5" entrytime="00:01:43.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.65" />
                    <SPLIT distance="100" swimtime="00:00:50.12" />
                    <SPLIT distance="150" swimtime="00:01:17.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3484" number="1" />
                    <RELAYPOSITION athleteid="3349" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="3419" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="3339" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="3">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1395" points="767" swimtime="00:02:01.03" resultid="3518" heatid="4684" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                    <SPLIT distance="100" swimtime="00:01:02.84" />
                    <SPLIT distance="150" swimtime="00:01:30.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3349" number="1" />
                    <RELAYPOSITION athleteid="3446" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3484" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="3437" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1565" points="520" swimtime="00:02:02.16" resultid="3519" heatid="4728" lane="9" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:00:58.02" />
                    <SPLIT distance="150" swimtime="00:01:32.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3477" number="1" />
                    <RELAYPOSITION athleteid="3334" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="3356" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="3446" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1395" points="429" swimtime="00:02:26.85" resultid="3520" heatid="4684" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:17.95" />
                    <SPLIT distance="150" swimtime="00:01:51.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3398" number="1" />
                    <RELAYPOSITION athleteid="3497" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="3477" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="3356" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1371" points="828" swimtime="00:02:10.28" resultid="3521" heatid="4682" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:09.00" />
                    <SPLIT distance="150" swimtime="00:01:39.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3341" number="1" />
                    <RELAYPOSITION athleteid="3377" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3422" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="3413" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1541" points="920" swimtime="00:01:52.08" resultid="3522" heatid="4726" lane="5" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="100" swimtime="00:00:56.51" />
                    <SPLIT distance="150" swimtime="00:01:24.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3465" number="1" />
                    <RELAYPOSITION athleteid="3341" number="2" reactiontime="+4" />
                    <RELAYPOSITION athleteid="3377" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="3422" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1371" points="479" swimtime="00:02:39.38" resultid="3523" heatid="4682" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                    <SPLIT distance="100" swimtime="00:01:25.58" />
                    <SPLIT distance="150" swimtime="00:02:04.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3454" number="1" />
                    <RELAYPOSITION athleteid="3368" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="3458" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="3405" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1541" points="480" swimtime="00:02:18.46" resultid="3524" heatid="4726" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="150" swimtime="00:01:47.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3454" number="1" />
                    <RELAYPOSITION athleteid="3330" number="2" reactiontime="+11" />
                    <RELAYPOSITION athleteid="3458" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3413" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1141" points="888" swimtime="00:01:45.26" resultid="3505" heatid="4630" lane="4" entrytime="00:01:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="100" swimtime="00:00:52.54" />
                    <SPLIT distance="150" swimtime="00:01:20.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3377" number="1" />
                    <RELAYPOSITION athleteid="3364" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3422" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3315" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1718" points="759" swimtime="00:02:02.77" resultid="3506" heatid="4765" lane="4" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="100" swimtime="00:00:58.66" />
                    <SPLIT distance="150" swimtime="00:01:29.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3383" number="1" />
                    <RELAYPOSITION athleteid="3315" number="2" reactiontime="+21" />
                    <RELAYPOSITION athleteid="3377" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="3330" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1141" points="589" swimtime="00:01:59.42" resultid="3507" heatid="4630" lane="6" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:06.20" />
                    <SPLIT distance="150" swimtime="00:01:31.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3405" number="1" />
                    <RELAYPOSITION athleteid="3458" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3387" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3429" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1718" points="652" swimtime="00:02:07.70" resultid="3508" heatid="4765" lane="3" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:04.71" />
                    <SPLIT distance="150" swimtime="00:01:39.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3334" number="1" />
                    <RELAYPOSITION athleteid="3429" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3413" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="3422" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="3">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1141" points="900" swimtime="00:01:45.91" resultid="3509" heatid="4630" lane="3" entrytime="00:01:52.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.35" />
                    <SPLIT distance="100" swimtime="00:00:54.48" />
                    <SPLIT distance="150" swimtime="00:01:19.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3349" number="1" />
                    <RELAYPOSITION athleteid="3341" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3484" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3465" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1718" points="689" swimtime="00:02:08.18" resultid="3510" heatid="4765" lane="5" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                    <SPLIT distance="100" swimtime="00:01:06.41" />
                    <SPLIT distance="150" swimtime="00:01:34.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3349" number="1" />
                    <RELAYPOSITION athleteid="3368" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3484" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="3405" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1141" points="598" swimtime="00:02:04.54" resultid="3511" heatid="4630" lane="7" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:05.84" />
                    <SPLIT distance="150" swimtime="00:01:36.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3368" number="1" />
                    <RELAYPOSITION athleteid="3437" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3413" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3446" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1718" status="DNS" swimtime="00:00:00.00" resultid="3512" heatid="4765" lane="7" entrytime="00:02:12.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3454" number="1" />
                    <RELAYPOSITION athleteid="3446" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3437" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3493" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="1141" points="339" swimtime="00:02:26.53" resultid="3513" heatid="4629" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                    <SPLIT distance="100" swimtime="00:01:19.90" />
                    <SPLIT distance="150" swimtime="00:01:57.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3454" number="1" />
                    <RELAYPOSITION athleteid="3321" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3497" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3477" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="1718" status="DNS" swimtime="00:00:00.00" resultid="3514" heatid="4765" lane="9" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3398" number="1" />
                    <RELAYPOSITION athleteid="3497" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3321" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3405" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="11314" nation="POL" region="14" clubid="3581" name="Fundacja HASTEN Warszawa" shortname="HASTEN Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Natalia" lastname="Pawlaczek" birthdate="1993-01-04" gender="F" nation="POL" license="111314600002" athleteid="3582">
              <RESULTS>
                <RESULT eventid="1059" points="773" swimtime="00:00:28.04" resultid="3583" heatid="4602" lane="4" entrytime="00:00:27.27" />
                <RESULT eventid="1439" points="769" swimtime="00:00:29.99" resultid="3584" heatid="4697" lane="4" entrytime="00:00:28.99" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="3779" name="KS WARTA Poznań" shortname="WARTA Poznań">
          <ATHLETES>
            <ATHLETE firstname="Błażej" lastname="Wachowski" birthdate="1980-10-08" gender="M" nation="POL" license="100115700545" athleteid="3808">
              <RESULTS>
                <RESULT eventid="1090" points="528" swimtime="00:00:28.70" resultid="3809" heatid="4612" lane="3" entrytime="00:00:28.90" />
                <RESULT eventid="1182" points="468" swimtime="00:11:04.25" resultid="3810" heatid="4635" lane="4" entrytime="00:10:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:18.50" />
                    <SPLIT distance="150" swimtime="00:02:00.81" />
                    <SPLIT distance="200" swimtime="00:02:43.20" />
                    <SPLIT distance="250" swimtime="00:03:25.46" />
                    <SPLIT distance="300" swimtime="00:04:07.80" />
                    <SPLIT distance="350" swimtime="00:04:50.15" />
                    <SPLIT distance="400" swimtime="00:05:32.84" />
                    <SPLIT distance="450" swimtime="00:06:15.15" />
                    <SPLIT distance="500" swimtime="00:06:57.04" />
                    <SPLIT distance="550" swimtime="00:07:39.00" />
                    <SPLIT distance="600" swimtime="00:08:21.15" />
                    <SPLIT distance="650" swimtime="00:09:03.43" />
                    <SPLIT distance="700" swimtime="00:09:45.27" />
                    <SPLIT distance="750" swimtime="00:10:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="402" swimtime="00:02:49.99" resultid="3811" heatid="4681" lane="0" entrytime="00:02:46.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:18.87" />
                    <SPLIT distance="150" swimtime="00:02:04.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="481" swimtime="00:02:25.01" resultid="3812" heatid="4723" lane="2" entrytime="00:02:22.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:11.40" />
                    <SPLIT distance="150" swimtime="00:01:49.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" status="DNS" swimtime="00:00:00.00" resultid="3813" heatid="4740" lane="2" entrytime="00:01:12.15" />
                <RESULT eventid="1766" points="491" swimtime="00:05:12.74" resultid="3814" heatid="4796" lane="8" entrytime="00:05:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="150" swimtime="00:01:54.73" />
                    <SPLIT distance="200" swimtime="00:02:34.73" />
                    <SPLIT distance="250" swimtime="00:03:14.74" />
                    <SPLIT distance="300" swimtime="00:03:55.01" />
                    <SPLIT distance="350" swimtime="00:04:35.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Kuca" birthdate="1994-07-23" gender="M" nation="POL" license="100115700396" athleteid="3798">
              <RESULTS>
                <RESULT eventid="1090" points="752" swimtime="00:00:24.52" resultid="3799" heatid="4617" lane="2" entrytime="00:00:24.20" />
                <RESULT eventid="1354" points="711" swimtime="00:02:15.24" resultid="3800" heatid="4681" lane="4" entrytime="00:02:15.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                    <SPLIT distance="100" swimtime="00:01:01.76" />
                    <SPLIT distance="150" swimtime="00:01:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="743" swimtime="00:00:58.59" resultid="3801" heatid="4742" lane="5" entrytime="00:00:58.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Zawadka" birthdate="1978-12-30" gender="M" nation="POL" license="500115700748" athleteid="3831">
              <RESULTS>
                <RESULT eventid="1456" points="502" swimtime="00:00:31.74" resultid="3832" heatid="4701" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1633" points="386" swimtime="00:01:18.02" resultid="3991" heatid="4739" lane="4" entrytime="00:01:17.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Wiśniewska" birthdate="1997-10-01" gender="F" nation="POL" license="500115600544" athleteid="3822">
              <RESULTS>
                <RESULT eventid="1107" points="750" swimtime="00:02:34.83" resultid="3823" heatid="4621" lane="4" entrytime="00:02:35.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:13.55" />
                    <SPLIT distance="150" swimtime="00:01:56.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="521" swimtime="00:10:53.18" resultid="3824" heatid="4632" lane="3" entrytime="00:10:26.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:15.66" />
                    <SPLIT distance="150" swimtime="00:01:56.13" />
                    <SPLIT distance="200" swimtime="00:02:36.93" />
                    <SPLIT distance="250" swimtime="00:03:18.38" />
                    <SPLIT distance="300" swimtime="00:03:59.16" />
                    <SPLIT distance="350" swimtime="00:04:40.29" />
                    <SPLIT distance="400" swimtime="00:05:22.00" />
                    <SPLIT distance="450" swimtime="00:06:03.22" />
                    <SPLIT distance="500" swimtime="00:06:44.96" />
                    <SPLIT distance="550" swimtime="00:07:26.32" />
                    <SPLIT distance="600" swimtime="00:08:08.27" />
                    <SPLIT distance="650" swimtime="00:08:49.76" />
                    <SPLIT distance="700" swimtime="00:09:31.74" />
                    <SPLIT distance="750" swimtime="00:10:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="834" swimtime="00:02:44.05" resultid="3825" heatid="4654" lane="5" entrytime="00:02:49.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="150" swimtime="00:02:01.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="603" swimtime="00:01:07.39" resultid="3826" heatid="4663" lane="9" entrytime="00:01:07.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1404" points="838" swimtime="00:01:14.82" resultid="3827" heatid="4688" lane="5" entrytime="00:01:17.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="737" swimtime="00:05:35.18" resultid="3828" heatid="4785" lane="4" entrytime="00:05:34.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:14.16" />
                    <SPLIT distance="150" swimtime="00:02:00.38" />
                    <SPLIT distance="200" swimtime="00:02:43.66" />
                    <SPLIT distance="250" swimtime="00:03:27.91" />
                    <SPLIT distance="300" swimtime="00:04:13.43" />
                    <SPLIT distance="350" swimtime="00:04:55.11" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1684" points="761" swimtime="00:00:34.61" resultid="3829" heatid="4755" lane="3" entrytime="00:00:35.68" />
                <RESULT eventid="1742" points="558" swimtime="00:05:14.01" resultid="3830" heatid="4791" lane="6" entrytime="00:05:06.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:54.58" />
                    <SPLIT distance="200" swimtime="00:02:34.88" />
                    <SPLIT distance="250" swimtime="00:03:14.85" />
                    <SPLIT distance="300" swimtime="00:03:55.18" />
                    <SPLIT distance="350" swimtime="00:04:35.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Skurczyńska" birthdate="1971-10-13" gender="F" nation="POL" license="500115600746" athleteid="3780">
              <RESULTS>
                <RESULT eventid="1059" points="296" swimtime="00:00:40.63" resultid="3781" heatid="4597" lane="4" entrytime="00:00:43.53" />
                <RESULT eventid="1269" points="286" swimtime="00:04:09.87" resultid="3782" heatid="4653" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.33" />
                    <SPLIT distance="100" swimtime="00:01:55.77" />
                    <SPLIT distance="150" swimtime="00:03:04.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="331" swimtime="00:01:48.97" resultid="3783" heatid="4686" lane="6" entrytime="00:01:54.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="350" swimtime="00:00:48.49" resultid="3784" heatid="4752" lane="5" entrytime="00:00:52.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Majchrzak" birthdate="1983-01-21" gender="M" nation="POL" license="100115700630" athleteid="3802">
              <RESULTS>
                <RESULT eventid="1090" points="584" swimtime="00:00:27.75" resultid="3803" heatid="4615" lane="2" entrytime="00:00:26.40" />
                <RESULT eventid="1320" points="593" swimtime="00:01:00.93" resultid="3804" heatid="4673" lane="5" entrytime="00:00:59.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="554" swimtime="00:00:29.60" resultid="3805" heatid="4704" lane="0" entrytime="00:00:28.40" />
                <RESULT eventid="1633" points="555" swimtime="00:01:08.34" resultid="3806" heatid="4741" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="3807" heatid="4802" lane="8" />
                <RESULT eventid="1524" points="550" swimtime="00:02:18.63" resultid="3990" heatid="4724" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="150" swimtime="00:01:44.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Krupińska" birthdate="1953-05-24" gender="F" nation="POL" license="500115600520" athleteid="3785">
              <RESULTS>
                <RESULT eventid="1059" points="227" swimtime="00:00:50.36" resultid="3786" heatid="4596" lane="4" entrytime="00:00:58.00" />
                <RESULT eventid="1303" points="167" swimtime="00:02:01.34" resultid="3787" heatid="4659" lane="2" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="474" swimtime="00:02:02.96" resultid="3788" heatid="4686" lane="1" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="180" swimtime="00:04:25.10" resultid="3789" heatid="4714" lane="4" entrytime="00:04:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.89" />
                    <SPLIT distance="100" swimtime="00:02:09.33" />
                    <SPLIT distance="150" swimtime="00:03:20.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="408" swimtime="00:00:56.17" resultid="3790" heatid="4752" lane="3" entrytime="00:00:54.50" />
                <RESULT eventid="1269" points="460" swimtime="00:04:30.90" resultid="3989" heatid="4652" lane="3" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.65" />
                    <SPLIT distance="100" swimtime="00:02:13.34" />
                    <SPLIT distance="150" swimtime="00:03:25.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Janyga" birthdate="1966-03-27" gender="M" nation="POL" license="100115700346" athleteid="3791">
              <RESULTS>
                <RESULT eventid="1090" points="596" swimtime="00:00:29.04" resultid="3792" heatid="4611" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1252" points="672" swimtime="00:00:33.14" resultid="3793" heatid="4649" lane="2" entrytime="00:00:34.50" />
                <RESULT eventid="1490" points="668" swimtime="00:01:12.62" resultid="3794" heatid="4712" lane="6" entrytime="00:01:13.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="583" swimtime="00:02:28.44" resultid="3795" heatid="4723" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                    <SPLIT distance="150" swimtime="00:01:51.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="604" swimtime="00:02:46.55" resultid="3796" heatid="4749" lane="7" entrytime="00:02:45.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:21.53" />
                    <SPLIT distance="150" swimtime="00:02:05.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Witt" birthdate="1991-08-11" gender="M" nation="POL" license="500115700645" athleteid="3815">
              <RESULTS>
                <RESULT eventid="1090" points="705" swimtime="00:00:24.86" resultid="3816" heatid="4616" lane="4" entrytime="00:00:24.82" />
                <RESULT eventid="1320" points="698" swimtime="00:00:56.12" resultid="3817" heatid="4675" lane="8" entrytime="00:00:55.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="655" swimtime="00:00:26.78" resultid="3818" heatid="4704" lane="4" entrytime="00:00:26.69" />
                <RESULT eventid="1524" points="603" swimtime="00:02:09.62" resultid="3819" heatid="4725" lane="9" entrytime="00:02:10.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                    <SPLIT distance="100" swimtime="00:01:02.14" />
                    <SPLIT distance="150" swimtime="00:01:36.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="575" swimtime="00:01:03.84" resultid="3820" heatid="4741" lane="4" entrytime="00:01:04.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="568" swimtime="00:04:47.52" resultid="3821" heatid="4796" lane="4" entrytime="00:04:47.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:05.79" />
                    <SPLIT distance="150" swimtime="00:01:42.48" />
                    <SPLIT distance="200" swimtime="00:02:19.49" />
                    <SPLIT distance="250" swimtime="00:02:56.96" />
                    <SPLIT distance="300" swimtime="00:03:35.11" />
                    <SPLIT distance="350" swimtime="00:04:12.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="579" swimtime="00:02:06.51" resultid="3833" heatid="4684" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:37.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3791" number="1" />
                    <RELAYPOSITION athleteid="3802" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3815" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="3808" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="643" swimtime="00:01:49.96" resultid="3834" heatid="4728" lane="6" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.17" />
                    <SPLIT distance="100" swimtime="00:00:52.95" />
                    <SPLIT distance="150" swimtime="00:01:21.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3815" number="1" />
                    <RELAYPOSITION athleteid="3808" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="3791" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3802" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="11614" nation="POL" region="14" clubid="2686" name="5STYL Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Łatkowska" birthdate="1965-06-10" gender="F" nation="POL" athleteid="2745">
              <RESULTS>
                <RESULT eventid="1107" points="246" swimtime="00:04:01.76" resultid="2746" heatid="4619" lane="8" entrytime="00:03:58.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.64" />
                    <SPLIT distance="100" swimtime="00:01:57.11" />
                    <SPLIT distance="150" swimtime="00:03:05.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="242" swimtime="00:29:48.89" resultid="2747" heatid="4637" lane="6" entrytime="00:28:48.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                    <SPLIT distance="100" swimtime="00:01:44.75" />
                    <SPLIT distance="150" swimtime="00:02:41.51" />
                    <SPLIT distance="200" swimtime="00:03:40.53" />
                    <SPLIT distance="250" swimtime="00:04:38.73" />
                    <SPLIT distance="300" swimtime="00:05:39.10" />
                    <SPLIT distance="350" swimtime="00:06:36.04" />
                    <SPLIT distance="400" swimtime="00:07:37.25" />
                    <SPLIT distance="450" swimtime="00:08:36.55" />
                    <SPLIT distance="500" swimtime="00:09:37.20" />
                    <SPLIT distance="550" swimtime="00:10:35.25" />
                    <SPLIT distance="600" swimtime="00:11:35.83" />
                    <SPLIT distance="650" swimtime="00:12:33.60" />
                    <SPLIT distance="700" swimtime="00:13:35.24" />
                    <SPLIT distance="750" swimtime="00:14:35.19" />
                    <SPLIT distance="800" swimtime="00:15:37.58" />
                    <SPLIT distance="850" swimtime="00:16:38.90" />
                    <SPLIT distance="900" swimtime="00:17:41.09" />
                    <SPLIT distance="950" swimtime="00:18:41.54" />
                    <SPLIT distance="1000" swimtime="00:19:42.99" />
                    <SPLIT distance="1050" swimtime="00:20:44.57" />
                    <SPLIT distance="1100" swimtime="00:21:45.66" />
                    <SPLIT distance="1150" swimtime="00:22:45.68" />
                    <SPLIT distance="1200" swimtime="00:23:47.48" />
                    <SPLIT distance="1250" swimtime="00:24:47.56" />
                    <SPLIT distance="1300" swimtime="00:25:50.19" />
                    <SPLIT distance="1350" swimtime="00:26:49.19" />
                    <SPLIT distance="1400" swimtime="00:27:51.01" />
                    <SPLIT distance="1450" swimtime="00:28:49.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="230" swimtime="00:00:52.21" resultid="2748" heatid="4641" lane="0" entrytime="00:00:52.68" entrycourse="LCM" />
                <RESULT eventid="1303" points="257" swimtime="00:01:37.51" resultid="2749" heatid="4660" lane="9" entrytime="00:01:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="174" swimtime="00:00:54.61" resultid="2750" heatid="4694" lane="5" entrytime="00:00:54.90" entrycourse="LCM" />
                <RESULT eventid="1507" points="247" swimtime="00:03:37.04" resultid="2751" heatid="4715" lane="8" entrytime="00:03:28.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.39" />
                    <SPLIT distance="100" swimtime="00:01:45.54" />
                    <SPLIT distance="150" swimtime="00:02:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="257" swimtime="00:00:56.46" resultid="2752" heatid="4752" lane="1" entrytime="00:00:55.60" entrycourse="LCM" />
                <RESULT eventid="1742" points="240" swimtime="00:07:35.52" resultid="2753" heatid="4793" lane="9" entrytime="00:07:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="100" swimtime="00:01:45.67" />
                    <SPLIT distance="150" swimtime="00:02:42.52" />
                    <SPLIT distance="200" swimtime="00:03:42.03" />
                    <SPLIT distance="250" swimtime="00:04:39.95" />
                    <SPLIT distance="300" swimtime="00:05:41.52" />
                    <SPLIT distance="350" swimtime="00:06:40.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Broniszewski" birthdate="1980-09-26" gender="M" nation="POL" athleteid="2693">
              <RESULTS>
                <RESULT eventid="1090" points="351" swimtime="00:00:32.88" resultid="2694" heatid="4608" lane="7" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1320" points="318" swimtime="00:01:14.96" resultid="2695" heatid="4668" lane="1" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="362" swimtime="00:01:29.17" resultid="2696" heatid="4691" lane="3" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="314" swimtime="00:02:47.09" resultid="2697" heatid="4721" lane="7" entrytime="00:02:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:02:02.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="372" swimtime="00:00:40.09" resultid="2698" heatid="4758" lane="4" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1766" points="320" swimtime="00:06:00.47" resultid="2699" heatid="4799" lane="6" entrytime="00:06:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:10.45" />
                    <SPLIT distance="200" swimtime="00:02:56.84" />
                    <SPLIT distance="250" swimtime="00:03:42.34" />
                    <SPLIT distance="300" swimtime="00:04:28.85" />
                    <SPLIT distance="350" swimtime="00:05:14.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Barnasiuk" birthdate="1992-02-04" gender="M" nation="POL" athleteid="2711">
              <RESULTS>
                <RESULT eventid="1124" points="645" swimtime="00:02:21.38" resultid="2712" heatid="4628" lane="3" entrytime="00:02:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="100" swimtime="00:01:06.75" />
                    <SPLIT distance="150" swimtime="00:01:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="691" swimtime="00:02:36.10" resultid="2713" heatid="4658" lane="2" entrytime="00:02:37.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:01:56.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="631" swimtime="00:01:11.40" resultid="2714" heatid="4693" lane="1" entrytime="00:01:11.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="587" swimtime="00:05:11.33" resultid="2715" heatid="4787" lane="3" entrytime="00:05:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                    <SPLIT distance="100" swimtime="00:01:08.32" />
                    <SPLIT distance="150" swimtime="00:01:52.35" />
                    <SPLIT distance="200" swimtime="00:02:35.64" />
                    <SPLIT distance="250" swimtime="00:03:18.50" />
                    <SPLIT distance="300" swimtime="00:04:01.65" />
                    <SPLIT distance="350" swimtime="00:04:37.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="576" swimtime="00:01:03.80" resultid="2716" heatid="4741" lane="6" entrytime="00:01:05.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="628" swimtime="00:00:32.39" resultid="2717" heatid="4762" lane="9" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Niedźwiadek" birthdate="1993-10-18" gender="M" nation="POL" athleteid="2687">
              <RESULTS>
                <RESULT eventid="1090" points="425" swimtime="00:00:29.42" resultid="2688" heatid="4612" lane="7" entrytime="00:00:29.37" entrycourse="LCM" />
                <RESULT eventid="1182" points="459" swimtime="00:10:33.20" resultid="2689" heatid="4636" lane="9" entrytime="00:10:41.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:50.04" />
                    <SPLIT distance="200" swimtime="00:02:29.07" />
                    <SPLIT distance="250" swimtime="00:03:08.35" />
                    <SPLIT distance="300" swimtime="00:03:48.15" />
                    <SPLIT distance="350" swimtime="00:04:28.03" />
                    <SPLIT distance="400" swimtime="00:05:07.89" />
                    <SPLIT distance="450" swimtime="00:05:48.15" />
                    <SPLIT distance="500" swimtime="00:06:29.19" />
                    <SPLIT distance="550" swimtime="00:07:09.93" />
                    <SPLIT distance="600" swimtime="00:07:50.81" />
                    <SPLIT distance="650" swimtime="00:08:32.06" />
                    <SPLIT distance="700" swimtime="00:09:13.65" />
                    <SPLIT distance="750" swimtime="00:09:55.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="458" swimtime="00:01:04.56" resultid="2690" heatid="4671" lane="3" entrytime="00:01:05.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="462" swimtime="00:02:21.66" resultid="2691" heatid="4723" lane="7" entrytime="00:02:22.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:09.10" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="508" swimtime="00:04:58.27" resultid="2692" heatid="4796" lane="6" entrytime="00:04:57.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:11.63" />
                    <SPLIT distance="150" swimtime="00:01:49.21" />
                    <SPLIT distance="200" swimtime="00:02:27.24" />
                    <SPLIT distance="250" swimtime="00:03:05.39" />
                    <SPLIT distance="300" swimtime="00:03:44.07" />
                    <SPLIT distance="350" swimtime="00:04:21.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Butscher" birthdate="1975-01-18" gender="M" nation="POL" athleteid="2760">
              <RESULTS>
                <RESULT eventid="1090" points="345" swimtime="00:00:33.57" resultid="2761" heatid="4609" lane="1" entrytime="00:00:32.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Korzeniowski" birthdate="1985-07-09" gender="M" nation="POL" athleteid="2726">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1090" points="918" swimtime="00:00:23.41" resultid="2727" heatid="4617" lane="4" entrytime="00:00:23.80" entrycourse="LCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1124" points="917" swimtime="00:02:09.30" resultid="2728" heatid="4628" lane="4" entrytime="00:02:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                    <SPLIT distance="100" swimtime="00:01:00.48" />
                    <SPLIT distance="150" swimtime="00:01:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="837" swimtime="00:00:53.88" resultid="2729" heatid="4675" lane="4" entrytime="00:00:52.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="943" swimtime="00:00:24.61" resultid="2730" heatid="4705" lane="5" entrytime="00:00:24.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Krawczyk" birthdate="1978-09-10" gender="M" nation="POL" athleteid="2737">
              <RESULTS>
                <RESULT eventid="1090" points="390" swimtime="00:00:32.21" resultid="2738" heatid="4609" lane="0" entrytime="00:00:32.50" entrycourse="LCM" />
                <RESULT eventid="1182" points="318" swimtime="00:12:42.48" resultid="2739" heatid="4634" lane="5" entrytime="00:12:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="100" swimtime="00:01:24.68" />
                    <SPLIT distance="200" swimtime="00:03:01.53" />
                    <SPLIT distance="250" swimtime="00:03:50.47" />
                    <SPLIT distance="300" swimtime="00:04:39.97" />
                    <SPLIT distance="350" swimtime="00:05:28.47" />
                    <SPLIT distance="400" swimtime="00:06:18.05" />
                    <SPLIT distance="450" swimtime="00:07:06.76" />
                    <SPLIT distance="500" swimtime="00:07:55.40" />
                    <SPLIT distance="550" swimtime="00:08:43.84" />
                    <SPLIT distance="600" swimtime="00:09:32.62" />
                    <SPLIT distance="650" swimtime="00:10:22.33" />
                    <SPLIT distance="700" swimtime="00:11:09.37" />
                    <SPLIT distance="750" swimtime="00:11:56.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="377" swimtime="00:01:12.29" resultid="2740" heatid="4668" lane="5" entrytime="00:01:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="344" swimtime="00:05:58.18" resultid="2741" heatid="4799" lane="2" entrytime="00:06:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:19.37" />
                    <SPLIT distance="150" swimtime="00:02:04.77" />
                    <SPLIT distance="200" swimtime="00:02:51.85" />
                    <SPLIT distance="250" swimtime="00:03:39.18" />
                    <SPLIT distance="300" swimtime="00:04:26.90" />
                    <SPLIT distance="350" swimtime="00:05:14.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Dubiel" birthdate="1993-12-12" gender="M" nation="POL" athleteid="2718">
              <RESULTS>
                <RESULT eventid="1320" points="830" swimtime="00:00:52.99" resultid="2719" heatid="4675" lane="3" entrytime="00:00:54.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.60" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1524" points="836" swimtime="00:01:56.28" resultid="2720" heatid="4725" lane="5" entrytime="00:01:56.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                    <SPLIT distance="100" swimtime="00:00:57.49" />
                    <SPLIT distance="150" swimtime="00:01:27.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Wziątek" birthdate="1988-01-14" gender="M" nation="POL" athleteid="2703">
              <RESULTS>
                <RESULT eventid="1320" points="410" swimtime="00:01:08.34" resultid="2704" heatid="4670" lane="5" entrytime="00:01:09.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="366" swimtime="00:02:37.64" resultid="2705" heatid="4722" lane="2" entrytime="00:02:35.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                    <SPLIT distance="150" swimtime="00:01:55.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="314" swimtime="00:01:18.86" resultid="2706" heatid="4739" lane="5" entrytime="00:01:18.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="363" swimtime="00:05:44.63" resultid="2707" heatid="4798" lane="5" entrytime="00:05:34.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="100" swimtime="00:01:16.25" />
                    <SPLIT distance="150" swimtime="00:01:59.59" />
                    <SPLIT distance="200" swimtime="00:02:44.04" />
                    <SPLIT distance="250" swimtime="00:03:30.18" />
                    <SPLIT distance="300" swimtime="00:04:16.79" />
                    <SPLIT distance="350" swimtime="00:05:02.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Cieślak" birthdate="1992-01-07" gender="M" nation="POL" athleteid="2708">
              <RESULTS>
                <RESULT eventid="1090" points="794" swimtime="00:00:23.89" resultid="2709" heatid="4617" lane="3" entrytime="00:00:24.00" entrycourse="LCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1456" points="818" swimtime="00:00:24.87" resultid="2710" heatid="4705" lane="4" entrytime="00:00:24.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Wiśniewski" birthdate="1977-02-19" gender="M" nation="POL" athleteid="2762">
              <RESULTS>
                <RESULT eventid="1090" points="349" swimtime="00:00:33.42" resultid="2763" heatid="4608" lane="3" entrytime="00:00:33.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Kozyra" birthdate="1959-12-25" gender="M" nation="POL" athleteid="2731">
              <RESULTS>
                <RESULT eventid="1090" points="346" swimtime="00:00:35.93" resultid="2732" heatid="4607" lane="7" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1124" points="267" swimtime="00:03:40.36" resultid="2733" heatid="4624" lane="8" entrytime="00:03:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                    <SPLIT distance="100" swimtime="00:01:42.90" />
                    <SPLIT distance="150" swimtime="00:02:52.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="350" swimtime="00:01:21.81" resultid="2734" heatid="4666" lane="4" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="262" swimtime="00:00:43.18" resultid="2735" heatid="4698" lane="4" entrytime="00:00:42.00" entrycourse="LCM" />
                <RESULT eventid="1524" points="301" swimtime="00:03:10.50" resultid="2736" heatid="4720" lane="0" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:01:27.22" />
                    <SPLIT distance="150" swimtime="00:02:19.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Dzikiewicz" birthdate="1990-10-27" gender="M" nation="POL" athleteid="2754">
              <RESULTS>
                <RESULT eventid="1090" points="296" swimtime="00:00:33.19" resultid="2755" heatid="4608" lane="0" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1320" points="230" swimtime="00:01:21.25" resultid="2756" heatid="4667" lane="0" entrytime="00:01:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Budzis" birthdate="1990-03-04" gender="F" nation="POL" athleteid="2766">
              <RESULTS>
                <RESULT eventid="1059" points="639" swimtime="00:00:29.88" resultid="2767" heatid="4602" lane="9" entrytime="00:00:29.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Serafin" birthdate="1979-03-06" gender="M" nation="POL" athleteid="2764">
              <RESULTS>
                <RESULT eventid="1090" points="296" swimtime="00:00:34.80" resultid="2765" heatid="4606" lane="7" entrytime="00:00:38.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Pilarska" birthdate="1997-02-16" gender="F" nation="POL" athleteid="2742">
              <RESULTS>
                <RESULT eventid="1059" points="696" swimtime="00:00:28.68" resultid="2743" heatid="4601" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1439" points="630" swimtime="00:00:30.69" resultid="2744" heatid="4697" lane="7" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Dubiel" birthdate="1987-01-15" gender="M" nation="POL" athleteid="2721">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1090" points="792" swimtime="00:00:24.59" resultid="2722" heatid="4616" lane="2" entrytime="00:00:25.50" entrycourse="LCM" />
                <RESULT eventid="1252" points="807" swimtime="00:00:28.11" resultid="2723" heatid="4651" lane="1" entrytime="00:00:28.50" entrycourse="LCM" />
                <RESULT eventid="1320" points="734" swimtime="00:00:56.28" resultid="2724" heatid="4675" lane="9" entrytime="00:00:56.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G1 - Pływak nie złamał powierzchni wody głową przed lub na linii 15 m po starcie lub nawrocie." eventid="1490" status="DSQ" swimtime="00:01:02.46" resultid="2725" heatid="4713" lane="3" entrytime="00:01:02.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Kamiński" birthdate="1986-02-11" gender="M" nation="POL" athleteid="2700">
              <RESULTS>
                <RESULT eventid="1090" points="316" swimtime="00:00:33.41" resultid="2701" heatid="4607" lane="6" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1320" points="254" swimtime="00:01:20.16" resultid="2702" heatid="4668" lane="9" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Kulik" birthdate="1981-04-10" gender="M" nation="POL" athleteid="2757">
              <RESULTS>
                <RESULT eventid="1090" points="402" swimtime="00:00:31.42" resultid="2758" heatid="4609" lane="3" entrytime="00:00:31.89" entrycourse="LCM" />
                <RESULT eventid="1320" points="337" swimtime="00:01:13.54" resultid="2759" heatid="4670" lane="0" entrytime="00:01:11.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1395" points="872" swimtime="00:01:47.07" resultid="4410" heatid="4683" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                    <SPLIT distance="100" swimtime="00:00:58.65" />
                    <SPLIT distance="150" swimtime="00:01:23.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2721" number="1" />
                    <RELAYPOSITION athleteid="2708" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="2726" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="2718" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1565" points="891" swimtime="00:01:36.46" resultid="4411" heatid="4727" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.71" />
                    <SPLIT distance="100" swimtime="00:00:47.55" />
                    <SPLIT distance="150" swimtime="00:01:12.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2726" number="1" />
                    <RELAYPOSITION athleteid="2708" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2718" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2721" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1565" points="488" swimtime="00:01:57.90" resultid="4412" heatid="4727" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.35" />
                    <SPLIT distance="100" swimtime="00:00:58.04" />
                    <SPLIT distance="150" swimtime="00:01:27.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2711" number="1" />
                    <RELAYPOSITION athleteid="2693" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="2687" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="2703" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1141" points="835" swimtime="00:01:46.32" resultid="4409" heatid="4629" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.14" />
                    <SPLIT distance="100" swimtime="00:00:48.21" />
                    <SPLIT distance="150" swimtime="00:01:17.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2708" number="1" />
                    <RELAYPOSITION athleteid="2726" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2766" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2742" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="01" clubid="1910" name="UKS ENERGETYK Zgorzelec" shortname="ENERGETYK Zgorzelec">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Daszyński" birthdate="1948-11-29" gender="M" nation="POL" athleteid="1911">
              <RESULTS>
                <RESULT eventid="1124" points="239" swimtime="00:04:45.99" resultid="1912" heatid="4623" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.71" />
                    <SPLIT distance="100" swimtime="00:02:21.26" />
                    <SPLIT distance="150" swimtime="00:03:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="225" swimtime="00:18:16.83" resultid="1913" heatid="4633" lane="2" entrytime="00:17:26.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.46" />
                    <SPLIT distance="100" swimtime="00:02:09.96" />
                    <SPLIT distance="150" swimtime="00:03:20.63" />
                    <SPLIT distance="200" swimtime="00:04:31.10" />
                    <SPLIT distance="250" swimtime="00:05:41.77" />
                    <SPLIT distance="300" swimtime="00:06:52.58" />
                    <SPLIT distance="350" swimtime="00:08:01.53" />
                    <SPLIT distance="400" swimtime="00:09:10.98" />
                    <SPLIT distance="450" swimtime="00:10:19.58" />
                    <SPLIT distance="500" swimtime="00:11:29.19" />
                    <SPLIT distance="550" swimtime="00:12:39.86" />
                    <SPLIT distance="600" swimtime="00:13:49.19" />
                    <SPLIT distance="650" swimtime="00:14:59.16" />
                    <SPLIT distance="700" swimtime="00:16:10.11" />
                    <SPLIT distance="750" swimtime="00:17:13.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="244" swimtime="00:00:55.11" resultid="1914" heatid="4646" lane="8" entrytime="00:00:56.00" />
                <RESULT eventid="1354" points="158" swimtime="00:05:53.64" resultid="1915" heatid="4679" lane="8" entrytime="00:05:32.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.06" />
                    <SPLIT distance="100" swimtime="00:02:42.04" />
                    <SPLIT distance="150" swimtime="00:04:15.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="254" swimtime="00:02:01.83" resultid="1916" heatid="4709" lane="4" entrytime="00:02:01.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="259" swimtime="00:10:19.48" resultid="1917" heatid="4789" lane="8" entrytime="00:09:48.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.59" />
                    <SPLIT distance="100" swimtime="00:02:45.86" />
                    <SPLIT distance="150" swimtime="00:04:03.31" />
                    <SPLIT distance="200" swimtime="00:05:17.70" />
                    <SPLIT distance="250" swimtime="00:06:46.39" />
                    <SPLIT distance="300" swimtime="00:08:12.10" />
                    <SPLIT distance="350" swimtime="00:09:16.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="131" swimtime="00:02:38.67" resultid="1918" heatid="4738" lane="0" entrytime="00:02:32.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="1919" heatid="4801" lane="8" entrytime="00:08:22.58" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03706" nation="POL" region="06" clubid="3883" name="St. SIEMACHA Kraków">
          <ATHLETES>
            <ATHLETE firstname="Paulina" lastname="Palmowska-Latuszek" birthdate="1985-08-01" gender="F" nation="POL" license="503706600141" athleteid="2629">
              <RESULTS>
                <RESULT eventid="1059" points="598" swimtime="00:00:30.83" resultid="2630" heatid="4601" lane="8" entrytime="00:00:30.62" />
                <RESULT eventid="1234" points="559" swimtime="00:00:34.75" resultid="2631" heatid="4643" lane="7" entrytime="00:00:34.80" />
                <RESULT eventid="1303" points="624" swimtime="00:01:07.97" resultid="2632" heatid="4662" lane="5" entrytime="00:01:08.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="564" swimtime="00:01:14.73" resultid="2633" heatid="4708" lane="7" entrytime="00:01:15.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="523" swimtime="00:02:36.32" resultid="2634" heatid="4717" lane="9" entrytime="00:02:36.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="100" swimtime="00:01:14.46" />
                    <SPLIT distance="150" swimtime="00:01:55.49" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1650" points="590" swimtime="00:02:44.73" resultid="2635" heatid="4745" lane="2" entrytime="00:02:44.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:20.56" />
                    <SPLIT distance="150" swimtime="00:02:03.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="484" swimtime="00:05:38.95" resultid="2636" heatid="4792" lane="5" entrytime="00:05:41.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:18.73" />
                    <SPLIT distance="150" swimtime="00:02:02.85" />
                    <SPLIT distance="200" swimtime="00:02:46.17" />
                    <SPLIT distance="250" swimtime="00:03:29.88" />
                    <SPLIT distance="300" swimtime="00:04:14.27" />
                    <SPLIT distance="350" swimtime="00:04:58.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="3835" name="KU AZS UAM Poznań" shortname="AZS UAM Poznań">
          <ATHLETES>
            <ATHLETE firstname="Bartosz" lastname="Kaczmarek" birthdate="1983-07-27" gender="M" nation="POL" license="503315700216" athleteid="3836">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1090" status="DSQ" swimtime="00:00:00.00" resultid="3837" heatid="4604" lane="0" />
                <RESULT eventid="1252" points="482" swimtime="00:00:34.60" resultid="3838" heatid="4645" lane="1" />
                <RESULT eventid="1320" points="489" swimtime="00:01:04.98" resultid="3839" heatid="4664" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="410" swimtime="00:01:18.65" resultid="3840" heatid="4709" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="385" swimtime="00:02:36.21" resultid="3841" heatid="4718" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:14.03" />
                    <SPLIT distance="150" swimtime="00:01:55.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00201" nation="POL" region="01" clubid="3737" name="KS AZS AWF Wrocław" shortname="AZS AWF Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Rytter" birthdate="2001-10-17" gender="M" nation="POL" license="100201700226" athleteid="3745">
              <RESULTS>
                <RESULT eventid="1090" swimtime="00:00:25.38" resultid="3746" heatid="4604" lane="2" />
                <RESULT eventid="1320" swimtime="00:00:55.83" resultid="3747" heatid="4664" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" status="DNS" swimtime="00:00:00.00" resultid="3748" heatid="4756" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Sasin" birthdate="1994-05-29" gender="F" nation="POL" license="100201600097" athleteid="3738">
              <RESULTS>
                <RESULT eventid="1059" points="741" swimtime="00:00:28.09" resultid="3739" heatid="4602" lane="6" entrytime="00:00:27.88" />
                <RESULT eventid="1107" points="791" swimtime="00:02:32.14" resultid="3740" heatid="4621" lane="5" entrytime="00:02:36.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:57.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="789" swimtime="00:01:01.63" resultid="3741" heatid="4663" lane="5" entrytime="00:01:00.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="671" swimtime="00:00:30.06" resultid="3742" heatid="4697" lane="5" entrytime="00:00:29.08" />
                <RESULT eventid="1507" points="717" swimtime="00:02:19.11" resultid="3743" heatid="4717" lane="4" entrytime="00:02:14.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:06.44" />
                    <SPLIT distance="150" swimtime="00:01:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1615" points="716" swimtime="00:01:07.03" resultid="3744" heatid="4736" lane="4" entrytime="00:01:05.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02611" nation="POL" region="11" clubid="1880" name="WETERAN Zabrze">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Twardysko" birthdate="1956-01-16" gender="M" nation="POL" license="102611700035" athleteid="1881">
              <RESULTS>
                <RESULT eventid="1090" points="397" swimtime="00:00:35.66" resultid="1882" heatid="4607" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1182" points="413" swimtime="00:13:28.16" resultid="1883" heatid="4634" lane="2" entrytime="00:13:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:28.75" />
                    <SPLIT distance="150" swimtime="00:02:17.48" />
                    <SPLIT distance="200" swimtime="00:03:08.15" />
                    <SPLIT distance="250" swimtime="00:03:59.25" />
                    <SPLIT distance="300" swimtime="00:04:50.78" />
                    <SPLIT distance="350" swimtime="00:05:42.50" />
                    <SPLIT distance="400" swimtime="00:06:34.15" />
                    <SPLIT distance="450" swimtime="00:07:26.68" />
                    <SPLIT distance="500" swimtime="00:08:18.27" />
                    <SPLIT distance="550" swimtime="00:09:10.87" />
                    <SPLIT distance="600" swimtime="00:10:03.34" />
                    <SPLIT distance="650" swimtime="00:10:55.91" />
                    <SPLIT distance="700" swimtime="00:11:48.17" />
                    <SPLIT distance="750" swimtime="00:12:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="375" swimtime="00:00:42.91" resultid="1884" heatid="4648" lane="1" entrytime="00:00:39.50" />
                <RESULT eventid="1320" points="404" swimtime="00:01:20.41" resultid="1885" heatid="4668" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="340" swimtime="00:01:37.58" resultid="1886" heatid="4711" lane="0" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="385" swimtime="00:02:57.71" resultid="1887" heatid="4721" lane="8" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:25.34" />
                    <SPLIT distance="150" swimtime="00:02:12.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="330" swimtime="00:03:39.31" resultid="1888" heatid="4747" lane="5" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.66" />
                    <SPLIT distance="100" swimtime="00:01:47.11" />
                    <SPLIT distance="150" swimtime="00:02:45.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="363" swimtime="00:06:29.10" resultid="1889" heatid="4799" lane="8" entrytime="00:06:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                    <SPLIT distance="100" swimtime="00:01:29.86" />
                    <SPLIT distance="150" swimtime="00:02:19.37" />
                    <SPLIT distance="200" swimtime="00:03:09.62" />
                    <SPLIT distance="250" swimtime="00:04:00.34" />
                    <SPLIT distance="300" swimtime="00:04:51.19" />
                    <SPLIT distance="350" swimtime="00:05:42.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Genowefa" lastname="Drużyńska" birthdate="1951-02-19" gender="F" nation="POL" license="102611600033" athleteid="1897">
              <RESULTS>
                <RESULT eventid="1059" points="176" swimtime="00:00:54.82" resultid="1898" heatid="4596" lane="5" entrytime="00:00:58.00" />
                <RESULT eventid="1234" points="148" swimtime="00:01:05.36" resultid="1899" heatid="4640" lane="3" entrytime="00:01:06.00" />
                <RESULT eventid="1404" points="182" swimtime="00:02:49.06" resultid="1900" heatid="4685" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="136" swimtime="00:01:07.90" resultid="1901" heatid="4694" lane="2" />
                <RESULT eventid="1684" points="198" swimtime="00:01:11.49" resultid="1902" heatid="4751" lane="5" entrytime="00:01:06.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beata" lastname="Sulewska" birthdate="1972-11-02" gender="F" nation="POL" license="102611600016" athleteid="1890">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="1891" heatid="4600" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1158" points="653" swimtime="00:11:01.48" resultid="1892" heatid="4632" lane="6" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="150" swimtime="00:01:59.50" />
                    <SPLIT distance="200" swimtime="00:02:40.69" />
                    <SPLIT distance="250" swimtime="00:03:22.06" />
                    <SPLIT distance="300" swimtime="00:04:03.65" />
                    <SPLIT distance="350" swimtime="00:04:45.59" />
                    <SPLIT distance="400" swimtime="00:05:27.30" />
                    <SPLIT distance="450" swimtime="00:06:09.44" />
                    <SPLIT distance="500" swimtime="00:06:51.44" />
                    <SPLIT distance="550" swimtime="00:07:33.37" />
                    <SPLIT distance="600" swimtime="00:08:15.51" />
                    <SPLIT distance="650" swimtime="00:08:57.69" />
                    <SPLIT distance="700" swimtime="00:09:39.86" />
                    <SPLIT distance="750" swimtime="00:10:17.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1269" points="674" swimtime="00:03:07.75" resultid="1893" heatid="4654" lane="8" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                    <SPLIT distance="100" swimtime="00:01:31.26" />
                    <SPLIT distance="150" swimtime="00:02:20.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="657" swimtime="00:01:26.77" resultid="1894" heatid="4688" lane="9" entrytime="00:01:26.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="651" swimtime="00:02:33.64" resultid="1895" heatid="4717" lane="0" entrytime="00:02:31.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                    <SPLIT distance="150" swimtime="00:01:55.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="648" swimtime="00:05:24.22" resultid="1896" heatid="4791" lane="8" entrytime="00:05:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:17.26" />
                    <SPLIT distance="150" swimtime="00:01:58.19" />
                    <SPLIT distance="200" swimtime="00:02:39.84" />
                    <SPLIT distance="250" swimtime="00:03:21.56" />
                    <SPLIT distance="300" swimtime="00:04:03.23" />
                    <SPLIT distance="350" swimtime="00:04:44.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01203" nation="POL" region="03" clubid="1833" name="UKS TRÓJKA Puławy" shortname="TRÓJKA Puławy">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Maciejczak" birthdate="1960-07-08" gender="M" nation="POL" athleteid="1838">
              <RESULTS>
                <RESULT eventid="1216" points="292" swimtime="00:27:01.52" resultid="1839" heatid="4638" lane="2" entrytime="00:27:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:35.47" />
                    <SPLIT distance="150" swimtime="00:02:27.35" />
                    <SPLIT distance="200" swimtime="00:03:21.05" />
                    <SPLIT distance="250" swimtime="00:04:14.74" />
                    <SPLIT distance="300" swimtime="00:05:09.66" />
                    <SPLIT distance="350" swimtime="00:06:01.64" />
                    <SPLIT distance="400" swimtime="00:06:56.74" />
                    <SPLIT distance="450" swimtime="00:07:49.38" />
                    <SPLIT distance="500" swimtime="00:08:44.91" />
                    <SPLIT distance="550" swimtime="00:09:38.35" />
                    <SPLIT distance="600" swimtime="00:10:33.44" />
                    <SPLIT distance="650" swimtime="00:11:28.40" />
                    <SPLIT distance="700" swimtime="00:12:22.96" />
                    <SPLIT distance="750" swimtime="00:13:18.31" />
                    <SPLIT distance="800" swimtime="00:14:12.50" />
                    <SPLIT distance="850" swimtime="00:15:07.58" />
                    <SPLIT distance="900" swimtime="00:16:01.29" />
                    <SPLIT distance="950" swimtime="00:16:56.07" />
                    <SPLIT distance="1000" swimtime="00:17:50.46" />
                    <SPLIT distance="1050" swimtime="00:18:45.63" />
                    <SPLIT distance="1100" swimtime="00:19:40.69" />
                    <SPLIT distance="1150" swimtime="00:20:36.90" />
                    <SPLIT distance="1200" swimtime="00:21:29.36" />
                    <SPLIT distance="1250" swimtime="00:22:26.49" />
                    <SPLIT distance="1300" swimtime="00:23:20.51" />
                    <SPLIT distance="1350" swimtime="00:24:16.32" />
                    <SPLIT distance="1400" swimtime="00:25:11.35" />
                    <SPLIT distance="1450" swimtime="00:26:06.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="305" swimtime="00:01:25.64" resultid="1840" heatid="4667" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="186" swimtime="00:08:59.50" resultid="1841" heatid="4789" lane="1" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.69" />
                    <SPLIT distance="100" swimtime="00:02:05.57" />
                    <SPLIT distance="150" swimtime="00:03:21.94" />
                    <SPLIT distance="200" swimtime="00:04:33.16" />
                    <SPLIT distance="250" swimtime="00:06:01.06" />
                    <SPLIT distance="300" swimtime="00:07:24.13" />
                    <SPLIT distance="350" swimtime="00:08:11.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="320" swimtime="00:06:41.75" resultid="1842" heatid="4800" lane="1" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                    <SPLIT distance="150" swimtime="00:02:21.29" />
                    <SPLIT distance="200" swimtime="00:03:13.41" />
                    <SPLIT distance="250" swimtime="00:04:07.43" />
                    <SPLIT distance="300" swimtime="00:04:59.24" />
                    <SPLIT distance="350" swimtime="00:05:52.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" athleteid="1834">
              <RESULTS>
                <RESULT eventid="1216" points="518" swimtime="00:20:43.49" resultid="1835" heatid="4638" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                    <SPLIT distance="150" swimtime="00:01:58.39" />
                    <SPLIT distance="200" swimtime="00:02:40.60" />
                    <SPLIT distance="250" swimtime="00:03:22.64" />
                    <SPLIT distance="300" swimtime="00:04:04.48" />
                    <SPLIT distance="350" swimtime="00:04:45.69" />
                    <SPLIT distance="400" swimtime="00:05:27.30" />
                    <SPLIT distance="450" swimtime="00:06:08.49" />
                    <SPLIT distance="500" swimtime="00:06:49.63" />
                    <SPLIT distance="550" swimtime="00:07:31.31" />
                    <SPLIT distance="600" swimtime="00:08:12.86" />
                    <SPLIT distance="650" swimtime="00:08:54.40" />
                    <SPLIT distance="700" swimtime="00:09:35.93" />
                    <SPLIT distance="750" swimtime="00:10:17.59" />
                    <SPLIT distance="800" swimtime="00:10:59.01" />
                    <SPLIT distance="850" swimtime="00:11:40.27" />
                    <SPLIT distance="900" swimtime="00:12:21.83" />
                    <SPLIT distance="950" swimtime="00:13:03.76" />
                    <SPLIT distance="1000" swimtime="00:13:45.66" />
                    <SPLIT distance="1050" swimtime="00:14:28.03" />
                    <SPLIT distance="1100" swimtime="00:15:10.26" />
                    <SPLIT distance="1150" swimtime="00:15:52.09" />
                    <SPLIT distance="1200" swimtime="00:16:34.48" />
                    <SPLIT distance="1250" swimtime="00:17:16.74" />
                    <SPLIT distance="1300" swimtime="00:17:58.73" />
                    <SPLIT distance="1350" swimtime="00:18:40.95" />
                    <SPLIT distance="1400" swimtime="00:19:22.80" />
                    <SPLIT distance="1450" swimtime="00:20:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="557" swimtime="00:02:34.28" resultid="1836" heatid="4681" lane="1" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:14.99" />
                    <SPLIT distance="150" swimtime="00:01:55.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="589" swimtime="00:01:07.80" resultid="1837" heatid="4740" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01911" nation="POL" region="11" clubid="2301" name="RMKS Rybnik">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Duda" birthdate="1981-04-15" gender="F" nation="POL" athleteid="2302">
              <RESULTS>
                <RESULT eventid="1059" points="741" swimtime="00:00:29.21" resultid="2303" heatid="4601" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1107" points="603" swimtime="00:02:51.61" resultid="2304" heatid="4621" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:22.05" />
                    <SPLIT distance="150" swimtime="00:02:15.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="501" swimtime="00:00:37.29" resultid="2305" heatid="4642" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1303" points="657" swimtime="00:01:06.75" resultid="2306" heatid="4663" lane="0" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="757" swimtime="00:00:31.11" resultid="2307" heatid="4697" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1573" points="488" swimtime="00:06:33.53" resultid="2308" heatid="4786" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:01:29.45" />
                    <SPLIT distance="150" swimtime="00:02:24.55" />
                    <SPLIT distance="200" swimtime="00:03:15.94" />
                    <SPLIT distance="250" swimtime="00:04:13.50" />
                    <SPLIT distance="300" swimtime="00:05:09.74" />
                    <SPLIT distance="350" swimtime="00:05:54.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="545" swimtime="00:01:17.54" resultid="2309" heatid="4736" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="494" swimtime="00:00:41.00" resultid="2310" heatid="4754" lane="1" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAOPO" nation="POL" region="07" clubid="2995" name="T.P. MASTERS Opole" shortname="MASTERS Opole">
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Januszkiewicz" birthdate="1962-08-18" gender="M" nation="POL" athleteid="3001">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1490" points="874" swimtime="00:01:09.10" resultid="3002" heatid="4713" lane="9" entrytime="00:01:09.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1667" points="921" swimtime="00:02:30.15" resultid="3003" heatid="4750" lane="1" entrytime="00:02:32.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:13.05" />
                    <SPLIT distance="150" swimtime="00:01:51.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Mandziuk" birthdate="1965-04-11" gender="M" nation="POL" athleteid="2996">
              <RESULTS>
                <RESULT eventid="1090" points="326" swimtime="00:00:35.49" resultid="2997" heatid="4607" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1320" points="325" swimtime="00:01:21.45" resultid="2998" heatid="4667" lane="7" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="175" swimtime="00:02:00.86" resultid="2999" heatid="4691" lane="9" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="170" swimtime="00:00:54.09" resultid="3000" heatid="4757" lane="6" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05911" nation="POL" region="11" clubid="1810" name="UKS KARLIK Katowice" shortname="KARLIK Katowice">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Szczypiński" birthdate="1986-12-05" gender="M" nation="POL" athleteid="1811">
              <RESULTS>
                <RESULT eventid="1090" points="615" swimtime="00:00:26.76" resultid="1812" heatid="4615" lane="9" entrytime="00:00:26.80" />
                <RESULT eventid="1182" points="576" swimtime="00:09:59.01" resultid="1813" heatid="4636" lane="7" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:07.91" />
                    <SPLIT distance="150" swimtime="00:01:46.19" />
                    <SPLIT distance="200" swimtime="00:02:24.75" />
                    <SPLIT distance="250" swimtime="00:03:03.41" />
                    <SPLIT distance="300" swimtime="00:03:42.31" />
                    <SPLIT distance="350" swimtime="00:04:20.70" />
                    <SPLIT distance="400" swimtime="00:04:58.98" />
                    <SPLIT distance="450" swimtime="00:05:37.26" />
                    <SPLIT distance="500" swimtime="00:06:15.52" />
                    <SPLIT distance="550" swimtime="00:06:53.24" />
                    <SPLIT distance="600" swimtime="00:07:31.17" />
                    <SPLIT distance="650" swimtime="00:08:08.90" />
                    <SPLIT distance="700" swimtime="00:08:46.23" />
                    <SPLIT distance="750" swimtime="00:09:23.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MALUB" nation="POL" region="03" clubid="2231" name="MASTERS Lublin">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Wójcicka" birthdate="1975-04-28" gender="F" nation="POL" license="103503600002" athleteid="2232">
              <RESULTS>
                <RESULT eventid="1234" points="447" swimtime="00:00:40.55" resultid="2233" heatid="4642" lane="8" entrytime="00:00:40.48" entrycourse="LCM" />
                <RESULT eventid="1473" points="399" swimtime="00:01:31.00" resultid="2234" heatid="4707" lane="1" entrytime="00:01:40.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Ćwikła" birthdate="1975-11-07" gender="M" nation="POL" license="103503700005" athleteid="2239">
              <RESULTS>
                <RESULT eventid="1252" points="413" swimtime="00:00:37.06" resultid="2240" heatid="4649" lane="9" entrytime="00:00:36.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Molenda" birthdate="1971-12-11" gender="M" nation="POL" license="103503700012" athleteid="2241">
              <RESULTS>
                <RESULT eventid="1090" points="294" swimtime="00:00:36.19" resultid="2242" heatid="4606" lane="3" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1320" points="286" swimtime="00:01:22.12" resultid="2243" heatid="4667" lane="1" entrytime="00:01:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="250" swimtime="00:00:41.08" resultid="2244" heatid="4699" lane="0" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1524" points="238" swimtime="00:03:11.26" resultid="2245" heatid="4720" lane="6" entrytime="00:03:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:01:29.76" />
                    <SPLIT distance="150" swimtime="00:02:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="156" swimtime="00:01:46.25" resultid="2246" heatid="4738" lane="3" entrytime="00:01:48.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Dawidek" birthdate="1986-03-13" gender="M" nation="POL" license="103503700029" athleteid="2235">
              <RESULTS>
                <RESULT eventid="1124" points="357" swimtime="00:02:57.09" resultid="2236" heatid="4626" lane="8" entrytime="00:02:50.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:02:12.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="514" swimtime="00:01:03.36" resultid="2237" heatid="4672" lane="4" entrytime="00:01:02.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" status="DNS" swimtime="00:00:00.00" resultid="2238" heatid="4703" lane="1" entrytime="00:00:29.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Staszek" birthdate="1976-02-23" gender="M" nation="POL" license="103503700013" athleteid="2247">
              <RESULTS>
                <RESULT eventid="1090" points="328" swimtime="00:00:34.14" resultid="2248" heatid="4608" lane="5" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1320" points="288" swimtime="00:01:19.04" resultid="2249" heatid="4669" lane="4" entrytime="00:01:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="323" swimtime="00:01:34.36" resultid="2250" heatid="4691" lane="2" entrytime="00:01:33.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" status="DNS" swimtime="00:00:00.00" resultid="2251" heatid="4700" lane="9" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1701" points="336" swimtime="00:00:42.02" resultid="2252" heatid="4759" lane="3" entrytime="00:00:38.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="374" swimtime="00:02:26.29" resultid="2253" heatid="4684" lane="0" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:20.10" />
                    <SPLIT distance="150" swimtime="00:01:50.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2239" number="1" />
                    <RELAYPOSITION athleteid="2247" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="2235" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="2241" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MTM" nation="POL" region="14" clubid="2262" name="MASTERS Tomaszów Mazowiecki">
          <ATHLETES>
            <ATHLETE firstname="Barbara" lastname="Bucholz" birthdate="1973-12-01" gender="F" nation="POL" athleteid="2272">
              <RESULTS>
                <RESULT eventid="1107" points="176" swimtime="00:04:29.37" resultid="2273" heatid="4619" lane="9" entrytime="00:04:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.27" />
                    <SPLIT distance="100" swimtime="00:02:12.93" />
                    <SPLIT distance="150" swimtime="00:03:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="169" swimtime="00:04:57.61" resultid="2274" heatid="4652" lane="7" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.89" />
                    <SPLIT distance="100" swimtime="00:02:25.02" />
                    <SPLIT distance="150" swimtime="00:03:43.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="150" swimtime="00:01:53.47" resultid="2275" heatid="4659" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="182" swimtime="00:02:12.94" resultid="2276" heatid="4686" lane="9" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="174" swimtime="00:03:58.49" resultid="2277" heatid="4714" lane="5" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.71" />
                    <SPLIT distance="100" swimtime="00:01:56.04" />
                    <SPLIT distance="150" swimtime="00:02:58.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1615" points="127" swimtime="00:02:14.66" resultid="2278" heatid="4735" lane="7" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="177" swimtime="00:08:19.27" resultid="2279" heatid="4794" lane="4" entrytime="00:08:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.17" />
                    <SPLIT distance="100" swimtime="00:01:58.44" />
                    <SPLIT distance="150" swimtime="00:03:01.99" />
                    <SPLIT distance="200" swimtime="00:04:07.14" />
                    <SPLIT distance="250" swimtime="00:05:12.11" />
                    <SPLIT distance="300" swimtime="00:06:16.41" />
                    <SPLIT distance="350" swimtime="00:07:20.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Bucholz" birthdate="1972-01-26" gender="M" nation="POL" athleteid="2263">
              <RESULTS>
                <RESULT eventid="1124" points="388" swimtime="00:02:59.68" resultid="2264" heatid="4626" lane="0" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:28.41" />
                    <SPLIT distance="150" swimtime="00:02:19.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="539" swimtime="00:21:02.84" resultid="2265" heatid="4639" lane="7" entrytime="00:21:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:16.80" />
                    <SPLIT distance="150" swimtime="00:01:58.83" />
                    <SPLIT distance="200" swimtime="00:02:41.13" />
                    <SPLIT distance="250" swimtime="00:03:22.93" />
                    <SPLIT distance="300" swimtime="00:04:05.33" />
                    <SPLIT distance="350" swimtime="00:04:47.77" />
                    <SPLIT distance="400" swimtime="00:05:30.24" />
                    <SPLIT distance="450" swimtime="00:06:12.38" />
                    <SPLIT distance="500" swimtime="00:06:54.94" />
                    <SPLIT distance="550" swimtime="00:07:37.71" />
                    <SPLIT distance="600" swimtime="00:08:20.30" />
                    <SPLIT distance="650" swimtime="00:09:02.70" />
                    <SPLIT distance="700" swimtime="00:09:45.70" />
                    <SPLIT distance="750" swimtime="00:10:28.14" />
                    <SPLIT distance="800" swimtime="00:11:10.59" />
                    <SPLIT distance="850" swimtime="00:11:52.89" />
                    <SPLIT distance="900" swimtime="00:12:36.04" />
                    <SPLIT distance="950" swimtime="00:13:19.03" />
                    <SPLIT distance="1000" swimtime="00:14:02.12" />
                    <SPLIT distance="1050" swimtime="00:14:45.06" />
                    <SPLIT distance="1100" swimtime="00:15:27.52" />
                    <SPLIT distance="1150" swimtime="00:16:10.13" />
                    <SPLIT distance="1200" swimtime="00:16:52.66" />
                    <SPLIT distance="1250" swimtime="00:17:34.52" />
                    <SPLIT distance="1300" swimtime="00:18:17.31" />
                    <SPLIT distance="1350" swimtime="00:18:58.86" />
                    <SPLIT distance="1400" swimtime="00:19:41.59" />
                    <SPLIT distance="1450" swimtime="00:20:23.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="380" swimtime="00:03:19.34" resultid="2266" heatid="4656" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                    <SPLIT distance="100" swimtime="00:01:35.35" />
                    <SPLIT distance="150" swimtime="00:02:26.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="256" swimtime="00:03:29.83" resultid="2267" heatid="4679" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.35" />
                    <SPLIT distance="100" swimtime="00:01:40.97" />
                    <SPLIT distance="150" swimtime="00:02:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="297" swimtime="00:02:57.76" resultid="2268" heatid="4722" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:24.64" />
                    <SPLIT distance="150" swimtime="00:02:11.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="410" swimtime="00:06:24.40" resultid="2269" heatid="4788" lane="7" entrytime="00:07:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                    <SPLIT distance="100" swimtime="00:01:41.79" />
                    <SPLIT distance="150" swimtime="00:02:29.20" />
                    <SPLIT distance="200" swimtime="00:03:16.02" />
                    <SPLIT distance="250" swimtime="00:04:09.47" />
                    <SPLIT distance="300" swimtime="00:05:03.39" />
                    <SPLIT distance="350" swimtime="00:05:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" status="DNS" swimtime="00:00:00.00" resultid="2270" heatid="4738" lane="5" entrytime="00:01:42.00" />
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="2271" heatid="4797" lane="3" entrytime="00:05:16.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01304" nation="POL" region="04" clubid="2163" name="LANDSBERG CREW Gorzów Wlkp.">
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Kaczmarek" birthdate="1992-08-23" gender="F" nation="POL" license="501304600002" athleteid="2164">
              <RESULTS>
                <RESULT eventid="1059" points="714" swimtime="00:00:28.79" resultid="2165" heatid="4602" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1107" points="610" swimtime="00:02:37.86" resultid="2166" heatid="4621" lane="6" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:16.11" />
                    <SPLIT distance="150" swimtime="00:02:02.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="479" swimtime="00:03:10.24" resultid="2167" heatid="4654" lane="6" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                    <SPLIT distance="100" swimtime="00:01:34.19" />
                    <SPLIT distance="150" swimtime="00:02:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="690" swimtime="00:01:02.50" resultid="2168" heatid="4663" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" points="665" swimtime="00:02:20.15" resultid="2169" heatid="4717" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:45.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1573" points="667" swimtime="00:05:38.87" resultid="2170" heatid="4785" lane="5" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="150" swimtime="00:02:05.70" />
                    <SPLIT distance="200" swimtime="00:02:51.39" />
                    <SPLIT distance="250" swimtime="00:03:38.04" />
                    <SPLIT distance="300" swimtime="00:04:25.60" />
                    <SPLIT distance="350" swimtime="00:05:03.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1650" points="534" swimtime="00:02:49.56" resultid="2171" heatid="4745" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:23.27" />
                    <SPLIT distance="150" swimtime="00:02:06.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" points="597" swimtime="00:05:07.11" resultid="2172" heatid="4791" lane="5" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:01:53.56" />
                    <SPLIT distance="200" swimtime="00:02:32.93" />
                    <SPLIT distance="250" swimtime="00:03:11.60" />
                    <SPLIT distance="300" swimtime="00:03:51.07" />
                    <SPLIT distance="350" swimtime="00:04:30.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Kaczmarek" birthdate="1979-01-26" gender="M" nation="POL" license="501304600002" athleteid="2173">
              <RESULTS>
                <RESULT eventid="1124" points="636" swimtime="00:02:31.86" resultid="2174" heatid="4628" lane="8" entrytime="00:02:28.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:13.90" />
                    <SPLIT distance="150" swimtime="00:01:57.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="582" swimtime="00:10:17.52" resultid="2175" heatid="4636" lane="3" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="150" swimtime="00:01:52.29" />
                    <SPLIT distance="200" swimtime="00:02:31.25" />
                    <SPLIT distance="250" swimtime="00:03:10.71" />
                    <SPLIT distance="300" swimtime="00:03:49.91" />
                    <SPLIT distance="350" swimtime="00:04:29.15" />
                    <SPLIT distance="400" swimtime="00:05:08.25" />
                    <SPLIT distance="450" swimtime="00:05:47.37" />
                    <SPLIT distance="500" swimtime="00:06:26.26" />
                    <SPLIT distance="550" swimtime="00:07:05.67" />
                    <SPLIT distance="600" swimtime="00:07:44.69" />
                    <SPLIT distance="650" swimtime="00:08:23.84" />
                    <SPLIT distance="700" swimtime="00:09:02.10" />
                    <SPLIT distance="750" swimtime="00:09:39.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="526" swimtime="00:02:51.65" resultid="2176" heatid="4658" lane="8" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:26.08" />
                    <SPLIT distance="150" swimtime="00:02:10.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1354" points="473" swimtime="00:02:41.08" resultid="2177" heatid="4681" lane="6" entrytime="00:02:28.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                    <SPLIT distance="150" swimtime="00:01:57.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="593" swimtime="00:02:15.27" resultid="2178" heatid="4724" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="150" swimtime="00:01:41.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1597" points="604" swimtime="00:05:34.61" resultid="2179" heatid="4787" lane="6" entrytime="00:05:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                    <SPLIT distance="150" swimtime="00:01:59.82" />
                    <SPLIT distance="200" swimtime="00:02:45.42" />
                    <SPLIT distance="250" swimtime="00:03:33.03" />
                    <SPLIT distance="300" swimtime="00:04:20.87" />
                    <SPLIT distance="350" swimtime="00:04:58.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="508" swimtime="00:02:40.46" resultid="2180" heatid="4750" lane="0" entrytime="00:02:36.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:02:00.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="604" swimtime="00:04:51.86" resultid="2181" heatid="4795" lane="8" entrytime="00:04:44.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                    <SPLIT distance="150" swimtime="00:01:47.78" />
                    <SPLIT distance="200" swimtime="00:02:25.42" />
                    <SPLIT distance="250" swimtime="00:03:02.25" />
                    <SPLIT distance="300" swimtime="00:03:39.20" />
                    <SPLIT distance="350" swimtime="00:04:16.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04901" nation="POL" region="01" clubid="3764" name="KS NEPTUN Świdnica" shortname="NEPTUN Świdnica">
          <ATHLETES>
            <ATHLETE firstname="Bartłomiej" lastname="Żukowski" birthdate="1993-04-26" gender="M" nation="POL" license="104901700097" athleteid="3765">
              <RESULTS>
                <RESULT eventid="1090" points="749" swimtime="00:00:24.36" resultid="3766" heatid="4617" lane="8" entrytime="00:00:24.50" />
                <RESULT eventid="1422" points="784" swimtime="00:01:06.40" resultid="3767" heatid="4693" lane="5" entrytime="00:01:06.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="834" swimtime="00:00:29.47" resultid="3768" heatid="4762" lane="4" entrytime="00:00:28.91" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02211" nation="POL" region="11" clubid="3859" name="MUKS GILUS Gilowice" shortname="GILUS Gilowice">
          <ATHLETES>
            <ATHLETE firstname="Sławomir" lastname="Formas" birthdate="1969-11-05" gender="M" nation="POL" license="502211700187" athleteid="3860">
              <RESULTS>
                <RESULT eventid="1286" points="765" swimtime="00:02:37.89" resultid="3861" heatid="4658" lane="6" entrytime="00:02:36.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:16.45" />
                    <SPLIT distance="150" swimtime="00:01:57.83" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1422" points="854" swimtime="00:01:09.67" resultid="3862" heatid="4693" lane="2" entrytime="00:01:10.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="650" swimtime="00:01:06.04" resultid="3863" heatid="4740" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski MASTERS" eventid="1701" points="895" swimtime="00:00:31.02" resultid="3864" heatid="4762" lane="1" entrytime="00:00:31.04" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00303" nation="POL" region="03" clubid="2768" name="MASTERS AVIA Świdnik">
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Kędzierska" birthdate="1987-11-20" gender="F" nation="POL" license="504303600016" athleteid="2778">
              <RESULTS>
                <RESULT eventid="1404" points="500" swimtime="00:01:28.77" resultid="2779" heatid="4686" lane="7" entrytime="00:02:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Sitkowski" birthdate="1974-10-05" gender="M" nation="POL" license="504303700001" athleteid="2769">
              <RESULTS>
                <RESULT eventid="1090" points="610" swimtime="00:00:27.76" resultid="2770" heatid="4613" lane="7" entrytime="00:00:28.14" entrycourse="LCM" />
                <RESULT eventid="1252" points="552" swimtime="00:00:33.65" resultid="2771" heatid="4649" lane="4" entrytime="00:00:33.28" entrycourse="LCM" />
                <RESULT eventid="1490" points="529" swimtime="00:01:14.32" resultid="2772" heatid="4712" lane="7" entrytime="00:01:14.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="442" swimtime="00:02:52.70" resultid="2773" heatid="4749" lane="0" entrytime="00:02:54.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                    <SPLIT distance="150" swimtime="00:02:07.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Stypiński" birthdate="1956-04-17" gender="M" nation="POL" license="504303700015" athleteid="2800">
              <RESULTS>
                <RESULT eventid="1090" points="554" swimtime="00:00:31.90" resultid="2801" heatid="4609" lane="9" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1252" points="461" swimtime="00:00:40.04" resultid="2802" heatid="4648" lane="3" entrytime="00:00:38.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Lis" birthdate="1998-03-11" gender="M" nation="POL" license="104303700013" athleteid="2780">
              <RESULTS>
                <RESULT eventid="1090" points="661" swimtime="00:00:25.59" resultid="2781" heatid="4616" lane="7" entrytime="00:00:25.50" entrycourse="LCM" />
                <RESULT eventid="1252" points="574" swimtime="00:00:30.60" resultid="2782" heatid="4650" lane="7" entrytime="00:00:32.01" entrycourse="LCM" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2783" heatid="4674" lane="5" entrytime="00:00:56.70" entrycourse="LCM" />
                <RESULT eventid="1456" points="633" swimtime="00:00:27.61" resultid="2784" heatid="4705" lane="9" entrytime="00:00:26.50" entrycourse="LCM" />
                <RESULT eventid="1701" points="647" swimtime="00:00:31.46" resultid="2785" heatid="4762" lane="7" entrytime="00:00:31.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cezary" lastname="Lipiński" birthdate="1972-04-11" gender="M" nation="POL" license="104303700002" athleteid="2793">
              <RESULTS>
                <RESULT eventid="1090" points="574" swimtime="00:00:28.97" resultid="2794" heatid="4613" lane="8" entrytime="00:00:28.27" entrycourse="LCM" />
                <RESULT eventid="1216" points="581" swimtime="00:20:32.10" resultid="2795" heatid="4639" lane="5" entrytime="00:19:36.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                    <SPLIT distance="150" swimtime="00:01:54.45" />
                    <SPLIT distance="200" swimtime="00:02:34.60" />
                    <SPLIT distance="250" swimtime="00:03:15.62" />
                    <SPLIT distance="300" swimtime="00:03:55.56" />
                    <SPLIT distance="350" swimtime="00:04:36.47" />
                    <SPLIT distance="400" swimtime="00:05:16.99" />
                    <SPLIT distance="450" swimtime="00:05:57.03" />
                    <SPLIT distance="500" swimtime="00:06:38.17" />
                    <SPLIT distance="550" swimtime="00:07:19.16" />
                    <SPLIT distance="600" swimtime="00:08:00.33" />
                    <SPLIT distance="650" swimtime="00:08:41.40" />
                    <SPLIT distance="700" swimtime="00:09:22.87" />
                    <SPLIT distance="750" swimtime="00:10:03.74" />
                    <SPLIT distance="800" swimtime="00:10:45.23" />
                    <SPLIT distance="850" swimtime="00:11:26.51" />
                    <SPLIT distance="900" swimtime="00:12:08.05" />
                    <SPLIT distance="950" swimtime="00:12:50.09" />
                    <SPLIT distance="1000" swimtime="00:13:31.80" />
                    <SPLIT distance="1050" swimtime="00:14:13.36" />
                    <SPLIT distance="1100" swimtime="00:14:56.00" />
                    <SPLIT distance="1150" swimtime="00:15:38.72" />
                    <SPLIT distance="1200" swimtime="00:16:20.87" />
                    <SPLIT distance="1250" swimtime="00:17:02.77" />
                    <SPLIT distance="1300" swimtime="00:17:44.93" />
                    <SPLIT distance="1350" swimtime="00:18:26.94" />
                    <SPLIT distance="1400" swimtime="00:19:09.43" />
                    <SPLIT distance="1450" swimtime="00:19:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="609" swimtime="00:01:03.85" resultid="2796" heatid="4672" lane="6" entrytime="00:01:02.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="458" swimtime="00:00:33.56" resultid="2797" heatid="4701" lane="3" entrytime="00:00:32.81" entrycourse="LCM" />
                <RESULT eventid="1524" points="550" swimtime="00:02:24.76" resultid="2798" heatid="4723" lane="3" entrytime="00:02:20.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:10.76" />
                    <SPLIT distance="150" swimtime="00:01:48.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="562" swimtime="00:05:10.05" resultid="2799" heatid="4795" lane="9" entrytime="00:04:46.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                    <SPLIT distance="150" swimtime="00:01:52.13" />
                    <SPLIT distance="200" swimtime="00:02:31.39" />
                    <SPLIT distance="250" swimtime="00:03:10.76" />
                    <SPLIT distance="300" swimtime="00:03:51.13" />
                    <SPLIT distance="350" swimtime="00:04:31.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Mazur" birthdate="1995-03-13" gender="M" nation="POL" license="104303700009" athleteid="2774">
              <RESULTS>
                <RESULT eventid="1252" points="552" swimtime="00:00:31.01" resultid="2775" heatid="4650" lane="6" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1320" points="718" swimtime="00:00:56.32" resultid="2776" heatid="4675" lane="7" entrytime="00:00:55.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="620" swimtime="00:00:27.80" resultid="2777" heatid="4704" lane="5" entrytime="00:00:26.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Zielonka" birthdate="1986-05-26" gender="M" nation="POL" license="104303700006" athleteid="2786">
              <RESULTS>
                <RESULT eventid="1090" points="621" swimtime="00:00:26.67" resultid="2787" heatid="4615" lane="0" entrytime="00:00:26.52" entrycourse="LCM" />
                <RESULT eventid="1320" points="666" swimtime="00:00:58.14" resultid="2788" heatid="4674" lane="6" entrytime="00:00:57.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="576" swimtime="00:00:29.01" resultid="2789" heatid="4704" lane="9" entrytime="00:00:28.60" entrycourse="LCM" />
                <RESULT eventid="1524" points="593" swimtime="00:02:14.27" resultid="2790" heatid="4725" lane="8" entrytime="00:02:09.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="100" swimtime="00:01:05.21" />
                    <SPLIT distance="150" swimtime="00:01:39.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="480" swimtime="00:01:08.51" resultid="2791" heatid="4741" lane="1" entrytime="00:01:06.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" points="574" swimtime="00:04:55.86" resultid="2792" heatid="4795" lane="0" entrytime="00:04:44.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:11.17" />
                    <SPLIT distance="150" swimtime="00:01:48.56" />
                    <SPLIT distance="200" swimtime="00:02:26.78" />
                    <SPLIT distance="250" swimtime="00:03:04.75" />
                    <SPLIT distance="300" swimtime="00:03:42.74" />
                    <SPLIT distance="350" swimtime="00:04:20.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1565" points="637" swimtime="00:01:54.16" resultid="2803" heatid="4728" lane="1" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.63" />
                    <SPLIT distance="100" swimtime="00:00:58.68" />
                    <SPLIT distance="150" swimtime="00:01:28.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2769" number="1" />
                    <RELAYPOSITION athleteid="2800" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2793" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="2786" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT comment="K1 - Pływak wykonał kopnięcie delfinowe po pierwszym kopnięciu do stylu klasycznego (pierwszy ruch po starcie lub nawrocie)." eventid="1395" status="DSQ" swimtime="00:01:58.37" resultid="2804" heatid="4684" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:04.81" />
                    <SPLIT distance="150" swimtime="00:01:33.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2769" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2780" number="2" reactiontime="+24" status="DSQ" />
                    <RELAYPOSITION athleteid="2786" number="3" reactiontime="+36" status="DSQ" />
                    <RELAYPOSITION athleteid="2774" number="4" reactiontime="+7" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00116" nation="POL" region="16" clubid="1857" name="MKP Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Sławomir" lastname="Grzeszewski" birthdate="1953-09-25" gender="M" nation="POL" athleteid="1858">
              <RESULTS>
                <RESULT eventid="1124" points="399" swimtime="00:03:41.26" resultid="1859" heatid="4624" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:01:44.42" />
                    <SPLIT distance="150" swimtime="00:02:47.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="503" swimtime="00:03:52.31" resultid="1860" heatid="4657" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.71" />
                    <SPLIT distance="100" swimtime="00:01:53.22" />
                    <SPLIT distance="150" swimtime="00:02:54.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="492" swimtime="00:01:43.82" resultid="1861" heatid="4689" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1456" points="402" swimtime="00:00:40.61" resultid="1862" heatid="4699" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1701" points="580" swimtime="00:00:43.41" resultid="1863" heatid="4758" lane="6" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" region="14" clubid="1814" name="UKS DELFIN Legionowo" shortname="DELFIN Legionowo">
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Żbikowska" birthdate="1996-01-01" gender="F" nation="POL" license="S01414100028" athleteid="1821">
              <RESULTS>
                <RESULT eventid="1059" points="582" swimtime="00:00:30.43" resultid="1822" heatid="4601" lane="1" entrytime="00:00:30.58" />
                <RESULT eventid="1107" points="577" swimtime="00:02:48.96" resultid="1823" heatid="4620" lane="3" entrytime="00:02:56.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:20.60" />
                    <SPLIT distance="150" swimtime="00:02:06.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="590" swimtime="00:03:04.11" resultid="1824" heatid="4654" lane="9" entrytime="00:03:12.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                    <SPLIT distance="150" swimtime="00:02:18.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="555" swimtime="00:01:09.27" resultid="1825" heatid="4662" lane="3" entrytime="00:01:08.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="590" swimtime="00:01:24.12" resultid="1826" heatid="4688" lane="2" entrytime="00:01:23.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" status="DNS" swimtime="00:00:00.00" resultid="1827" heatid="4716" lane="4" entrytime="00:02:36.44" />
                <RESULT eventid="1684" points="589" swimtime="00:00:37.68" resultid="1828" heatid="4755" lane="1" entrytime="00:00:37.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Fajdasz" birthdate="1973-01-14" gender="M" nation="POL" license="101414700141" athleteid="1815">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="1816" heatid="4604" lane="1" />
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="1817" heatid="4644" lane="5" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="1818" heatid="4665" lane="0" />
                <RESULT eventid="1490" status="DNS" swimtime="00:00:00.00" resultid="1819" heatid="4709" lane="1" />
                <RESULT eventid="1667" status="DNS" swimtime="00:00:00.00" resultid="1820" heatid="4746" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Rapacki" birthdate="1978-05-18" gender="M" nation="POL" athleteid="1829">
              <RESULTS>
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)." eventid="1286" status="DSQ" swimtime="00:03:49.48" resultid="1830" heatid="4655" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.94" />
                    <SPLIT distance="100" swimtime="00:01:47.44" />
                    <SPLIT distance="150" swimtime="00:02:49.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="276" swimtime="00:01:39.38" resultid="1831" heatid="4690" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1701" points="341" swimtime="00:00:41.82" resultid="1832" heatid="4757" lane="9" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" region="11" clubid="3749" name="KS GÓRNIK Radlin" shortname="GÓRNIK Radlin">
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Kubica" birthdate="1972-02-22" gender="M" nation="POL" license="100211700343" athleteid="3750">
              <RESULTS>
                <RESULT eventid="1090" points="540" swimtime="00:00:29.57" resultid="3751" heatid="4604" lane="7" />
                <RESULT eventid="1216" points="415" swimtime="00:22:57.73" resultid="3752" heatid="4638" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:10.91" />
                    <SPLIT distance="200" swimtime="00:02:57.61" />
                    <SPLIT distance="250" swimtime="00:03:43.30" />
                    <SPLIT distance="300" swimtime="00:04:29.22" />
                    <SPLIT distance="350" swimtime="00:05:15.55" />
                    <SPLIT distance="400" swimtime="00:06:01.77" />
                    <SPLIT distance="450" swimtime="00:06:48.48" />
                    <SPLIT distance="500" swimtime="00:07:35.32" />
                    <SPLIT distance="550" swimtime="00:08:21.94" />
                    <SPLIT distance="600" swimtime="00:09:08.28" />
                    <SPLIT distance="650" swimtime="00:09:54.83" />
                    <SPLIT distance="700" swimtime="00:10:41.31" />
                    <SPLIT distance="750" swimtime="00:11:27.99" />
                    <SPLIT distance="800" swimtime="00:12:14.43" />
                    <SPLIT distance="850" swimtime="00:13:01.25" />
                    <SPLIT distance="900" swimtime="00:13:47.41" />
                    <SPLIT distance="950" swimtime="00:14:33.52" />
                    <SPLIT distance="1000" swimtime="00:15:19.99" />
                    <SPLIT distance="1050" swimtime="00:16:06.64" />
                    <SPLIT distance="1100" swimtime="00:16:52.97" />
                    <SPLIT distance="1150" swimtime="00:17:39.66" />
                    <SPLIT distance="1200" swimtime="00:18:25.72" />
                    <SPLIT distance="1250" swimtime="00:19:12.03" />
                    <SPLIT distance="1300" swimtime="00:19:57.67" />
                    <SPLIT distance="1350" swimtime="00:20:43.46" />
                    <SPLIT distance="1400" swimtime="00:21:28.81" />
                    <SPLIT distance="1450" swimtime="00:22:14.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="474" swimtime="00:00:36.65" resultid="3753" heatid="4644" lane="3" />
                <RESULT eventid="1354" status="DNS" swimtime="00:00:00.00" resultid="3754" heatid="4678" lane="3" />
                <RESULT eventid="1456" points="501" swimtime="00:00:32.57" resultid="3755" heatid="4698" lane="9" />
                <RESULT eventid="1490" points="457" swimtime="00:01:19.88" resultid="3756" heatid="4709" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1633" points="428" swimtime="00:01:15.93" resultid="3757" heatid="4737" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="398" swimtime="00:03:02.76" resultid="3758" heatid="4746" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:01:27.54" />
                    <SPLIT distance="150" swimtime="00:02:15.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" region="15" clubid="3902" name="UKS CITYZEN Poznań" shortname="CITYZEN Poznań">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Matyszczak" birthdate="1970-12-14" gender="M" nation="POL" license="503415700353" athleteid="3916">
              <RESULTS>
                <RESULT eventid="1090" points="463" swimtime="00:00:31.12" resultid="3917" heatid="4610" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1182" points="280" swimtime="00:13:37.02" resultid="3918" heatid="4634" lane="6" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:25.47" />
                    <SPLIT distance="150" swimtime="00:02:14.28" />
                    <SPLIT distance="200" swimtime="00:03:05.33" />
                    <SPLIT distance="250" swimtime="00:03:56.69" />
                    <SPLIT distance="300" swimtime="00:04:48.26" />
                    <SPLIT distance="350" swimtime="00:05:40.31" />
                    <SPLIT distance="400" swimtime="00:06:32.00" />
                    <SPLIT distance="450" swimtime="00:07:24.06" />
                    <SPLIT distance="500" swimtime="00:08:16.02" />
                    <SPLIT distance="550" swimtime="00:09:08.04" />
                    <SPLIT distance="600" swimtime="00:10:00.23" />
                    <SPLIT distance="650" swimtime="00:11:02.39" />
                    <SPLIT distance="700" swimtime="00:12:01.92" />
                    <SPLIT distance="750" swimtime="00:12:41.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="319" swimtime="00:00:41.82" resultid="3919" heatid="4648" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1320" points="406" swimtime="00:01:13.12" resultid="3920" heatid="4670" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="291" swimtime="00:01:32.89" resultid="3921" heatid="4711" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="315" swimtime="00:02:54.20" resultid="3922" heatid="4721" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:22.27" />
                    <SPLIT distance="150" swimtime="00:02:09.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="287" swimtime="00:03:23.82" resultid="3923" heatid="4748" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="100" swimtime="00:01:39.42" />
                    <SPLIT distance="150" swimtime="00:02:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1766" status="DNS" swimtime="00:00:00.00" resultid="3924" heatid="4798" lane="7" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rusłana" lastname="Dembecka" birthdate="1957-10-01" gender="F" nation="POL" license="503415600404" athleteid="3903">
              <RESULTS>
                <RESULT eventid="1059" points="144" swimtime="00:00:55.49" resultid="3904" heatid="4597" lane="2" entrytime="00:00:51.00" />
                <RESULT eventid="1234" points="127" swimtime="00:01:06.75" resultid="3905" heatid="4640" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1269" points="327" swimtime="00:04:39.44" resultid="3906" heatid="4652" lane="2" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.70" />
                    <SPLIT distance="100" swimtime="00:02:20.68" />
                    <SPLIT distance="150" swimtime="00:03:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="310" swimtime="00:02:13.15" resultid="3907" heatid="4686" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="127" swimtime="00:02:27.91" resultid="3908" heatid="4706" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="259" swimtime="00:01:02.86" resultid="3909" heatid="4752" lane="8" entrytime="00:00:56.00" />
                <RESULT eventid="1742" points="174" swimtime="00:09:19.70" resultid="3910" heatid="4794" lane="6" entrytime="00:09:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.11" />
                    <SPLIT distance="100" swimtime="00:02:08.97" />
                    <SPLIT distance="150" swimtime="00:03:19.82" />
                    <SPLIT distance="200" swimtime="00:04:31.29" />
                    <SPLIT distance="250" swimtime="00:05:43.15" />
                    <SPLIT distance="300" swimtime="00:06:55.29" />
                    <SPLIT distance="350" swimtime="00:08:08.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Łutowicz" birthdate="1950-08-23" gender="F" nation="POL" license="503415600183" athleteid="3911">
              <RESULTS>
                <RESULT eventid="1059" points="238" swimtime="00:00:49.57" resultid="3912" heatid="4597" lane="7" entrytime="00:00:52.00" />
                <RESULT eventid="1234" points="187" swimtime="00:01:00.57" resultid="3913" heatid="4640" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1303" points="181" swimtime="00:01:58.22" resultid="3914" heatid="4659" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1473" points="192" swimtime="00:02:13.84" resultid="3915" heatid="4706" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Boryski" birthdate="1951-03-05" gender="M" nation="POL" license="503415700180" athleteid="3938">
              <RESULTS>
                <RESULT eventid="1216" points="336" swimtime="00:29:23.00" resultid="3939" heatid="4638" lane="1" entrytime="00:29:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.18" />
                    <SPLIT distance="100" swimtime="00:01:48.94" />
                    <SPLIT distance="150" swimtime="00:02:49.55" />
                    <SPLIT distance="200" swimtime="00:03:49.43" />
                    <SPLIT distance="250" swimtime="00:04:48.24" />
                    <SPLIT distance="300" swimtime="00:05:48.97" />
                    <SPLIT distance="350" swimtime="00:06:47.42" />
                    <SPLIT distance="400" swimtime="00:07:45.34" />
                    <SPLIT distance="450" swimtime="00:08:45.18" />
                    <SPLIT distance="500" swimtime="00:09:44.30" />
                    <SPLIT distance="550" swimtime="00:10:43.78" />
                    <SPLIT distance="600" swimtime="00:11:43.14" />
                    <SPLIT distance="650" swimtime="00:12:42.86" />
                    <SPLIT distance="700" swimtime="00:13:42.72" />
                    <SPLIT distance="750" swimtime="00:14:41.68" />
                    <SPLIT distance="800" swimtime="00:15:39.62" />
                    <SPLIT distance="850" swimtime="00:16:38.58" />
                    <SPLIT distance="900" swimtime="00:17:38.19" />
                    <SPLIT distance="950" swimtime="00:18:37.65" />
                    <SPLIT distance="1000" swimtime="00:19:36.11" />
                    <SPLIT distance="1050" swimtime="00:20:34.91" />
                    <SPLIT distance="1100" swimtime="00:21:33.84" />
                    <SPLIT distance="1150" swimtime="00:22:32.97" />
                    <SPLIT distance="1200" swimtime="00:23:32.10" />
                    <SPLIT distance="1250" swimtime="00:24:31.48" />
                    <SPLIT distance="1300" swimtime="00:25:30.32" />
                    <SPLIT distance="1350" swimtime="00:26:30.09" />
                    <SPLIT distance="1400" swimtime="00:27:28.76" />
                    <SPLIT distance="1450" swimtime="00:28:27.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="339" swimtime="00:00:48.15" resultid="3940" heatid="4646" lane="4" entrytime="00:00:46.00" />
                <RESULT eventid="1490" points="300" swimtime="00:01:49.75" resultid="3941" heatid="4710" lane="1" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="303" swimtime="00:03:58.48" resultid="3942" heatid="4747" lane="1" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.26" />
                    <SPLIT distance="100" swimtime="00:02:00.99" />
                    <SPLIT distance="150" swimtime="00:03:03.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Rybak-Starczak" birthdate="1975-01-16" gender="F" nation="POL" license="503415600144" athleteid="3933">
              <RESULTS>
                <RESULT eventid="1107" points="409" swimtime="00:03:10.44" resultid="3934" heatid="4620" lane="1" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:34.79" />
                    <SPLIT distance="150" swimtime="00:02:28.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="471" swimtime="00:03:30.43" resultid="3935" heatid="4653" lane="3" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                    <SPLIT distance="100" swimtime="00:01:42.14" />
                    <SPLIT distance="150" swimtime="00:02:38.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1404" points="443" swimtime="00:01:34.85" resultid="3936" heatid="4687" lane="7" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1684" points="431" swimtime="00:00:44.42" resultid="3937" heatid="4754" lane="0" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Pietraszewski" birthdate="1955-04-07" gender="M" nation="POL" license="503415700182" athleteid="3925">
              <RESULTS>
                <RESULT eventid="1090" points="279" swimtime="00:00:40.10" resultid="3926" heatid="4605" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1252" points="185" swimtime="00:00:54.31" resultid="3927" heatid="4646" lane="7" entrytime="00:00:54.00" />
                <RESULT eventid="1320" points="239" swimtime="00:01:35.80" resultid="3928" heatid="4666" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1490" points="204" swimtime="00:01:55.62" resultid="3929" heatid="4710" lane="0" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="229" swimtime="00:03:31.44" resultid="3930" heatid="4720" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.65" />
                    <SPLIT distance="100" swimtime="00:01:41.05" />
                    <SPLIT distance="150" swimtime="00:02:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1667" points="230" swimtime="00:04:07.23" resultid="3931" heatid="4747" lane="0" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.30" />
                    <SPLIT distance="100" swimtime="00:02:02.48" />
                    <SPLIT distance="150" swimtime="00:03:05.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1141" points="399" swimtime="00:02:35.53" resultid="3944" heatid="4629" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.50" />
                    <SPLIT distance="100" swimtime="00:01:28.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3911" number="1" />
                    <RELAYPOSITION athleteid="3925" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3933" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3916" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1718" points="230" swimtime="00:03:28.94" resultid="3945" heatid="4764" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.63" />
                    <SPLIT distance="100" swimtime="00:02:05.79" />
                    <SPLIT distance="150" swimtime="00:02:45.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3911" number="1" />
                    <RELAYPOSITION athleteid="3903" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="3916" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="3925" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03508" nation="POL" region="08" clubid="3769" name="KS PRESTIGE Rzeszów" shortname="PRESTIGE Rzeszów">
          <ATHLETES>
            <ATHLETE firstname="Patrycja" lastname="Rupa" birthdate="1996-01-11" gender="F" nation="POL" license="103508600006" athleteid="3770">
              <RESULTS>
                <RESULT eventid="1059" points="571" swimtime="00:00:30.63" resultid="3771" heatid="4596" lane="3" />
                <RESULT comment="Przekroczony limit czasu" eventid="1158" status="OTL" swimtime="00:12:16.70" resultid="3772" heatid="4631" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="100" swimtime="00:01:23.95" />
                    <SPLIT distance="150" swimtime="00:02:09.82" />
                    <SPLIT distance="200" swimtime="00:02:56.44" />
                    <SPLIT distance="250" swimtime="00:03:43.56" />
                    <SPLIT distance="300" swimtime="00:04:30.79" />
                    <SPLIT distance="350" swimtime="00:05:17.68" />
                    <SPLIT distance="400" swimtime="00:06:05.01" />
                    <SPLIT distance="450" swimtime="00:06:52.07" />
                    <SPLIT distance="500" swimtime="00:07:39.14" />
                    <SPLIT distance="550" swimtime="00:08:26.60" />
                    <SPLIT distance="600" swimtime="00:09:13.77" />
                    <SPLIT distance="650" swimtime="00:10:00.94" />
                    <SPLIT distance="700" swimtime="00:10:47.36" />
                    <SPLIT distance="750" swimtime="00:11:33.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="608" swimtime="00:00:33.51" resultid="3773" heatid="4640" lane="7" />
                <RESULT eventid="1269" status="DNS" swimtime="00:00:00.00" resultid="3774" heatid="4652" lane="1" />
                <RESULT eventid="1473" points="601" swimtime="00:01:12.96" resultid="3775" heatid="4706" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1507" status="DNS" swimtime="00:00:00.00" resultid="3776" heatid="4714" lane="6" />
                <RESULT eventid="1650" points="563" swimtime="00:02:41.23" resultid="3777" heatid="4743" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:19.63" />
                    <SPLIT distance="150" swimtime="00:02:00.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1742" status="DNS" swimtime="00:00:00.00" resultid="3778" heatid="4794" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SMS SwimArt Myslenice" version="Build 27713">
    <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Kraków" name="Mistrzostwa Polski w Pływaniu Masters" course="SCM" deadline="2013-11-05" hostclub.url="http://www.swimart.pl" nation="POL" organizer="Małopolski OZP" organizer.url="http://www.mozp.pl" result.url="http://www.omegatiming.pl" timing="AUTOMATIC">
      <AGEDATE value="2013-11-17" type="YEAR" />
      <POOL name="ZKP AWF Kraków" lanemin="1" lanemax="8" />
      <POINTTABLE pointtableid="1121" name="DSV Master Performance Table" version="2013" />
      <CONTACT email="zawody@swimart.pl" name="Artur Żak" phone="501 689 458" />
      <SESSIONS>
        <SESSION date="2013-11-15" daytime="16:00" name="MP Masters BLOK I" number="1" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="1059" daytime="16:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2567" />
                    <RANKING order="2" place="2" resultid="5149" />
                    <RANKING order="3" place="3" resultid="1967" />
                    <RANKING order="4" place="4" resultid="2606" />
                    <RANKING order="5" place="5" resultid="3902" />
                    <RANKING order="6" place="6" resultid="3777" />
                    <RANKING order="7" place="7" resultid="2994" />
                    <RANKING order="8" place="8" resultid="2061" />
                    <RANKING order="9" place="9" resultid="5574" />
                    <RANKING order="10" place="10" resultid="5107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4047" />
                    <RANKING order="2" place="2" resultid="3540" />
                    <RANKING order="3" place="3" resultid="2921" />
                    <RANKING order="4" place="4" resultid="2647" />
                    <RANKING order="5" place="5" resultid="2334" />
                    <RANKING order="6" place="6" resultid="6292" />
                    <RANKING order="7" place="7" resultid="5307" />
                    <RANKING order="8" place="8" resultid="3125" />
                    <RANKING order="9" place="-1" resultid="5566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4041" />
                    <RANKING order="2" place="2" resultid="5872" />
                    <RANKING order="3" place="3" resultid="3589" />
                    <RANKING order="4" place="4" resultid="5098" />
                    <RANKING order="5" place="5" resultid="4352" />
                    <RANKING order="6" place="6" resultid="3493" />
                    <RANKING order="7" place="7" resultid="4096" />
                    <RANKING order="8" place="8" resultid="5928" />
                    <RANKING order="9" place="9" resultid="3681" />
                    <RANKING order="10" place="10" resultid="3753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5407" />
                    <RANKING order="2" place="2" resultid="2934" />
                    <RANKING order="3" place="3" resultid="2941" />
                    <RANKING order="4" place="4" resultid="5129" />
                    <RANKING order="5" place="5" resultid="6202" />
                    <RANKING order="6" place="6" resultid="2228" />
                    <RANKING order="7" place="7" resultid="6692" />
                    <RANKING order="8" place="8" resultid="2956" />
                    <RANKING order="9" place="9" resultid="4018" />
                    <RANKING order="10" place="10" resultid="3486" />
                    <RANKING order="11" place="11" resultid="5898" />
                    <RANKING order="12" place="12" resultid="5279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1060" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4547" />
                    <RANKING order="2" place="2" resultid="5035" />
                    <RANKING order="3" place="3" resultid="3888" />
                    <RANKING order="4" place="4" resultid="6457" />
                    <RANKING order="5" place="5" resultid="2946" />
                    <RANKING order="6" place="6" resultid="3746" />
                    <RANKING order="7" place="7" resultid="2952" />
                    <RANKING order="8" place="8" resultid="4694" />
                    <RANKING order="9" place="9" resultid="3067" />
                    <RANKING order="10" place="9" resultid="5978" />
                    <RANKING order="11" place="11" resultid="6126" />
                    <RANKING order="12" place="12" resultid="6304" />
                    <RANKING order="13" place="13" resultid="4753" />
                    <RANKING order="14" place="-1" resultid="2376" />
                    <RANKING order="15" place="-1" resultid="6098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3712" />
                    <RANKING order="2" place="2" resultid="4366" />
                    <RANKING order="3" place="3" resultid="6320" />
                    <RANKING order="4" place="4" resultid="2844" />
                    <RANKING order="5" place="5" resultid="5370" />
                    <RANKING order="6" place="6" resultid="5488" />
                    <RANKING order="7" place="7" resultid="6778" />
                    <RANKING order="8" place="8" resultid="3967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4992" />
                    <RANKING order="2" place="2" resultid="2135" />
                    <RANKING order="3" place="3" resultid="4985" />
                    <RANKING order="4" place="4" resultid="3596" />
                    <RANKING order="5" place="5" resultid="3883" />
                    <RANKING order="6" place="6" resultid="4617" />
                    <RANKING order="7" place="7" resultid="3322" />
                    <RANKING order="8" place="8" resultid="2262" />
                    <RANKING order="9" place="9" resultid="3570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2127" />
                    <RANKING order="2" place="2" resultid="3729" />
                    <RANKING order="3" place="3" resultid="3396" />
                    <RANKING order="4" place="4" resultid="3924" />
                    <RANKING order="5" place="5" resultid="4350" />
                    <RANKING order="6" place="6" resultid="3559" />
                    <RANKING order="7" place="7" resultid="3140" />
                    <RANKING order="8" place="-1" resultid="3437" />
                    <RANKING order="9" place="-1" resultid="4600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4340" />
                    <RANKING order="2" place="2" resultid="6314" />
                    <RANKING order="3" place="3" resultid="5499" />
                    <RANKING order="4" place="4" resultid="4285" />
                    <RANKING order="5" place="5" resultid="5003" />
                    <RANKING order="6" place="6" resultid="4595" />
                    <RANKING order="7" place="7" resultid="3355" />
                    <RANKING order="8" place="8" resultid="5387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4671" />
                    <RANKING order="2" place="2" resultid="5770" />
                    <RANKING order="3" place="3" resultid="5393" />
                    <RANKING order="4" place="4" resultid="4354" />
                    <RANKING order="5" place="5" resultid="4053" />
                    <RANKING order="6" place="6" resultid="3820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4289" />
                    <RANKING order="2" place="2" resultid="3431" />
                    <RANKING order="3" place="3" resultid="6342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1073" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7671" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7672" daytime="16:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7673" daytime="16:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7674" daytime="16:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7675" daytime="16:07" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7676" daytime="16:08" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7677" daytime="16:09" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7678" daytime="16:11" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7679" daytime="16:12" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7680" daytime="16:13" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7681" daytime="16:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7682" daytime="16:16" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7683" daytime="16:17" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="16:19" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3561" />
                    <RANKING order="2" place="2" resultid="2577" />
                    <RANKING order="3" place="3" resultid="6241" />
                    <RANKING order="4" place="4" resultid="6265" />
                    <RANKING order="5" place="5" resultid="2294" />
                    <RANKING order="6" place="6" resultid="4758" />
                    <RANKING order="7" place="-1" resultid="2223" />
                    <RANKING order="8" place="-1" resultid="6210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5952" />
                    <RANKING order="2" place="2" resultid="5135" />
                    <RANKING order="3" place="3" resultid="3837" />
                    <RANKING order="4" place="4" resultid="6274" />
                    <RANKING order="5" place="5" resultid="4073" />
                    <RANKING order="6" place="6" resultid="5733" />
                    <RANKING order="7" place="7" resultid="3250" />
                    <RANKING order="8" place="8" resultid="2074" />
                    <RANKING order="9" place="9" resultid="3895" />
                    <RANKING order="10" place="10" resultid="2028" />
                    <RANKING order="11" place="10" resultid="5350" />
                    <RANKING order="12" place="12" resultid="3426" />
                    <RANKING order="13" place="13" resultid="3423" />
                    <RANKING order="14" place="14" resultid="2325" />
                    <RANKING order="15" place="15" resultid="2316" />
                    <RANKING order="16" place="16" resultid="3429" />
                    <RANKING order="17" place="17" resultid="5431" />
                    <RANKING order="18" place="18" resultid="5114" />
                    <RANKING order="19" place="19" resultid="3734" />
                    <RANKING order="20" place="20" resultid="3687" />
                    <RANKING order="21" place="-1" resultid="4064" />
                    <RANKING order="22" place="-1" resultid="4774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1871" />
                    <RANKING order="2" place="2" resultid="1905" />
                    <RANKING order="3" place="3" resultid="5961" />
                    <RANKING order="4" place="4" resultid="2066" />
                    <RANKING order="5" place="5" resultid="5599" />
                    <RANKING order="6" place="6" resultid="4069" />
                    <RANKING order="7" place="7" resultid="3775" />
                    <RANKING order="8" place="8" resultid="4107" />
                    <RANKING order="9" place="9" resultid="1992" />
                    <RANKING order="10" place="10" resultid="3582" />
                    <RANKING order="11" place="10" resultid="5731" />
                    <RANKING order="12" place="12" resultid="3863" />
                    <RANKING order="13" place="12" resultid="4190" />
                    <RANKING order="14" place="14" resultid="3517" />
                    <RANKING order="15" place="15" resultid="5561" />
                    <RANKING order="16" place="16" resultid="3245" />
                    <RANKING order="17" place="17" resultid="5628" />
                    <RANKING order="18" place="18" resultid="3237" />
                    <RANKING order="19" place="19" resultid="4058" />
                    <RANKING order="20" place="20" resultid="6261" />
                    <RANKING order="21" place="21" resultid="4079" />
                    <RANKING order="22" place="22" resultid="4175" />
                    <RANKING order="23" place="23" resultid="3527" />
                    <RANKING order="24" place="24" resultid="4185" />
                    <RANKING order="25" place="25" resultid="4162" />
                    <RANKING order="26" place="26" resultid="3675" />
                    <RANKING order="27" place="27" resultid="2329" />
                    <RANKING order="28" place="28" resultid="4179" />
                    <RANKING order="29" place="29" resultid="3738" />
                    <RANKING order="30" place="30" resultid="4196" />
                    <RANKING order="31" place="31" resultid="5297" />
                    <RANKING order="32" place="32" resultid="3523" />
                    <RANKING order="33" place="33" resultid="4363" />
                    <RANKING order="34" place="-1" resultid="5327" />
                    <RANKING order="35" place="-1" resultid="2033" />
                    <RANKING order="36" place="-1" resultid="5773" />
                    <RANKING order="37" place="-1" resultid="6269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6048" />
                    <RANKING order="2" place="2" resultid="2782" />
                    <RANKING order="3" place="3" resultid="3337" />
                    <RANKING order="4" place="4" resultid="2307" />
                    <RANKING order="5" place="5" resultid="2877" />
                    <RANKING order="6" place="6" resultid="2964" />
                    <RANKING order="7" place="7" resultid="1945" />
                    <RANKING order="8" place="8" resultid="5539" />
                    <RANKING order="9" place="9" resultid="5787" />
                    <RANKING order="10" place="10" resultid="4704" />
                    <RANKING order="11" place="11" resultid="2914" />
                    <RANKING order="12" place="12" resultid="1926" />
                    <RANKING order="13" place="13" resultid="4736" />
                    <RANKING order="14" place="14" resultid="2835" />
                    <RANKING order="15" place="15" resultid="2970" />
                    <RANKING order="16" place="16" resultid="5145" />
                    <RANKING order="17" place="17" resultid="1912" />
                    <RANKING order="18" place="18" resultid="2983" />
                    <RANKING order="19" place="19" resultid="4102" />
                    <RANKING order="20" place="20" resultid="6134" />
                    <RANKING order="21" place="21" resultid="2974" />
                    <RANKING order="22" place="22" resultid="3353" />
                    <RANKING order="23" place="23" resultid="2320" />
                    <RANKING order="24" place="24" resultid="3700" />
                    <RANKING order="25" place="25" resultid="3946" />
                    <RANKING order="26" place="26" resultid="5980" />
                    <RANKING order="27" place="27" resultid="6226" />
                    <RANKING order="28" place="28" resultid="3120" />
                    <RANKING order="29" place="29" resultid="3850" />
                    <RANKING order="30" place="-1" resultid="4781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2790" />
                    <RANKING order="2" place="2" resultid="3328" />
                    <RANKING order="3" place="3" resultid="5414" />
                    <RANKING order="4" place="4" resultid="3942" />
                    <RANKING order="5" place="5" resultid="3576" />
                    <RANKING order="6" place="6" resultid="3602" />
                    <RANKING order="7" place="7" resultid="2091" />
                    <RANKING order="8" place="7" resultid="5736" />
                    <RANKING order="9" place="9" resultid="6112" />
                    <RANKING order="10" place="10" resultid="5188" />
                    <RANKING order="11" place="11" resultid="2773" />
                    <RANKING order="12" place="12" resultid="4666" />
                    <RANKING order="13" place="13" resultid="3546" />
                    <RANKING order="14" place="14" resultid="5207" />
                    <RANKING order="15" place="15" resultid="4700" />
                    <RANKING order="16" place="16" resultid="4428" />
                    <RANKING order="17" place="17" resultid="2960" />
                    <RANKING order="18" place="18" resultid="1976" />
                    <RANKING order="19" place="19" resultid="3403" />
                    <RANKING order="20" place="20" resultid="5740" />
                    <RANKING order="21" place="21" resultid="6027" />
                    <RANKING order="22" place="22" resultid="2233" />
                    <RANKING order="23" place="-1" resultid="2114" />
                    <RANKING order="24" place="-1" resultid="5492" />
                    <RANKING order="25" place="-1" resultid="5699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5122" />
                    <RANKING order="2" place="2" resultid="6191" />
                    <RANKING order="3" place="3" resultid="2853" />
                    <RANKING order="4" place="4" resultid="3635" />
                    <RANKING order="5" place="4" resultid="5883" />
                    <RANKING order="6" place="6" resultid="3014" />
                    <RANKING order="7" place="7" resultid="3866" />
                    <RANKING order="8" place="8" resultid="3392" />
                    <RANKING order="9" place="9" resultid="4491" />
                    <RANKING order="10" place="10" resultid="5705" />
                    <RANKING order="11" place="11" resultid="2167" />
                    <RANKING order="12" place="12" resultid="2366" />
                    <RANKING order="13" place="13" resultid="3091" />
                    <RANKING order="14" place="14" resultid="5376" />
                    <RANKING order="15" place="15" resultid="6397" />
                    <RANKING order="16" place="16" resultid="3915" />
                    <RANKING order="17" place="17" resultid="5272" />
                    <RANKING order="18" place="18" resultid="3764" />
                    <RANKING order="19" place="-1" resultid="2173" />
                    <RANKING order="20" place="-1" resultid="2184" />
                    <RANKING order="21" place="-1" resultid="3264" />
                    <RANKING order="22" place="-1" resultid="3477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5291" />
                    <RANKING order="2" place="2" resultid="3254" />
                    <RANKING order="3" place="3" resultid="2542" />
                    <RANKING order="4" place="4" resultid="4469" />
                    <RANKING order="5" place="5" resultid="4657" />
                    <RANKING order="6" place="6" resultid="3829" />
                    <RANKING order="7" place="7" resultid="3343" />
                    <RANKING order="8" place="8" resultid="2351" />
                    <RANKING order="9" place="9" resultid="2247" />
                    <RANKING order="10" place="10" resultid="2826" />
                    <RANKING order="11" place="11" resultid="2161" />
                    <RANKING order="12" place="12" resultid="3179" />
                    <RANKING order="13" place="13" resultid="3359" />
                    <RANKING order="14" place="14" resultid="3169" />
                    <RANKING order="15" place="15" resultid="1884" />
                    <RANKING order="16" place="16" resultid="4722" />
                    <RANKING order="17" place="17" resultid="2194" />
                    <RANKING order="18" place="18" resultid="5265" />
                    <RANKING order="19" place="19" resultid="5286" />
                    <RANKING order="20" place="20" resultid="5316" />
                    <RANKING order="21" place="21" resultid="3259" />
                    <RANKING order="22" place="-1" resultid="2710" />
                    <RANKING order="23" place="-1" resultid="3647" />
                    <RANKING order="24" place="-1" resultid="4536" />
                    <RANKING order="25" place="-1" resultid="4443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5182" />
                    <RANKING order="2" place="2" resultid="5947" />
                    <RANKING order="3" place="3" resultid="1863" />
                    <RANKING order="4" place="4" resultid="3621" />
                    <RANKING order="5" place="5" resultid="4483" />
                    <RANKING order="6" place="6" resultid="4461" />
                    <RANKING order="7" place="7" resultid="6284" />
                    <RANKING order="8" place="8" resultid="2150" />
                    <RANKING order="9" place="9" resultid="3421" />
                    <RANKING order="10" place="10" resultid="3314" />
                    <RANKING order="11" place="11" resultid="5195" />
                    <RANKING order="12" place="12" resultid="3195" />
                    <RANKING order="13" place="-1" resultid="5041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3511" />
                    <RANKING order="2" place="2" resultid="4300" />
                    <RANKING order="3" place="3" resultid="5646" />
                    <RANKING order="4" place="4" resultid="4609" />
                    <RANKING order="5" place="5" resultid="3406" />
                    <RANKING order="6" place="6" resultid="2808" />
                    <RANKING order="7" place="7" resultid="2650" />
                    <RANKING order="8" place="8" resultid="4976" />
                    <RANKING order="9" place="9" resultid="5535" />
                    <RANKING order="10" place="10" resultid="2144" />
                    <RANKING order="11" place="11" resultid="2046" />
                    <RANKING order="12" place="12" resultid="4541" />
                    <RANKING order="13" place="13" resultid="4447" />
                    <RANKING order="14" place="14" resultid="4688" />
                    <RANKING order="15" place="-1" resultid="1984" />
                    <RANKING order="16" place="-1" resultid="2668" />
                    <RANKING order="17" place="-1" resultid="5865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2705" />
                    <RANKING order="2" place="2" resultid="2237" />
                    <RANKING order="3" place="3" resultid="3811" />
                    <RANKING order="4" place="4" resultid="5022" />
                    <RANKING order="5" place="5" resultid="4347" />
                    <RANKING order="6" place="6" resultid="2404" />
                    <RANKING order="7" place="7" resultid="2197" />
                    <RANKING order="8" place="8" resultid="6443" />
                    <RANKING order="9" place="9" resultid="4359" />
                    <RANKING order="10" place="10" resultid="4502" />
                    <RANKING order="11" place="11" resultid="3799" />
                    <RANKING order="12" place="12" resultid="4507" />
                    <RANKING order="13" place="13" resultid="3300" />
                    <RANKING order="14" place="14" resultid="6246" />
                    <RANKING order="15" place="15" resultid="3969" />
                    <RANKING order="16" place="16" resultid="3149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6251" />
                    <RANKING order="2" place="2" resultid="4312" />
                    <RANKING order="3" place="3" resultid="4568" />
                    <RANKING order="4" place="4" resultid="4436" />
                    <RANKING order="5" place="5" resultid="3551" />
                    <RANKING order="6" place="6" resultid="3791" />
                    <RANKING order="7" place="-1" resultid="6232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4452" />
                    <RANKING order="2" place="2" resultid="5325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2613" />
                    <RANKING order="2" place="2" resultid="2660" />
                    <RANKING order="3" place="3" resultid="3310" />
                    <RANKING order="4" place="4" resultid="2360" />
                    <RANKING order="5" place="5" resultid="1954" />
                    <RANKING order="6" place="-1" resultid="4493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7684" daytime="16:19" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7685" daytime="16:23" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7686" daytime="16:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7687" daytime="16:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7688" daytime="16:27" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7689" daytime="16:29" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7690" daytime="16:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7691" daytime="16:31" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7692" daytime="16:33" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7693" daytime="16:34" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7694" daytime="16:35" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7695" daytime="16:36" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7696" daytime="16:38" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7697" daytime="16:39" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7698" daytime="16:40" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7699" daytime="16:41" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7700" daytime="16:43" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7701" daytime="16:44" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7702" daytime="16:45" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7703" daytime="16:46" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="7704" daytime="16:48" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="7705" daytime="16:49" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="7706" daytime="16:50" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="7707" daytime="16:51" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="7708" daytime="16:53" number="25" order="25" status="OFFICIAL" />
                <HEAT heatid="7709" daytime="16:54" number="26" order="26" status="OFFICIAL" />
                <HEAT heatid="7710" daytime="16:55" number="27" order="27" status="OFFICIAL" />
                <HEAT heatid="7711" daytime="16:56" number="28" order="28" status="OFFICIAL" />
                <HEAT heatid="7712" daytime="16:57" number="29" order="29" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="16:59" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2568" />
                    <RANKING order="2" place="2" resultid="3955" />
                    <RANKING order="3" place="3" resultid="1968" />
                    <RANKING order="4" place="4" resultid="2213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3842" />
                    <RANKING order="2" place="2" resultid="4730" />
                    <RANKING order="3" place="3" resultid="6020" />
                    <RANKING order="4" place="4" resultid="3072" />
                    <RANKING order="5" place="-1" resultid="3804" />
                    <RANKING order="6" place="-1" resultid="4793" />
                    <RANKING order="7" place="-1" resultid="5567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5583" />
                    <RANKING order="2" place="2" resultid="5099" />
                    <RANKING order="3" place="3" resultid="3590" />
                    <RANKING order="4" place="4" resultid="4739" />
                    <RANKING order="5" place="5" resultid="6462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1940" />
                    <RANKING order="2" place="2" resultid="3383" />
                    <RANKING order="3" place="3" resultid="3616" />
                    <RANKING order="4" place="4" resultid="4019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5030" />
                    <RANKING order="2" place="2" resultid="4304" />
                    <RANKING order="3" place="-1" resultid="6099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5170" />
                    <RANKING order="2" place="2" resultid="3879" />
                    <RANKING order="3" place="3" resultid="2845" />
                    <RANKING order="4" place="4" resultid="4651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3036" />
                    <RANKING order="2" place="2" resultid="2136" />
                    <RANKING order="3" place="3" resultid="3933" />
                    <RANKING order="4" place="4" resultid="2263" />
                    <RANKING order="5" place="5" resultid="4553" />
                    <RANKING order="6" place="6" resultid="3131" />
                    <RANKING order="7" place="7" resultid="4625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2128" />
                    <RANKING order="2" place="2" resultid="4601" />
                    <RANKING order="3" place="3" resultid="2254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4269" />
                    <RANKING order="2" place="2" resultid="5257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1105" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1106" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1107" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7713" daytime="16:59" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7714" daytime="17:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7715" daytime="17:11" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7716" daytime="17:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7717" daytime="17:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7718" daytime="17:24" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1108" daytime="17:28" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1109" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3562" />
                    <RANKING order="2" place="2" resultid="5155" />
                    <RANKING order="3" place="3" resultid="6406" />
                    <RANKING order="4" place="4" resultid="2295" />
                    <RANKING order="5" place="5" resultid="2578" />
                    <RANKING order="6" place="6" resultid="2206" />
                    <RANKING order="7" place="7" resultid="3659" />
                    <RANKING order="8" place="-1" resultid="3532" />
                    <RANKING order="9" place="-1" resultid="6211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2021" />
                    <RANKING order="2" place="2" resultid="5141" />
                    <RANKING order="3" place="3" resultid="5824" />
                    <RANKING order="4" place="4" resultid="6275" />
                    <RANKING order="5" place="5" resultid="2052" />
                    <RANKING order="6" place="6" resultid="5807" />
                    <RANKING order="7" place="7" resultid="4775" />
                    <RANKING order="8" place="8" resultid="3735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5600" />
                    <RANKING order="2" place="2" resultid="2067" />
                    <RANKING order="3" place="3" resultid="5962" />
                    <RANKING order="4" place="4" resultid="4800" />
                    <RANKING order="5" place="5" resultid="5629" />
                    <RANKING order="6" place="6" resultid="3518" />
                    <RANKING order="7" place="7" resultid="3062" />
                    <RANKING order="8" place="8" resultid="5588" />
                    <RANKING order="9" place="9" resultid="4163" />
                    <RANKING order="10" place="10" resultid="4715" />
                    <RANKING order="11" place="11" resultid="5241" />
                    <RANKING order="12" place="12" resultid="4213" />
                    <RANKING order="13" place="-1" resultid="5774" />
                    <RANKING order="14" place="-1" resultid="4153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2308" />
                    <RANKING order="2" place="2" resultid="1899" />
                    <RANKING order="3" place="3" resultid="2861" />
                    <RANKING order="4" place="4" resultid="2783" />
                    <RANKING order="5" place="5" resultid="6049" />
                    <RANKING order="6" place="6" resultid="5916" />
                    <RANKING order="7" place="7" resultid="5201" />
                    <RANKING order="8" place="8" resultid="2836" />
                    <RANKING order="9" place="9" resultid="4207" />
                    <RANKING order="10" place="10" resultid="2869" />
                    <RANKING order="11" place="11" resultid="1913" />
                    <RANKING order="12" place="-1" resultid="1946" />
                    <RANKING order="13" place="-1" resultid="4763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2791" />
                    <RANKING order="2" place="2" resultid="5415" />
                    <RANKING order="3" place="3" resultid="6173" />
                    <RANKING order="4" place="4" resultid="3603" />
                    <RANKING order="5" place="5" resultid="5208" />
                    <RANKING order="6" place="6" resultid="2088" />
                    <RANKING order="7" place="7" resultid="4319" />
                    <RANKING order="8" place="8" resultid="5216" />
                    <RANKING order="9" place="9" resultid="2727" />
                    <RANKING order="10" place="10" resultid="3464" />
                    <RANKING order="11" place="11" resultid="5741" />
                    <RANKING order="12" place="-1" resultid="3361" />
                    <RANKING order="13" place="-1" resultid="4329" />
                    <RANKING order="14" place="-1" resultid="4590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3654" />
                    <RANKING order="2" place="2" resultid="6192" />
                    <RANKING order="3" place="3" resultid="6057" />
                    <RANKING order="4" place="4" resultid="5528" />
                    <RANKING order="5" place="5" resultid="5706" />
                    <RANKING order="6" place="6" resultid="3092" />
                    <RANKING order="7" place="7" resultid="6398" />
                    <RANKING order="8" place="8" resultid="3719" />
                    <RANKING order="9" place="-1" resultid="3478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4035" />
                    <RANKING order="2" place="2" resultid="2543" />
                    <RANKING order="3" place="3" resultid="2827" />
                    <RANKING order="4" place="4" resultid="3224" />
                    <RANKING order="5" place="5" resultid="2248" />
                    <RANKING order="6" place="6" resultid="3180" />
                    <RANKING order="7" place="7" resultid="3768" />
                    <RANKING order="8" place="8" resultid="2156" />
                    <RANKING order="9" place="9" resultid="5317" />
                    <RANKING order="10" place="-1" resultid="2689" />
                    <RANKING order="11" place="-1" resultid="5016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6005" />
                    <RANKING order="2" place="2" resultid="5042" />
                    <RANKING order="3" place="3" resultid="2552" />
                    <RANKING order="4" place="4" resultid="2622" />
                    <RANKING order="5" place="5" resultid="4134" />
                    <RANKING order="6" place="6" resultid="5637" />
                    <RANKING order="7" place="7" resultid="5520" />
                    <RANKING order="8" place="8" resultid="4484" />
                    <RANKING order="9" place="9" resultid="3201" />
                    <RANKING order="10" place="-1" resultid="3173" />
                    <RANKING order="11" place="-1" resultid="3045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4420" />
                    <RANKING order="2" place="2" resultid="5647" />
                    <RANKING order="3" place="3" resultid="6182" />
                    <RANKING order="4" place="4" resultid="2809" />
                    <RANKING order="5" place="5" resultid="3407" />
                    <RANKING order="6" place="6" resultid="3446" />
                    <RANKING order="7" place="7" resultid="4582" />
                    <RANKING order="8" place="8" resultid="5654" />
                    <RANKING order="9" place="9" resultid="3455" />
                    <RANKING order="10" place="-1" resultid="4977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2684" />
                    <RANKING order="2" place="2" resultid="2238" />
                    <RANKING order="3" place="3" resultid="5506" />
                    <RANKING order="4" place="4" resultid="2736" />
                    <RANKING order="5" place="5" resultid="3290" />
                    <RANKING order="6" place="6" resultid="4503" />
                    <RANKING order="7" place="7" resultid="3301" />
                    <RANKING order="8" place="-1" resultid="6247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4295" />
                    <RANKING order="2" place="2" resultid="4569" />
                    <RANKING order="3" place="3" resultid="6233" />
                    <RANKING order="4" place="-1" resultid="3792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4453" />
                    <RANKING order="2" place="2" resultid="5249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1123" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7719" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7720" daytime="17:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7721" daytime="17:39" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7722" daytime="17:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7723" daytime="17:49" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7724" daytime="17:53" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7725" daytime="17:57" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7726" daytime="18:01" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7727" daytime="18:05" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7728" daytime="18:08" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7729" daytime="18:12" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7730" daytime="18:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7731" daytime="18:19" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7732" daytime="18:22" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7733" daytime="18:25" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="18:29" gender="X" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="96" agemin="80" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="1126" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4114" />
                    <RANKING order="2" place="2" resultid="4808" />
                    <RANKING order="3" place="3" resultid="6450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4806" />
                    <RANKING order="2" place="2" resultid="3976" />
                    <RANKING order="3" place="3" resultid="2998" />
                    <RANKING order="4" place="4" resultid="3084" />
                    <RANKING order="5" place="5" resultid="3502" />
                    <RANKING order="6" place="6" resultid="3706" />
                    <RANKING order="7" place="-1" resultid="5661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3975" />
                    <RANKING order="2" place="2" resultid="4115" />
                    <RANKING order="3" place="3" resultid="2999" />
                    <RANKING order="4" place="4" resultid="6083" />
                    <RANKING order="5" place="5" resultid="6451" />
                    <RANKING order="6" place="6" resultid="4711" />
                    <RANKING order="7" place="-1" resultid="5797" />
                    <RANKING order="8" place="-1" resultid="3083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5048" />
                    <RANKING order="2" place="2" resultid="2188" />
                    <RANKING order="3" place="3" resultid="3978" />
                    <RANKING order="4" place="4" resultid="5049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4379" />
                    <RANKING order="2" place="2" resultid="3980" />
                    <RANKING order="3" place="3" resultid="4632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="400" agemin="280" name="Kategoria F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4378" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7734" daytime="18:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7735" daytime="18:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7736" daytime="18:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7737" daytime="18:38" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="18:41" gender="F" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3907" />
                    <RANKING order="2" place="2" resultid="3956" />
                    <RANKING order="3" place="3" resultid="5575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4048" />
                    <RANKING order="2" place="2" resultid="4409" />
                    <RANKING order="3" place="3" resultid="3073" />
                    <RANKING order="4" place="4" resultid="5308" />
                    <RANKING order="5" place="5" resultid="3078" />
                    <RANKING order="6" place="6" resultid="3126" />
                    <RANKING order="7" place="-1" resultid="4794" />
                    <RANKING order="8" place="-1" resultid="6309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2272" />
                    <RANKING order="2" place="2" resultid="4787" />
                    <RANKING order="3" place="3" resultid="5873" />
                    <RANKING order="4" place="4" resultid="4027" />
                    <RANKING order="5" place="5" resultid="6013" />
                    <RANKING order="6" place="-1" resultid="5783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3693" />
                    <RANKING order="2" place="2" resultid="3859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="44" agemin="40" name="Kategoria D" />
                <AGEGROUP agegroupid="1146" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3104" />
                    <RANKING order="2" place="2" resultid="6070" />
                    <RANKING order="3" place="3" resultid="4146" />
                    <RANKING order="4" place="4" resultid="3216" />
                    <RANKING order="5" place="5" resultid="3613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3037" />
                    <RANKING order="2" place="2" resultid="4681" />
                    <RANKING order="3" place="3" resultid="3934" />
                    <RANKING order="4" place="4" resultid="4554" />
                    <RANKING order="5" place="5" resultid="4562" />
                    <RANKING order="6" place="6" resultid="3132" />
                    <RANKING order="7" place="7" resultid="6108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3925" />
                    <RANKING order="2" place="-1" resultid="6141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1149" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5004" />
                    <RANKING order="2" place="2" resultid="5388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="1151" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4270" />
                    <RANKING order="2" place="-1" resultid="3432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1153" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1155" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8712" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8713" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8714" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8715" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8716" number="5" order="5" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1729" />
                <TIMESTANDARDREF timestandardlistid="1739" />
                <TIMESTANDARDREF timestandardlistid="1743" />
                <TIMESTANDARDREF timestandardlistid="1747" />
                <TIMESTANDARDREF timestandardlistid="1751" />
                <TIMESTANDARDREF timestandardlistid="1755" />
                <TIMESTANDARDREF timestandardlistid="1759" />
                <TIMESTANDARDREF timestandardlistid="1763" />
                <TIMESTANDARDREF timestandardlistid="1767" />
                <TIMESTANDARDREF timestandardlistid="1775" />
                <TIMESTANDARDREF timestandardlistid="1771" />
                <TIMESTANDARDREF timestandardlistid="1779" />
                <TIMESTANDARDREF timestandardlistid="1783" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1156" daytime="20:05" gender="M" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1157" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5953" />
                    <RANKING order="2" place="2" resultid="3896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3241" />
                    <RANKING order="2" place="2" resultid="4801" />
                    <RANKING order="3" place="3" resultid="4227" />
                    <RANKING order="4" place="4" resultid="3586" />
                    <RANKING order="5" place="5" resultid="3739" />
                    <RANKING order="6" place="-1" resultid="4154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5555" />
                    <RANKING order="2" place="2" resultid="3110" />
                    <RANKING order="3" place="3" resultid="3757" />
                    <RANKING order="4" place="4" resultid="4208" />
                    <RANKING order="5" place="5" resultid="5917" />
                    <RANKING order="6" place="6" resultid="3054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6174" />
                    <RANKING order="2" place="2" resultid="3854" />
                    <RANKING order="3" place="3" resultid="5189" />
                    <RANKING order="4" place="4" resultid="2774" />
                    <RANKING order="5" place="5" resultid="6187" />
                    <RANKING order="6" place="6" resultid="2004" />
                    <RANKING order="7" place="7" resultid="6378" />
                    <RANKING order="8" place="8" resultid="6311" />
                    <RANKING order="9" place="9" resultid="3465" />
                    <RANKING order="10" place="10" resultid="3471" />
                    <RANKING order="11" place="11" resultid="5095" />
                    <RANKING order="12" place="12" resultid="2979" />
                    <RANKING order="13" place="13" resultid="4747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2180" />
                    <RANKING order="2" place="2" resultid="5884" />
                    <RANKING order="3" place="3" resultid="2347" />
                    <RANKING order="4" place="4" resultid="2694" />
                    <RANKING order="5" place="5" resultid="2038" />
                    <RANKING order="6" place="6" resultid="3231" />
                    <RANKING order="7" place="7" resultid="3015" />
                    <RANKING order="8" place="8" resultid="6058" />
                    <RANKING order="9" place="9" resultid="3724" />
                    <RANKING order="10" place="10" resultid="3916" />
                    <RANKING order="11" place="11" resultid="3720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5496" />
                    <RANKING order="2" place="2" resultid="3648" />
                    <RANKING order="3" place="3" resultid="2602" />
                    <RANKING order="4" place="4" resultid="3769" />
                    <RANKING order="5" place="5" resultid="3210" />
                    <RANKING order="6" place="6" resultid="2195" />
                    <RANKING order="7" place="7" resultid="4723" />
                    <RANKING order="8" place="-1" resultid="5287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3608" />
                    <RANKING order="2" place="2" resultid="2639" />
                    <RANKING order="3" place="3" resultid="6285" />
                    <RANKING order="4" place="4" resultid="5423" />
                    <RANKING order="5" place="5" resultid="6118" />
                    <RANKING order="6" place="6" resultid="5196" />
                    <RANKING order="7" place="-1" resultid="1864" />
                    <RANKING order="8" place="-1" resultid="4462" />
                    <RANKING order="9" place="-1" resultid="3046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4610" />
                    <RANKING order="2" place="2" resultid="3447" />
                    <RANKING order="3" place="3" resultid="2651" />
                    <RANKING order="4" place="4" resultid="2669" />
                    <RANKING order="5" place="5" resultid="5514" />
                    <RANKING order="6" place="6" resultid="3456" />
                    <RANKING order="7" place="-1" resultid="1985" />
                    <RANKING order="8" place="-1" resultid="3630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3812" />
                    <RANKING order="2" place="2" resultid="2198" />
                    <RANKING order="3" place="3" resultid="2405" />
                    <RANKING order="4" place="-1" resultid="3291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3552" />
                    <RANKING order="2" place="2" resultid="3893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5164" />
                    <RANKING order="2" place="-1" resultid="1955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1171" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8717" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8718" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8719" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8720" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8721" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8722" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8723" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8724" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8725" number="9" order="9" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1785" />
                <TIMESTANDARDREF timestandardlistid="1789" />
                <TIMESTANDARDREF timestandardlistid="1793" />
                <TIMESTANDARDREF timestandardlistid="1797" />
                <TIMESTANDARDREF timestandardlistid="1801" />
                <TIMESTANDARDREF timestandardlistid="1805" />
                <TIMESTANDARDREF timestandardlistid="1809" />
                <TIMESTANDARDREF timestandardlistid="1813" />
                <TIMESTANDARDREF timestandardlistid="1817" />
                <TIMESTANDARDREF timestandardlistid="1821" />
                <TIMESTANDARDREF timestandardlistid="1825" />
                <TIMESTANDARDREF timestandardlistid="1829" />
                <TIMESTANDARDREF timestandardlistid="1833" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="8925" />
            <JUDGE officialid="8910" />
            <JUDGE officialid="8924" />
            <JUDGE officialid="8926" />
            <JUDGE officialid="8906" />
            <JUDGE officialid="8919" />
            <JUDGE officialid="8923" />
            <JUDGE officialid="8909" />
            <JUDGE officialid="8921" />
            <JUDGE officialid="8914" />
            <JUDGE officialid="8915" />
            <JUDGE officialid="8918" />
            <JUDGE officialid="8922" />
            <JUDGE officialid="8917" />
            <JUDGE officialid="8920" />
            <JUDGE officialid="8928" />
            <JUDGE officialid="8912" />
            <JUDGE officialid="8916" />
            <JUDGE officialid="8916" />
            <JUDGE officialid="8908" />
            <JUDGE officialid="8908" />
            <JUDGE officialid="8911" />
            <JUDGE officialid="8911" />
            <JUDGE officialid="8913" />
            <JUDGE officialid="8927" />
            <JUDGE officialid="8905" />
            <JUDGE officialid="8904" />
            <JUDGE officialid="8903" />
            <JUDGE officialid="8907" />
            <JUDGE officialid="8941" />
            <JUDGE officialid="8901" />
            <JUDGE officialid="8902" />
          </JUDGES>
        </SESSION>
        <SESSION date="2013-11-16" daytime="09:00" name="MP Masters BLOK II" number="2" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1173" daytime="09:00" gender="F" number="8" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1175" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6199" />
                    <RANKING order="2" place="2" resultid="2628" />
                    <RANKING order="3" place="3" resultid="5150" />
                    <RANKING order="4" place="4" resultid="3903" />
                    <RANKING order="5" place="5" resultid="2062" />
                    <RANKING order="6" place="6" resultid="3029" />
                    <RANKING order="7" place="7" resultid="2214" />
                    <RANKING order="8" place="8" resultid="1987" />
                    <RANKING order="9" place="-1" resultid="2001" />
                    <RANKING order="10" place="-1" resultid="5839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3843" />
                    <RANKING order="2" place="2" resultid="6350" />
                    <RANKING order="3" place="3" resultid="4731" />
                    <RANKING order="4" place="4" resultid="6021" />
                    <RANKING order="5" place="5" resultid="6293" />
                    <RANKING order="6" place="-1" resultid="2922" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5584" />
                    <RANKING order="2" place="2" resultid="3591" />
                    <RANKING order="3" place="3" resultid="6032" />
                    <RANKING order="4" place="4" resultid="3494" />
                    <RANKING order="5" place="5" resultid="5929" />
                    <RANKING order="6" place="-1" resultid="3682" />
                    <RANKING order="7" place="-1" resultid="4788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2927" />
                    <RANKING order="2" place="2" resultid="2229" />
                    <RANKING order="3" place="3" resultid="6203" />
                    <RANKING order="4" place="4" resultid="5280" />
                    <RANKING order="5" place="5" resultid="4020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5036" />
                    <RANKING order="2" place="2" resultid="5493" />
                    <RANKING order="3" place="3" resultid="3889" />
                    <RANKING order="4" place="4" resultid="6458" />
                    <RANKING order="5" place="5" resultid="6382" />
                    <RANKING order="6" place="6" resultid="3641" />
                    <RANKING order="7" place="7" resultid="3747" />
                    <RANKING order="8" place="8" resultid="2947" />
                    <RANKING order="9" place="9" resultid="4695" />
                    <RANKING order="10" place="10" resultid="3872" />
                    <RANKING order="11" place="11" resultid="6305" />
                    <RANKING order="12" place="12" resultid="2377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4367" />
                    <RANKING order="2" place="2" resultid="5489" />
                    <RANKING order="3" place="3" resultid="6779" />
                    <RANKING order="4" place="4" resultid="3217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4986" />
                    <RANKING order="2" place="2" resultid="2137" />
                    <RANKING order="3" place="3" resultid="5177" />
                    <RANKING order="4" place="4" resultid="4563" />
                    <RANKING order="5" place="5" resultid="3417" />
                    <RANKING order="6" place="-1" resultid="4555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3397" />
                    <RANKING order="2" place="2" resultid="3926" />
                    <RANKING order="3" place="3" resultid="2007" />
                    <RANKING order="4" place="4" resultid="3141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4341" />
                    <RANKING order="2" place="2" resultid="6315" />
                    <RANKING order="3" place="3" resultid="3378" />
                    <RANKING order="4" place="4" resultid="3356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5771" />
                    <RANKING order="2" place="2" resultid="4672" />
                    <RANKING order="3" place="3" resultid="4054" />
                    <RANKING order="4" place="4" resultid="4355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4290" />
                    <RANKING order="2" place="2" resultid="6343" />
                    <RANKING order="3" place="3" resultid="5258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1187" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7753" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7754" daytime="09:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7755" daytime="09:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7756" daytime="09:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7757" daytime="09:07" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7758" daytime="09:09" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7759" daytime="09:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7760" daytime="09:12" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7761" daytime="09:13" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1190" daytime="09:15" gender="M" number="9" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1191" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3563" />
                    <RANKING order="2" place="2" resultid="6242" />
                    <RANKING order="3" place="3" resultid="5687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5954" />
                    <RANKING order="2" place="2" resultid="6139" />
                    <RANKING order="3" place="3" resultid="6276" />
                    <RANKING order="4" place="4" resultid="6326" />
                    <RANKING order="5" place="5" resultid="2587" />
                    <RANKING order="6" place="6" resultid="5402" />
                    <RANKING order="7" place="7" resultid="2075" />
                    <RANKING order="8" place="8" resultid="4512" />
                    <RANKING order="9" place="9" resultid="3427" />
                    <RANKING order="10" place="10" resultid="5115" />
                    <RANKING order="11" place="11" resultid="3688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4108" />
                    <RANKING order="2" place="2" resultid="3238" />
                    <RANKING order="3" place="3" resultid="5963" />
                    <RANKING order="4" place="4" resultid="4059" />
                    <RANKING order="5" place="5" resultid="4802" />
                    <RANKING order="6" place="6" resultid="3529" />
                    <RANKING order="7" place="7" resultid="4164" />
                    <RANKING order="8" place="8" resultid="4180" />
                    <RANKING order="9" place="9" resultid="4716" />
                    <RANKING order="10" place="10" resultid="4214" />
                    <RANKING order="11" place="-1" resultid="3740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1900" />
                    <RANKING order="2" place="2" resultid="2784" />
                    <RANKING order="3" place="3" resultid="6333" />
                    <RANKING order="4" place="4" resultid="6065" />
                    <RANKING order="5" place="5" resultid="1914" />
                    <RANKING order="6" place="6" resultid="2837" />
                    <RANKING order="7" place="7" resultid="2915" />
                    <RANKING order="8" place="8" resultid="3758" />
                    <RANKING order="9" place="9" resultid="2988" />
                    <RANKING order="10" place="10" resultid="3947" />
                    <RANKING order="11" place="11" resultid="4764" />
                    <RANKING order="12" place="12" resultid="3851" />
                    <RANKING order="13" place="-1" resultid="2396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5416" />
                    <RANKING order="2" place="2" resultid="4330" />
                    <RANKING order="3" place="3" resultid="4667" />
                    <RANKING order="4" place="4" resultid="3943" />
                    <RANKING order="5" place="5" resultid="2094" />
                    <RANKING order="6" place="6" resultid="3604" />
                    <RANKING order="7" place="7" resultid="5209" />
                    <RANKING order="8" place="8" resultid="6370" />
                    <RANKING order="9" place="9" resultid="3362" />
                    <RANKING order="10" place="10" resultid="5700" />
                    <RANKING order="11" place="11" resultid="4429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4373" />
                    <RANKING order="2" place="2" resultid="5345" />
                    <RANKING order="3" place="3" resultid="6337" />
                    <RANKING order="4" place="4" resultid="3232" />
                    <RANKING order="5" place="5" resultid="5885" />
                    <RANKING order="6" place="6" resultid="2854" />
                    <RANKING order="7" place="7" resultid="5707" />
                    <RANKING order="8" place="8" resultid="2039" />
                    <RANKING order="9" place="9" resultid="3721" />
                    <RANKING order="10" place="-1" resultid="2174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4036" />
                    <RANKING order="2" place="2" resultid="4470" />
                    <RANKING order="3" place="3" resultid="4658" />
                    <RANKING order="4" place="4" resultid="3344" />
                    <RANKING order="5" place="5" resultid="2690" />
                    <RANKING order="6" place="6" resultid="3830" />
                    <RANKING order="7" place="7" resultid="5477" />
                    <RANKING order="8" place="8" resultid="3181" />
                    <RANKING order="9" place="9" resultid="4336" />
                    <RANKING order="10" place="10" resultid="1885" />
                    <RANKING order="11" place="11" resultid="5266" />
                    <RANKING order="12" place="-1" resultid="2162" />
                    <RANKING order="13" place="-1" resultid="4444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5183" />
                    <RANKING order="2" place="2" resultid="3317" />
                    <RANKING order="3" place="3" resultid="5043" />
                    <RANKING order="4" place="4" resultid="2623" />
                    <RANKING order="5" place="5" resultid="4463" />
                    <RANKING order="6" place="6" resultid="2151" />
                    <RANKING order="7" place="7" resultid="5521" />
                    <RANKING order="8" place="8" resultid="3174" />
                    <RANKING order="9" place="9" resultid="5424" />
                    <RANKING order="10" place="10" resultid="3202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3512" />
                    <RANKING order="2" place="2" resultid="2652" />
                    <RANKING order="3" place="3" resultid="4978" />
                    <RANKING order="4" place="4" resultid="3448" />
                    <RANKING order="5" place="5" resultid="3408" />
                    <RANKING order="6" place="6" resultid="2810" />
                    <RANKING order="7" place="7" resultid="2670" />
                    <RANKING order="8" place="8" resultid="5515" />
                    <RANKING order="9" place="9" resultid="4448" />
                    <RANKING order="10" place="10" resultid="5608" />
                    <RANKING order="11" place="-1" resultid="2145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4281" />
                    <RANKING order="2" place="2" resultid="2680" />
                    <RANKING order="3" place="3" resultid="3439" />
                    <RANKING order="4" place="4" resultid="2723" />
                    <RANKING order="5" place="5" resultid="4348" />
                    <RANKING order="6" place="6" resultid="4508" />
                    <RANKING order="7" place="7" resultid="3292" />
                    <RANKING order="8" place="8" resultid="3800" />
                    <RANKING order="9" place="9" resultid="3413" />
                    <RANKING order="10" place="10" resultid="6444" />
                    <RANKING order="11" place="11" resultid="3150" />
                    <RANKING order="12" place="-1" resultid="6248" />
                    <RANKING order="13" place="-1" resultid="5615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4313" />
                    <RANKING order="2" place="2" resultid="4570" />
                    <RANKING order="3" place="3" resultid="3553" />
                    <RANKING order="4" place="4" resultid="4437" />
                    <RANKING order="5" place="5" resultid="5623" />
                    <RANKING order="6" place="-1" resultid="3793" />
                    <RANKING order="7" place="-1" resultid="6234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4454" />
                    <RANKING order="2" place="2" resultid="4577" />
                    <RANKING order="3" place="3" resultid="5970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2615" />
                    <RANKING order="2" place="2" resultid="2661" />
                    <RANKING order="3" place="3" resultid="2013" />
                    <RANKING order="4" place="4" resultid="1956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7762" daytime="09:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7763" daytime="09:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7764" daytime="09:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7765" daytime="09:21" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7766" daytime="09:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7767" daytime="09:24" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7768" daytime="09:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7769" daytime="09:27" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7770" daytime="09:28" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7771" daytime="09:30" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7772" daytime="09:31" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7773" daytime="09:32" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7774" daytime="09:34" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7775" daytime="09:35" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7776" daytime="09:36" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7777" daytime="09:38" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1206" daytime="09:39" gender="F" number="10" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1207" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5576" />
                    <RANKING order="2" place="2" resultid="5108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5568" />
                    <RANKING order="2" place="2" resultid="3960" />
                    <RANKING order="3" place="3" resultid="3805" />
                    <RANKING order="4" place="4" resultid="1963" />
                    <RANKING order="5" place="5" resultid="5234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4042" />
                    <RANKING order="2" place="2" resultid="5100" />
                    <RANKING order="3" place="3" resultid="4740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5408" />
                    <RANKING order="2" place="2" resultid="5130" />
                    <RANKING order="3" place="3" resultid="3617" />
                    <RANKING order="4" place="4" resultid="3487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4305" />
                    <RANKING order="2" place="2" resultid="6127" />
                    <RANKING order="3" place="3" resultid="5880" />
                    <RANKING order="4" place="4" resultid="3068" />
                    <RANKING order="5" place="5" resultid="3873" />
                    <RANKING order="6" place="-1" resultid="6100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5171" />
                    <RANKING order="2" place="2" resultid="5371" />
                    <RANKING order="3" place="3" resultid="6071" />
                    <RANKING order="4" place="4" resultid="2846" />
                    <RANKING order="5" place="5" resultid="6466" />
                    <RANKING order="6" place="6" resultid="2370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3884" />
                    <RANKING order="2" place="2" resultid="6363" />
                    <RANKING order="3" place="3" resultid="5936" />
                    <RANKING order="4" place="4" resultid="4682" />
                    <RANKING order="5" place="5" resultid="3571" />
                    <RANKING order="6" place="6" resultid="2264" />
                    <RANKING order="7" place="7" resultid="4626" />
                    <RANKING order="8" place="8" resultid="3161" />
                    <RANKING order="9" place="9" resultid="2761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4602" />
                    <RANKING order="2" place="2" resultid="2255" />
                    <RANKING order="3" place="3" resultid="2530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6168" />
                    <RANKING order="2" place="2" resultid="3786" />
                    <RANKING order="3" place="3" resultid="5078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4271" />
                    <RANKING order="2" place="-1" resultid="6344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3116" />
                    <RANKING order="2" place="-1" resultid="2122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1220" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1221" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7778" daytime="09:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7779" daytime="09:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7780" daytime="09:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7781" daytime="09:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7782" daytime="10:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7783" daytime="10:04" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1222" daytime="10:09" gender="M" number="11" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1223" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5157" />
                    <RANKING order="2" place="2" resultid="2207" />
                    <RANKING order="3" place="3" resultid="2560" />
                    <RANKING order="4" place="4" resultid="5688" />
                    <RANKING order="5" place="-1" resultid="2287" />
                    <RANKING order="6" place="-1" resultid="3533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5816" />
                    <RANKING order="2" place="2" resultid="5381" />
                    <RANKING order="3" place="3" resultid="2022" />
                    <RANKING order="4" place="4" resultid="5808" />
                    <RANKING order="5" place="5" resultid="5351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4085" />
                    <RANKING order="2" place="2" resultid="5601" />
                    <RANKING order="3" place="3" resultid="6043" />
                    <RANKING order="4" place="4" resultid="4186" />
                    <RANKING order="5" place="5" resultid="5630" />
                    <RANKING order="6" place="6" resultid="4155" />
                    <RANKING order="7" place="7" resultid="2330" />
                    <RANKING order="8" place="8" resultid="4165" />
                    <RANKING order="9" place="-1" resultid="5595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2862" />
                    <RANKING order="2" place="2" resultid="2878" />
                    <RANKING order="3" place="3" resultid="3349" />
                    <RANKING order="4" place="4" resultid="2870" />
                    <RANKING order="5" place="5" resultid="2321" />
                    <RANKING order="6" place="6" resultid="3055" />
                    <RANKING order="7" place="7" resultid="5912" />
                    <RANKING order="8" place="8" resultid="5925" />
                    <RANKING order="9" place="-1" resultid="4782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3664" />
                    <RANKING order="2" place="2" resultid="2714" />
                    <RANKING order="3" place="3" resultid="6357" />
                    <RANKING order="4" place="4" resultid="2729" />
                    <RANKING order="5" place="5" resultid="2980" />
                    <RANKING order="6" place="6" resultid="3472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5123" />
                    <RANKING order="2" place="2" resultid="3016" />
                    <RANKING order="3" place="3" resultid="5529" />
                    <RANKING order="4" place="4" resultid="2168" />
                    <RANKING order="5" place="5" resultid="5377" />
                    <RANKING order="6" place="6" resultid="5273" />
                    <RANKING order="7" place="7" resultid="3917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4659" />
                    <RANKING order="2" place="2" resultid="3225" />
                    <RANKING order="3" place="3" resultid="5892" />
                    <RANKING order="4" place="4" resultid="2249" />
                    <RANKING order="5" place="5" resultid="2157" />
                    <RANKING order="6" place="6" resultid="3770" />
                    <RANKING order="7" place="7" resultid="5012" />
                    <RANKING order="8" place="8" resultid="5318" />
                    <RANKING order="9" place="9" resultid="3260" />
                    <RANKING order="10" place="-1" resultid="5017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4958" />
                    <RANKING order="2" place="2" resultid="4135" />
                    <RANKING order="3" place="3" resultid="2553" />
                    <RANKING order="4" place="4" resultid="4498" />
                    <RANKING order="5" place="5" resultid="3626" />
                    <RANKING order="6" place="6" resultid="3203" />
                    <RANKING order="7" place="7" resultid="6119" />
                    <RANKING order="8" place="8" resultid="2751" />
                    <RANKING order="9" place="9" resultid="3196" />
                    <RANKING order="10" place="10" resultid="4090" />
                    <RANKING order="11" place="-1" resultid="2536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4421" />
                    <RANKING order="2" place="2" resultid="4476" />
                    <RANKING order="3" place="3" resultid="6183" />
                    <RANKING order="4" place="4" resultid="5642" />
                    <RANKING order="5" place="5" resultid="4611" />
                    <RANKING order="6" place="6" resultid="4583" />
                    <RANKING order="7" place="7" resultid="3188" />
                    <RANKING order="8" place="8" resultid="3457" />
                    <RANKING order="9" place="9" resultid="5655" />
                    <RANKING order="10" place="-1" resultid="3631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4999" />
                    <RANKING order="2" place="2" resultid="2685" />
                    <RANKING order="3" place="3" resultid="5507" />
                    <RANKING order="4" place="4" resultid="3302" />
                    <RANKING order="5" place="5" resultid="3151" />
                    <RANKING order="6" place="-1" resultid="5616" />
                    <RANKING order="7" place="-1" resultid="3970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4276" />
                    <RANKING order="2" place="2" resultid="2744" />
                    <RANKING order="3" place="3" resultid="4438" />
                    <RANKING order="4" place="4" resultid="4571" />
                    <RANKING order="5" place="5" resultid="1997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4578" />
                    <RANKING order="2" place="2" resultid="5250" />
                    <RANKING order="3" place="3" resultid="5971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2662" />
                    <RANKING order="2" place="2" resultid="2361" />
                    <RANKING order="3" place="3" resultid="5165" />
                    <RANKING order="4" place="4" resultid="4494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1237" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7784" daytime="10:09" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7785" daytime="10:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7786" daytime="10:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7787" daytime="10:27" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7788" daytime="10:31" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7789" daytime="10:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7790" daytime="10:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7791" daytime="10:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7792" daytime="10:48" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7793" daytime="10:52" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7794" daytime="10:56" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7795" daytime="11:00" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1238" daytime="11:04" gender="F" number="12" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1239" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2570" />
                    <RANKING order="2" place="2" resultid="5151" />
                    <RANKING order="3" place="3" resultid="2607" />
                    <RANKING order="4" place="4" resultid="1969" />
                    <RANKING order="5" place="5" resultid="3778" />
                    <RANKING order="6" place="6" resultid="3908" />
                    <RANKING order="7" place="7" resultid="5840" />
                    <RANKING order="8" place="8" resultid="2995" />
                    <RANKING order="9" place="9" resultid="3904" />
                    <RANKING order="10" place="10" resultid="5109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4049" />
                    <RANKING order="2" place="2" resultid="6351" />
                    <RANKING order="3" place="3" resultid="3541" />
                    <RANKING order="4" place="4" resultid="4410" />
                    <RANKING order="5" place="5" resultid="2335" />
                    <RANKING order="6" place="6" resultid="5309" />
                    <RANKING order="7" place="7" resultid="2584" />
                    <RANKING order="8" place="8" resultid="5361" />
                    <RANKING order="9" place="9" resultid="3127" />
                    <RANKING order="10" place="-1" resultid="5792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5442" />
                    <RANKING order="2" place="2" resultid="5874" />
                    <RANKING order="3" place="3" resultid="2273" />
                    <RANKING order="4" place="4" resultid="4028" />
                    <RANKING order="5" place="5" resultid="6014" />
                    <RANKING order="6" place="6" resultid="2298" />
                    <RANKING order="7" place="7" resultid="3495" />
                    <RANKING order="8" place="8" resultid="3683" />
                    <RANKING order="9" place="-1" resultid="4097" />
                    <RANKING order="10" place="-1" resultid="4789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2935" />
                    <RANKING order="2" place="2" resultid="2942" />
                    <RANKING order="3" place="3" resultid="3694" />
                    <RANKING order="4" place="4" resultid="2230" />
                    <RANKING order="5" place="5" resultid="2957" />
                    <RANKING order="6" place="6" resultid="5899" />
                    <RANKING order="7" place="7" resultid="5281" />
                    <RANKING order="8" place="8" resultid="3488" />
                    <RANKING order="9" place="9" resultid="3860" />
                    <RANKING order="10" place="-1" resultid="5764" />
                    <RANKING order="11" place="-1" resultid="6693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4306" />
                    <RANKING order="2" place="2" resultid="6383" />
                    <RANKING order="3" place="3" resultid="6459" />
                    <RANKING order="4" place="4" resultid="3525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3105" />
                    <RANKING order="2" place="2" resultid="6321" />
                    <RANKING order="3" place="3" resultid="3713" />
                    <RANKING order="4" place="4" resultid="4652" />
                    <RANKING order="5" place="5" resultid="3218" />
                    <RANKING order="6" place="6" resultid="2372" />
                    <RANKING order="7" place="-1" resultid="4147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4993" />
                    <RANKING order="2" place="2" resultid="6404" />
                    <RANKING order="3" place="3" resultid="5178" />
                    <RANKING order="4" place="4" resultid="3935" />
                    <RANKING order="5" place="5" resultid="4618" />
                    <RANKING order="6" place="6" resultid="4564" />
                    <RANKING order="7" place="7" resultid="3133" />
                    <RANKING order="8" place="8" resultid="3572" />
                    <RANKING order="9" place="9" resultid="3162" />
                    <RANKING order="10" place="10" resultid="2762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3730" />
                    <RANKING order="2" place="2" resultid="1980" />
                    <RANKING order="3" place="3" resultid="3142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6316" />
                    <RANKING order="2" place="2" resultid="5500" />
                    <RANKING order="3" place="3" resultid="4286" />
                    <RANKING order="4" place="4" resultid="5005" />
                    <RANKING order="5" place="5" resultid="5389" />
                    <RANKING order="6" place="6" resultid="3157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4673" />
                    <RANKING order="2" place="2" resultid="4055" />
                    <RANKING order="3" place="3" resultid="3822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1249" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1251" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7796" daytime="11:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7797" daytime="11:07" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7798" daytime="11:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7799" daytime="11:13" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7800" daytime="11:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7801" daytime="11:17" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7802" daytime="11:19" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7803" daytime="11:21" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7804" daytime="11:23" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7805" daytime="11:25" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1254" daytime="11:27" gender="M" number="13" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1255" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3564" />
                    <RANKING order="2" place="2" resultid="6392" />
                    <RANKING order="3" place="3" resultid="2579" />
                    <RANKING order="4" place="4" resultid="5750" />
                    <RANKING order="5" place="5" resultid="6212" />
                    <RANKING order="6" place="6" resultid="6266" />
                    <RANKING order="7" place="7" resultid="4759" />
                    <RANKING order="8" place="-1" resultid="2224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5955" />
                    <RANKING order="2" place="2" resultid="5136" />
                    <RANKING order="3" place="3" resultid="5728" />
                    <RANKING order="4" place="4" resultid="5825" />
                    <RANKING order="5" place="5" resultid="4074" />
                    <RANKING order="6" place="6" resultid="3838" />
                    <RANKING order="7" place="7" resultid="5403" />
                    <RANKING order="8" place="8" resultid="6327" />
                    <RANKING order="9" place="9" resultid="3897" />
                    <RANKING order="10" place="10" resultid="5352" />
                    <RANKING order="11" place="11" resultid="3424" />
                    <RANKING order="12" place="12" resultid="4776" />
                    <RANKING order="13" place="13" resultid="2326" />
                    <RANKING order="14" place="14" resultid="5432" />
                    <RANKING order="15" place="15" resultid="2317" />
                    <RANKING order="16" place="16" resultid="5116" />
                    <RANKING order="17" place="17" resultid="3689" />
                    <RANKING order="18" place="-1" resultid="4065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1872" />
                    <RANKING order="2" place="2" resultid="1906" />
                    <RANKING order="3" place="3" resultid="2068" />
                    <RANKING order="4" place="4" resultid="5328" />
                    <RANKING order="5" place="5" resultid="5602" />
                    <RANKING order="6" place="6" resultid="4070" />
                    <RANKING order="7" place="7" resultid="3583" />
                    <RANKING order="8" place="8" resultid="4191" />
                    <RANKING order="9" place="9" resultid="1993" />
                    <RANKING order="10" place="10" resultid="3864" />
                    <RANKING order="11" place="11" resultid="6262" />
                    <RANKING order="12" place="12" resultid="5562" />
                    <RANKING order="13" place="13" resultid="4060" />
                    <RANKING order="14" place="14" resultid="6270" />
                    <RANKING order="15" place="15" resultid="4080" />
                    <RANKING order="16" place="16" resultid="2389" />
                    <RANKING order="17" place="17" resultid="4176" />
                    <RANKING order="18" place="18" resultid="3676" />
                    <RANKING order="19" place="19" resultid="4181" />
                    <RANKING order="20" place="20" resultid="5242" />
                    <RANKING order="21" place="21" resultid="5298" />
                    <RANKING order="22" place="22" resultid="4364" />
                    <RANKING order="23" place="-1" resultid="2034" />
                    <RANKING order="24" place="-1" resultid="3741" />
                    <RANKING order="25" place="-1" resultid="5775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6050" />
                    <RANKING order="2" place="2" resultid="2309" />
                    <RANKING order="3" place="3" resultid="2785" />
                    <RANKING order="4" place="4" resultid="5398" />
                    <RANKING order="5" place="5" resultid="2879" />
                    <RANKING order="6" place="6" resultid="3111" />
                    <RANKING order="7" place="7" resultid="2916" />
                    <RANKING order="8" place="8" resultid="2965" />
                    <RANKING order="9" place="9" resultid="5540" />
                    <RANKING order="10" place="10" resultid="4705" />
                    <RANKING order="11" place="11" resultid="5788" />
                    <RANKING order="12" place="12" resultid="1947" />
                    <RANKING order="13" place="13" resultid="3759" />
                    <RANKING order="14" place="14" resultid="4200" />
                    <RANKING order="15" place="15" resultid="4737" />
                    <RANKING order="16" place="16" resultid="2200" />
                    <RANKING order="17" place="17" resultid="6135" />
                    <RANKING order="18" place="18" resultid="2975" />
                    <RANKING order="19" place="19" resultid="3166" />
                    <RANKING order="20" place="20" resultid="5981" />
                    <RANKING order="21" place="21" resultid="3948" />
                    <RANKING order="22" place="22" resultid="3701" />
                    <RANKING order="23" place="23" resultid="4765" />
                    <RANKING order="24" place="24" resultid="5694" />
                    <RANKING order="25" place="25" resultid="3121" />
                    <RANKING order="26" place="26" resultid="3670" />
                    <RANKING order="27" place="-1" resultid="1927" />
                    <RANKING order="28" place="-1" resultid="2397" />
                    <RANKING order="29" place="-1" resultid="4103" />
                    <RANKING order="30" place="-1" resultid="4783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3329" />
                    <RANKING order="2" place="2" resultid="6175" />
                    <RANKING order="3" place="3" resultid="5737" />
                    <RANKING order="4" place="4" resultid="3577" />
                    <RANKING order="5" place="5" resultid="5190" />
                    <RANKING order="6" place="6" resultid="2775" />
                    <RANKING order="7" place="7" resultid="5217" />
                    <RANKING order="8" place="8" resultid="4430" />
                    <RANKING order="9" place="9" resultid="4701" />
                    <RANKING order="10" place="10" resultid="2115" />
                    <RANKING order="11" place="11" resultid="6207" />
                    <RANKING order="12" place="12" resultid="1977" />
                    <RANKING order="13" place="13" resultid="3466" />
                    <RANKING order="14" place="14" resultid="4748" />
                    <RANKING order="15" place="15" resultid="6358" />
                    <RANKING order="16" place="16" resultid="5701" />
                    <RANKING order="17" place="17" resultid="2234" />
                    <RANKING order="18" place="-1" resultid="3404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5124" />
                    <RANKING order="2" place="2" resultid="6193" />
                    <RANKING order="3" place="3" resultid="3636" />
                    <RANKING order="4" place="4" resultid="5886" />
                    <RANKING order="5" place="5" resultid="2855" />
                    <RANKING order="6" place="6" resultid="3233" />
                    <RANKING order="7" place="7" resultid="2367" />
                    <RANKING order="8" place="8" resultid="3393" />
                    <RANKING order="9" place="9" resultid="2040" />
                    <RANKING order="10" place="10" resultid="3093" />
                    <RANKING order="11" place="11" resultid="6228" />
                    <RANKING order="12" place="12" resultid="3918" />
                    <RANKING order="13" place="-1" resultid="5714" />
                    <RANKING order="14" place="-1" resultid="2185" />
                    <RANKING order="15" place="-1" resultid="3479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5292" />
                    <RANKING order="2" place="2" resultid="3255" />
                    <RANKING order="3" place="3" resultid="4471" />
                    <RANKING order="4" place="4" resultid="2544" />
                    <RANKING order="5" place="5" resultid="2352" />
                    <RANKING order="6" place="6" resultid="2828" />
                    <RANKING order="7" place="7" resultid="3182" />
                    <RANKING order="8" place="8" resultid="3649" />
                    <RANKING order="9" place="9" resultid="6038" />
                    <RANKING order="10" place="10" resultid="3170" />
                    <RANKING order="11" place="11" resultid="4724" />
                    <RANKING order="12" place="12" resultid="5288" />
                    <RANKING order="13" place="-1" resultid="2163" />
                    <RANKING order="14" place="-1" resultid="4537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5044" />
                    <RANKING order="2" place="2" resultid="5948" />
                    <RANKING order="3" place="3" resultid="1865" />
                    <RANKING order="4" place="4" resultid="4485" />
                    <RANKING order="5" place="5" resultid="6286" />
                    <RANKING order="6" place="6" resultid="5425" />
                    <RANKING order="7" place="7" resultid="5197" />
                    <RANKING order="8" place="8" resultid="6120" />
                    <RANKING order="9" place="9" resultid="4091" />
                    <RANKING order="10" place="-1" resultid="2640" />
                    <RANKING order="11" place="-1" resultid="3047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3513" />
                    <RANKING order="2" place="2" resultid="5648" />
                    <RANKING order="3" place="3" resultid="5866" />
                    <RANKING order="4" place="4" resultid="3409" />
                    <RANKING order="5" place="5" resultid="4301" />
                    <RANKING order="6" place="6" resultid="5536" />
                    <RANKING order="7" place="7" resultid="4542" />
                    <RANKING order="8" place="-1" resultid="2671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2706" />
                    <RANKING order="2" place="2" resultid="3813" />
                    <RANKING order="3" place="3" resultid="5023" />
                    <RANKING order="4" place="4" resultid="2406" />
                    <RANKING order="5" place="5" resultid="6445" />
                    <RANKING order="6" place="6" resultid="6249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4314" />
                    <RANKING order="2" place="2" resultid="5624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4455" />
                    <RANKING order="2" place="2" resultid="5620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2014" />
                    <RANKING order="2" place="2" resultid="1957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1269" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7806" daytime="11:27" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7807" daytime="11:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7808" daytime="11:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7809" daytime="11:37" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7810" daytime="11:39" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7811" daytime="11:41" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7812" daytime="11:43" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7813" daytime="11:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7814" daytime="11:47" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7815" daytime="11:49" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7816" daytime="11:51" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7817" daytime="11:53" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7818" daytime="11:55" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7819" daytime="11:56" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7820" daytime="11:58" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7821" daytime="12:00" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7822" daytime="12:02" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7823" daytime="12:04" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7824" daytime="12:05" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7825" daytime="12:07" number="20" order="20" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1270" daytime="12:09" gender="F" number="14" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1271" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2571" />
                    <RANKING order="2" place="2" resultid="1970" />
                    <RANKING order="3" place="3" resultid="2215" />
                    <RANKING order="4" place="4" resultid="2063" />
                    <RANKING order="5" place="5" resultid="2996" />
                    <RANKING order="6" place="6" resultid="2629" />
                    <RANKING order="7" place="7" resultid="3779" />
                    <RANKING order="8" place="8" resultid="2608" />
                    <RANKING order="9" place="9" resultid="3030" />
                    <RANKING order="10" place="10" resultid="5577" />
                    <RANKING order="11" place="11" resultid="3951" />
                    <RANKING order="12" place="12" resultid="1988" />
                    <RANKING order="13" place="-1" resultid="2002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3844" />
                    <RANKING order="2" place="2" resultid="4732" />
                    <RANKING order="3" place="3" resultid="5235" />
                    <RANKING order="4" place="4" resultid="3961" />
                    <RANKING order="5" place="5" resultid="4795" />
                    <RANKING order="6" place="6" resultid="3074" />
                    <RANKING order="7" place="7" resultid="3806" />
                    <RANKING order="8" place="8" resultid="1964" />
                    <RANKING order="9" place="9" resultid="6294" />
                    <RANKING order="10" place="10" resultid="3079" />
                    <RANKING order="11" place="11" resultid="5366" />
                    <RANKING order="12" place="-1" resultid="5793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5443" />
                    <RANKING order="2" place="2" resultid="3592" />
                    <RANKING order="3" place="3" resultid="5101" />
                    <RANKING order="4" place="4" resultid="4741" />
                    <RANKING order="5" place="5" resultid="6033" />
                    <RANKING order="6" place="6" resultid="4029" />
                    <RANKING order="7" place="7" resultid="6463" />
                    <RANKING order="8" place="8" resultid="5930" />
                    <RANKING order="9" place="9" resultid="2299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2928" />
                    <RANKING order="2" place="2" resultid="2936" />
                    <RANKING order="3" place="3" resultid="5409" />
                    <RANKING order="4" place="4" resultid="2943" />
                    <RANKING order="5" place="5" resultid="3384" />
                    <RANKING order="6" place="6" resultid="3695" />
                    <RANKING order="7" place="7" resultid="4021" />
                    <RANKING order="8" place="8" resultid="5900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5037" />
                    <RANKING order="2" place="2" resultid="5031" />
                    <RANKING order="3" place="3" resultid="3890" />
                    <RANKING order="4" place="4" resultid="3642" />
                    <RANKING order="5" place="5" resultid="5484" />
                    <RANKING order="6" place="6" resultid="2948" />
                    <RANKING order="7" place="7" resultid="3748" />
                    <RANKING order="8" place="8" resultid="4696" />
                    <RANKING order="9" place="9" resultid="6128" />
                    <RANKING order="10" place="10" resultid="6306" />
                    <RANKING order="11" place="11" resultid="4754" />
                    <RANKING order="12" place="-1" resultid="4548" />
                    <RANKING order="13" place="-1" resultid="6101" />
                    <RANKING order="14" place="-1" resultid="6218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4368" />
                    <RANKING order="2" place="2" resultid="3880" />
                    <RANKING order="3" place="3" resultid="2847" />
                    <RANKING order="4" place="4" resultid="6072" />
                    <RANKING order="5" place="5" resultid="6780" />
                    <RANKING order="6" place="6" resultid="3614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2138" />
                    <RANKING order="2" place="2" resultid="3039" />
                    <RANKING order="3" place="3" resultid="4994" />
                    <RANKING order="4" place="4" resultid="4987" />
                    <RANKING order="5" place="5" resultid="3597" />
                    <RANKING order="6" place="6" resultid="4619" />
                    <RANKING order="7" place="7" resultid="6364" />
                    <RANKING order="8" place="8" resultid="4683" />
                    <RANKING order="9" place="9" resultid="2265" />
                    <RANKING order="10" place="10" resultid="5937" />
                    <RANKING order="11" place="-1" resultid="3418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3398" />
                    <RANKING order="2" place="2" resultid="2129" />
                    <RANKING order="3" place="3" resultid="3731" />
                    <RANKING order="4" place="4" resultid="2256" />
                    <RANKING order="5" place="5" resultid="2008" />
                    <RANKING order="6" place="6" resultid="2531" />
                    <RANKING order="7" place="-1" resultid="4603" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4342" />
                    <RANKING order="2" place="2" resultid="5501" />
                    <RANKING order="3" place="3" resultid="5006" />
                    <RANKING order="4" place="4" resultid="3787" />
                    <RANKING order="5" place="5" resultid="3379" />
                    <RANKING order="6" place="6" resultid="4596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5394" />
                    <RANKING order="2" place="2" resultid="4325" />
                    <RANKING order="3" place="3" resultid="4356" />
                    <RANKING order="4" place="4" resultid="3823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4291" />
                    <RANKING order="2" place="2" resultid="5259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1284" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1285" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7826" daytime="12:09" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7827" daytime="12:13" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7828" daytime="12:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7829" daytime="12:19" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7830" daytime="12:21" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7831" daytime="12:23" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7832" daytime="12:26" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7833" daytime="12:28" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7834" daytime="12:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7835" daytime="12:32" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7836" daytime="12:34" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7837" daytime="12:36" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="12:39" gender="M" number="15" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1287" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6407" />
                    <RANKING order="2" place="2" resultid="2594" />
                    <RANKING order="3" place="3" resultid="6393" />
                    <RANKING order="4" place="4" resultid="2580" />
                    <RANKING order="5" place="5" resultid="2208" />
                    <RANKING order="6" place="6" resultid="2288" />
                    <RANKING order="7" place="7" resultid="3660" />
                    <RANKING order="8" place="-1" resultid="5689" />
                    <RANKING order="9" place="-1" resultid="6213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5357" />
                    <RANKING order="2" place="2" resultid="5826" />
                    <RANKING order="3" place="3" resultid="5142" />
                    <RANKING order="4" place="4" resultid="2023" />
                    <RANKING order="5" place="5" resultid="6328" />
                    <RANKING order="6" place="6" resultid="2588" />
                    <RANKING order="7" place="7" resultid="5809" />
                    <RANKING order="8" place="8" resultid="4513" />
                    <RANKING order="9" place="9" resultid="3520" />
                    <RANKING order="10" place="10" resultid="4777" />
                    <RANKING order="11" place="-1" resultid="2056" />
                    <RANKING order="12" place="-1" resultid="3251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5964" />
                    <RANKING order="2" place="2" resultid="2069" />
                    <RANKING order="3" place="3" resultid="4109" />
                    <RANKING order="4" place="4" resultid="4086" />
                    <RANKING order="5" place="5" resultid="4803" />
                    <RANKING order="6" place="6" resultid="5631" />
                    <RANKING order="7" place="7" resultid="4156" />
                    <RANKING order="8" place="8" resultid="3063" />
                    <RANKING order="9" place="9" resultid="2390" />
                    <RANKING order="10" place="10" resultid="3677" />
                    <RANKING order="11" place="11" resultid="4197" />
                    <RANKING order="12" place="12" resultid="5243" />
                    <RANKING order="13" place="13" resultid="4171" />
                    <RANKING order="14" place="14" resultid="4215" />
                    <RANKING order="15" place="-1" resultid="5776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1901" />
                    <RANKING order="2" place="2" resultid="2310" />
                    <RANKING order="3" place="3" resultid="2863" />
                    <RANKING order="4" place="4" resultid="6051" />
                    <RANKING order="5" place="5" resultid="2354" />
                    <RANKING order="6" place="6" resultid="6066" />
                    <RANKING order="7" place="7" resultid="2966" />
                    <RANKING order="8" place="8" resultid="2838" />
                    <RANKING order="9" place="9" resultid="5918" />
                    <RANKING order="10" place="10" resultid="1915" />
                    <RANKING order="11" place="11" resultid="4201" />
                    <RANKING order="12" place="12" resultid="2201" />
                    <RANKING order="13" place="13" resultid="2984" />
                    <RANKING order="14" place="14" resultid="1948" />
                    <RANKING order="15" place="15" resultid="5302" />
                    <RANKING order="16" place="16" resultid="2301" />
                    <RANKING order="17" place="17" resultid="3702" />
                    <RANKING order="18" place="-1" resultid="4706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2792" />
                    <RANKING order="2" place="2" resultid="5417" />
                    <RANKING order="3" place="3" resultid="6113" />
                    <RANKING order="4" place="4" resultid="3605" />
                    <RANKING order="5" place="5" resultid="3578" />
                    <RANKING order="6" place="6" resultid="5210" />
                    <RANKING order="7" place="7" resultid="5481" />
                    <RANKING order="8" place="8" resultid="2776" />
                    <RANKING order="9" place="9" resultid="6371" />
                    <RANKING order="10" place="10" resultid="6176" />
                    <RANKING order="11" place="11" resultid="2089" />
                    <RANKING order="12" place="12" resultid="5218" />
                    <RANKING order="13" place="13" resultid="2770" />
                    <RANKING order="14" place="14" resultid="2991" />
                    <RANKING order="15" place="15" resultid="2116" />
                    <RANKING order="16" place="16" resultid="3363" />
                    <RANKING order="17" place="17" resultid="5742" />
                    <RANKING order="18" place="18" resultid="2961" />
                    <RANKING order="19" place="19" resultid="3467" />
                    <RANKING order="20" place="20" resultid="4749" />
                    <RANKING order="21" place="21" resultid="6028" />
                    <RANKING order="22" place="22" resultid="3473" />
                    <RANKING order="23" place="-1" resultid="4331" />
                    <RANKING order="24" place="-1" resultid="4591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3655" />
                    <RANKING order="2" place="2" resultid="4374" />
                    <RANKING order="3" place="3" resultid="6194" />
                    <RANKING order="4" place="4" resultid="6338" />
                    <RANKING order="5" place="5" resultid="5346" />
                    <RANKING order="6" place="6" resultid="3867" />
                    <RANKING order="7" place="7" resultid="6059" />
                    <RANKING order="8" place="8" resultid="5708" />
                    <RANKING order="9" place="9" resultid="3094" />
                    <RANKING order="10" place="10" resultid="3725" />
                    <RANKING order="11" place="11" resultid="6205" />
                    <RANKING order="12" place="-1" resultid="2176" />
                    <RANKING order="13" place="-1" resultid="3265" />
                    <RANKING order="14" place="-1" resultid="3722" />
                    <RANKING order="15" place="-1" resultid="6399" />
                    <RANKING order="16" place="-1" resultid="3480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5293" />
                    <RANKING order="2" place="2" resultid="4037" />
                    <RANKING order="3" place="3" resultid="1921" />
                    <RANKING order="4" place="4" resultid="2545" />
                    <RANKING order="5" place="5" resultid="3831" />
                    <RANKING order="6" place="6" resultid="2357" />
                    <RANKING order="7" place="6" resultid="5893" />
                    <RANKING order="8" place="8" resultid="2250" />
                    <RANKING order="9" place="9" resultid="3226" />
                    <RANKING order="10" place="10" resultid="6039" />
                    <RANKING order="11" place="11" resultid="1886" />
                    <RANKING order="12" place="12" resultid="3771" />
                    <RANKING order="13" place="13" resultid="5267" />
                    <RANKING order="14" place="-1" resultid="3345" />
                    <RANKING order="15" place="-1" resultid="4660" />
                    <RANKING order="16" place="-1" resultid="4725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6006" />
                    <RANKING order="2" place="2" resultid="5184" />
                    <RANKING order="3" place="3" resultid="2537" />
                    <RANKING order="4" place="4" resultid="3318" />
                    <RANKING order="5" place="5" resultid="2624" />
                    <RANKING order="6" place="6" resultid="5638" />
                    <RANKING order="7" place="7" resultid="3609" />
                    <RANKING order="8" place="8" resultid="3622" />
                    <RANKING order="9" place="9" resultid="1866" />
                    <RANKING order="10" place="10" resultid="5522" />
                    <RANKING order="11" place="11" resultid="4486" />
                    <RANKING order="12" place="-1" resultid="2152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4422" />
                    <RANKING order="2" place="2" resultid="5649" />
                    <RANKING order="3" place="3" resultid="4612" />
                    <RANKING order="4" place="4" resultid="2811" />
                    <RANKING order="5" place="5" resultid="5656" />
                    <RANKING order="6" place="6" resultid="2047" />
                    <RANKING order="7" place="7" resultid="2146" />
                    <RANKING order="8" place="8" resultid="4689" />
                    <RANKING order="9" place="-1" resultid="3449" />
                    <RANKING order="10" place="-1" resultid="5609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2239" />
                    <RANKING order="2" place="2" resultid="5508" />
                    <RANKING order="3" place="3" resultid="5024" />
                    <RANKING order="4" place="4" resultid="3801" />
                    <RANKING order="5" place="5" resultid="4504" />
                    <RANKING order="6" place="6" resultid="4360" />
                    <RANKING order="7" place="7" resultid="3303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4296" />
                    <RANKING order="2" place="2" resultid="3554" />
                    <RANKING order="3" place="3" resultid="3794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1298" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1299" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2616" />
                    <RANKING order="2" place="2" resultid="2663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1300" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1301" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7838" daytime="12:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7839" daytime="12:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7840" daytime="12:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7841" daytime="12:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7842" daytime="12:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7843" daytime="12:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7844" daytime="12:54" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7845" daytime="12:57" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7846" daytime="12:59" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7847" daytime="13:01" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7848" daytime="13:03" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7849" daytime="13:05" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7850" daytime="13:07" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7851" daytime="13:09" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7852" daytime="13:11" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7853" daytime="13:13" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7854" daytime="13:15" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7855" daytime="13:17" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7856" daytime="13:18" number="19" order="19" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="13:21" gender="F" number="16" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1303" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6022" />
                    <RANKING order="2" place="2" resultid="5310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="34" agemin="30" name="Kategoria B" />
                <AGEGROUP agegroupid="1306" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="44" agemin="40" name="Kategoria D" />
                <AGEGROUP agegroupid="1308" agemax="49" agemin="45" name="Kategoria E" />
                <AGEGROUP agegroupid="1309" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3936" />
                    <RANKING order="2" place="2" resultid="3134" />
                    <RANKING order="3" place="3" resultid="4556" />
                    <RANKING order="4" place="-1" resultid="4627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="64" agemin="60" name="Kategoria H" />
                <AGEGROUP agegroupid="1312" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="1313" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="1314" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1315" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1316" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1317" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7857" daytime="13:21" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7858" daytime="13:29" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1318" daytime="13:35" gender="M" number="17" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1319" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5158" />
                    <RANKING order="2" place="2" resultid="2561" />
                    <RANKING order="3" place="-1" resultid="3534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1320" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6277" />
                    <RANKING order="2" place="2" resultid="2277" />
                    <RANKING order="3" place="3" resultid="2029" />
                    <RANKING order="4" place="-1" resultid="2635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1321" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1907" />
                    <RANKING order="2" place="2" resultid="3246" />
                    <RANKING order="3" place="3" resultid="4228" />
                    <RANKING order="4" place="4" resultid="5820" />
                    <RANKING order="5" place="-1" resultid="4717" />
                    <RANKING order="6" place="-1" resultid="5589" />
                    <RANKING order="7" place="-1" resultid="5777" />
                    <RANKING order="8" place="-1" resultid="3497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1322" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2971" />
                    <RANKING order="2" place="2" resultid="5202" />
                    <RANKING order="3" place="3" resultid="2871" />
                    <RANKING order="4" place="4" resultid="5695" />
                    <RANKING order="5" place="-1" resultid="5919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1323" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2793" />
                    <RANKING order="2" place="2" resultid="3855" />
                    <RANKING order="3" place="3" resultid="6299" />
                    <RANKING order="4" place="4" resultid="4320" />
                    <RANKING order="5" place="5" resultid="5743" />
                    <RANKING order="6" place="-1" resultid="2730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1324" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1325" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2829" />
                    <RANKING order="2" place="2" resultid="3211" />
                    <RANKING order="3" place="3" resultid="5018" />
                    <RANKING order="4" place="4" resultid="5319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1326" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2554" />
                    <RANKING order="2" place="2" resultid="4464" />
                    <RANKING order="3" place="3" resultid="2752" />
                    <RANKING order="4" place="-1" resultid="6007" />
                    <RANKING order="5" place="-1" resultid="3048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4477" />
                    <RANKING order="2" place="2" resultid="5867" />
                    <RANKING order="3" place="3" resultid="3189" />
                    <RANKING order="4" place="4" resultid="2653" />
                    <RANKING order="5" place="5" resultid="4584" />
                    <RANKING order="6" place="6" resultid="3458" />
                    <RANKING order="7" place="-1" resultid="4979" />
                    <RANKING order="8" place="-1" resultid="5610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1328" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2240" />
                    <RANKING order="2" place="2" resultid="2737" />
                    <RANKING order="3" place="3" resultid="5025" />
                    <RANKING order="4" place="4" resultid="3814" />
                    <RANKING order="5" place="5" resultid="3293" />
                    <RANKING order="6" place="6" resultid="1895" />
                    <RANKING order="7" place="-1" resultid="6223" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1329" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2745" />
                    <RANKING order="2" place="2" resultid="6235" />
                    <RANKING order="3" place="-1" resultid="6252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1330" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1331" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1332" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1333" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7859" daytime="13:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7860" daytime="13:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7861" daytime="13:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7862" daytime="13:51" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7863" daytime="13:56" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7864" daytime="13:59" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7865" daytime="14:03" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1334" daytime="14:07" gender="F" number="18" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1350" agemax="96" agemin="80" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="1351" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3973" />
                    <RANKING order="2" place="2" resultid="3001" />
                    <RANKING order="3" place="3" resultid="6079" />
                    <RANKING order="4" place="4" resultid="4118" />
                    <RANKING order="5" place="5" resultid="5987" />
                    <RANKING order="6" place="6" resultid="3088" />
                    <RANKING order="7" place="-1" resultid="6452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5050" />
                    <RANKING order="2" place="-1" resultid="5799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3987" />
                    <RANKING order="2" place="2" resultid="4631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1355" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1356" agemax="400" agemin="280" name="Kategoria F" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7866" daytime="14:07" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7867" daytime="14:11" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1357" daytime="14:15" gender="M" number="19" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1358" agemax="96" agemin="80" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="1359" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6449" />
                    <RANKING order="2" place="-1" resultid="6409" />
                    <RANKING order="3" place="-1" resultid="2077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1360" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3269" />
                    <RANKING order="2" place="2" resultid="4120" />
                    <RANKING order="3" place="3" resultid="5754" />
                    <RANKING order="4" place="4" resultid="4812" />
                    <RANKING order="5" place="5" resultid="4122" />
                    <RANKING order="6" place="6" resultid="3982" />
                    <RANKING order="7" place="7" resultid="6453" />
                    <RANKING order="8" place="8" resultid="4245" />
                    <RANKING order="9" place="9" resultid="4247" />
                    <RANKING order="10" place="10" resultid="2336" />
                    <RANKING order="11" place="11" resultid="4248" />
                    <RANKING order="12" place="-1" resultid="3709" />
                    <RANKING order="13" place="-1" resultid="2043" />
                    <RANKING order="14" place="-1" resultid="3086" />
                    <RANKING order="15" place="-1" resultid="5667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1361" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2884" />
                    <RANKING order="2" place="2" resultid="6081" />
                    <RANKING order="3" place="3" resultid="5224" />
                    <RANKING order="4" place="4" resultid="3271" />
                    <RANKING order="5" place="5" resultid="4518" />
                    <RANKING order="6" place="6" resultid="2096" />
                    <RANKING order="7" place="7" resultid="4814" />
                    <RANKING order="8" place="8" resultid="5717" />
                    <RANKING order="9" place="-1" resultid="8769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1362" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3985" />
                    <RANKING order="2" place="2" resultid="4382" />
                    <RANKING order="3" place="3" resultid="5988" />
                    <RANKING order="4" place="4" resultid="2379" />
                    <RANKING order="5" place="5" resultid="3501" />
                    <RANKING order="6" place="-1" resultid="2189" />
                    <RANKING order="7" place="-1" resultid="8761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1363" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5052" />
                    <RANKING order="2" place="2" resultid="5544" />
                    <RANKING order="3" place="3" resultid="4516" />
                    <RANKING order="4" place="4" resultid="5663" />
                    <RANKING order="5" place="-1" resultid="4633" />
                    <RANKING order="6" place="-1" resultid="8782" />
                    <RANKING order="7" place="-1" resultid="2645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1364" agemax="400" agemin="280" name="Kategoria F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4381" />
                    <RANKING order="2" place="-1" resultid="5665" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7868" daytime="14:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7869" daytime="14:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7870" daytime="14:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7871" daytime="14:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7872" daytime="14:29" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="8925" />
            <JUDGE officialid="8910" />
            <JUDGE officialid="8924" />
            <JUDGE officialid="8926" />
            <JUDGE officialid="8906" />
            <JUDGE officialid="8919" />
            <JUDGE officialid="8923" />
            <JUDGE officialid="8909" />
            <JUDGE officialid="8921" />
            <JUDGE officialid="8914" />
            <JUDGE officialid="8915" />
            <JUDGE officialid="8918" />
            <JUDGE officialid="8922" />
            <JUDGE officialid="8917" />
            <JUDGE officialid="8920" />
            <JUDGE officialid="8928" />
            <JUDGE officialid="8912" />
            <JUDGE officialid="8916" />
            <JUDGE officialid="8916" />
            <JUDGE officialid="8908" />
            <JUDGE officialid="8908" />
            <JUDGE officialid="8911" />
            <JUDGE officialid="8911" />
            <JUDGE officialid="8913" />
            <JUDGE officialid="8927" />
            <JUDGE officialid="8905" />
            <JUDGE officialid="8904" />
            <JUDGE officialid="8903" />
            <JUDGE officialid="8907" />
            <JUDGE officialid="8941" />
            <JUDGE officialid="8901" />
            <JUDGE officialid="8902" />
          </JUDGES>
        </SESSION>
        <SESSION date="2013-11-16" daytime="16:15" name="MP Masters BLOK III" number="3" warmupfrom="15:00" warmupuntil="15:55">
          <EVENTS>
            <EVENT eventid="1366" daytime="16:15" gender="F" number="20" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1368" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2572" />
                    <RANKING order="2" place="2" resultid="2216" />
                    <RANKING order="3" place="3" resultid="5578" />
                    <RANKING order="4" place="4" resultid="5110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1369" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5569" />
                    <RANKING order="2" place="2" resultid="3542" />
                    <RANKING order="3" place="3" resultid="3962" />
                    <RANKING order="4" place="4" resultid="3807" />
                    <RANKING order="5" place="5" resultid="1965" />
                    <RANKING order="6" place="6" resultid="4411" />
                    <RANKING order="7" place="-1" resultid="6296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1370" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4043" />
                    <RANKING order="2" place="2" resultid="5102" />
                    <RANKING order="3" place="3" resultid="5931" />
                    <RANKING order="4" place="-1" resultid="4098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1371" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2929" />
                    <RANKING order="2" place="2" resultid="5410" />
                    <RANKING order="3" place="3" resultid="5131" />
                    <RANKING order="4" place="4" resultid="3489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1372" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2677" />
                    <RANKING order="2" place="2" resultid="4307" />
                    <RANKING order="3" place="3" resultid="6384" />
                    <RANKING order="4" place="4" resultid="2953" />
                    <RANKING order="5" place="5" resultid="4697" />
                    <RANKING order="6" place="6" resultid="5881" />
                    <RANKING order="7" place="7" resultid="3069" />
                    <RANKING order="8" place="8" resultid="3874" />
                    <RANKING order="9" place="-1" resultid="6102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1373" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5172" />
                    <RANKING order="2" place="2" resultid="5372" />
                    <RANKING order="3" place="3" resultid="2848" />
                    <RANKING order="4" place="4" resultid="6469" />
                    <RANKING order="5" place="5" resultid="6467" />
                    <RANKING order="6" place="-1" resultid="6781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1374" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4995" />
                    <RANKING order="2" place="2" resultid="3885" />
                    <RANKING order="3" place="3" resultid="6365" />
                    <RANKING order="4" place="4" resultid="4620" />
                    <RANKING order="5" place="5" resultid="3598" />
                    <RANKING order="6" place="6" resultid="5938" />
                    <RANKING order="7" place="7" resultid="3573" />
                    <RANKING order="8" place="8" resultid="4684" />
                    <RANKING order="9" place="9" resultid="2266" />
                    <RANKING order="10" place="10" resultid="2763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1375" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2257" />
                    <RANKING order="2" place="2" resultid="4604" />
                    <RANKING order="3" place="3" resultid="2532" />
                    <RANKING order="4" place="-1" resultid="3143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1376" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6169" />
                    <RANKING order="2" place="2" resultid="3788" />
                    <RANKING order="3" place="3" resultid="4597" />
                    <RANKING order="4" place="4" resultid="3158" />
                    <RANKING order="5" place="-1" resultid="5007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1377" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1378" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4272" />
                    <RANKING order="2" place="2" resultid="6345" />
                    <RANKING order="3" place="3" resultid="5260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1379" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3117" />
                    <RANKING order="2" place="2" resultid="2124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1380" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1381" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1382" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7873" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7874" daytime="16:19" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7875" daytime="16:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7876" daytime="16:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7877" daytime="16:28" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7878" daytime="16:31" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7879" daytime="16:33" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7880" daytime="16:36" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1383" daytime="16:38" gender="M" number="21" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1384" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5159" />
                    <RANKING order="2" place="2" resultid="2283" />
                    <RANKING order="3" place="3" resultid="6243" />
                    <RANKING order="4" place="4" resultid="3549" />
                    <RANKING order="5" place="5" resultid="2209" />
                    <RANKING order="6" place="6" resultid="2289" />
                    <RANKING order="7" place="7" resultid="2562" />
                    <RANKING order="8" place="-1" resultid="3535" />
                    <RANKING order="9" place="-1" resultid="5690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1385" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5358" />
                    <RANKING order="2" place="2" resultid="5817" />
                    <RANKING order="3" place="3" resultid="2024" />
                    <RANKING order="4" place="4" resultid="5810" />
                    <RANKING order="5" place="5" resultid="5813" />
                    <RANKING order="6" place="6" resultid="5353" />
                    <RANKING order="7" place="7" resultid="2327" />
                    <RANKING order="8" place="-1" resultid="5382" />
                    <RANKING order="9" place="-1" resultid="2057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1386" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5965" />
                    <RANKING order="2" place="2" resultid="4087" />
                    <RANKING order="3" place="3" resultid="6044" />
                    <RANKING order="4" place="4" resultid="4110" />
                    <RANKING order="5" place="5" resultid="4187" />
                    <RANKING order="6" place="6" resultid="3064" />
                    <RANKING order="7" place="7" resultid="3678" />
                    <RANKING order="8" place="8" resultid="2331" />
                    <RANKING order="9" place="9" resultid="4166" />
                    <RANKING order="10" place="10" resultid="4172" />
                    <RANKING order="11" place="11" resultid="4216" />
                    <RANKING order="12" place="12" resultid="2758" />
                    <RANKING order="13" place="-1" resultid="5596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1387" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2864" />
                    <RANKING order="2" place="2" resultid="2880" />
                    <RANKING order="3" place="3" resultid="3338" />
                    <RANKING order="4" place="4" resultid="3350" />
                    <RANKING order="5" place="5" resultid="5541" />
                    <RANKING order="6" place="6" resultid="5789" />
                    <RANKING order="7" place="7" resultid="2839" />
                    <RANKING order="8" place="8" resultid="2872" />
                    <RANKING order="9" place="9" resultid="2985" />
                    <RANKING order="10" place="10" resultid="2202" />
                    <RANKING order="11" place="11" resultid="2322" />
                    <RANKING order="12" place="12" resultid="5303" />
                    <RANKING order="13" place="13" resultid="6136" />
                    <RANKING order="14" place="14" resultid="5913" />
                    <RANKING order="15" place="15" resultid="5437" />
                    <RANKING order="16" place="16" resultid="5926" />
                    <RANKING order="17" place="17" resultid="3671" />
                    <RANKING order="18" place="-1" resultid="4784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1388" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2794" />
                    <RANKING order="2" place="2" resultid="2715" />
                    <RANKING order="3" place="3" resultid="3665" />
                    <RANKING order="4" place="4" resultid="6359" />
                    <RANKING order="5" place="5" resultid="2731" />
                    <RANKING order="6" place="6" resultid="3474" />
                    <RANKING order="7" place="-1" resultid="5211" />
                    <RANKING order="8" place="-1" resultid="6114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1389" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5125" />
                    <RANKING order="2" place="2" resultid="3017" />
                    <RANKING order="3" place="3" resultid="3868" />
                    <RANKING order="4" place="4" resultid="5530" />
                    <RANKING order="5" place="5" resultid="2169" />
                    <RANKING order="6" place="6" resultid="5378" />
                    <RANKING order="7" place="7" resultid="5709" />
                    <RANKING order="8" place="8" resultid="3389" />
                    <RANKING order="9" place="9" resultid="3095" />
                    <RANKING order="10" place="10" resultid="3726" />
                    <RANKING order="11" place="11" resultid="5274" />
                    <RANKING order="12" place="12" resultid="3765" />
                    <RANKING order="13" place="-1" resultid="3266" />
                    <RANKING order="14" place="-1" resultid="3481" />
                    <RANKING order="15" place="-1" resultid="3919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1390" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4661" />
                    <RANKING order="2" place="2" resultid="5894" />
                    <RANKING order="3" place="3" resultid="3227" />
                    <RANKING order="4" place="4" resultid="2251" />
                    <RANKING order="5" place="5" resultid="3325" />
                    <RANKING order="6" place="6" resultid="2158" />
                    <RANKING order="7" place="7" resultid="5013" />
                    <RANKING order="8" place="8" resultid="1887" />
                    <RANKING order="9" place="9" resultid="3261" />
                    <RANKING order="10" place="-1" resultid="2711" />
                    <RANKING order="11" place="-1" resultid="4538" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3334" />
                    <RANKING order="2" place="2" resultid="2555" />
                    <RANKING order="3" place="3" resultid="4959" />
                    <RANKING order="4" place="4" resultid="3624" />
                    <RANKING order="5" place="5" resultid="5639" />
                    <RANKING order="6" place="6" resultid="4499" />
                    <RANKING order="7" place="7" resultid="2153" />
                    <RANKING order="8" place="8" resultid="3627" />
                    <RANKING order="9" place="9" resultid="3204" />
                    <RANKING order="10" place="10" resultid="3197" />
                    <RANKING order="11" place="11" resultid="5426" />
                    <RANKING order="12" place="12" resultid="2753" />
                    <RANKING order="13" place="-1" resultid="4092" />
                    <RANKING order="14" place="-1" resultid="4136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1392" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4423" />
                    <RANKING order="2" place="2" resultid="4478" />
                    <RANKING order="3" place="3" resultid="2048" />
                    <RANKING order="4" place="4" resultid="6184" />
                    <RANKING order="5" place="5" resultid="5643" />
                    <RANKING order="6" place="6" resultid="4690" />
                    <RANKING order="7" place="7" resultid="3190" />
                    <RANKING order="8" place="8" resultid="4585" />
                    <RANKING order="9" place="9" resultid="5657" />
                    <RANKING order="10" place="10" resultid="3459" />
                    <RANKING order="11" place="-1" resultid="3632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1393" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5000" />
                    <RANKING order="2" place="2" resultid="2686" />
                    <RANKING order="3" place="3" resultid="2724" />
                    <RANKING order="4" place="4" resultid="5509" />
                    <RANKING order="5" place="5" resultid="3304" />
                    <RANKING order="6" place="6" resultid="3152" />
                    <RANKING order="7" place="-1" resultid="2738" />
                    <RANKING order="8" place="-1" resultid="5617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1394" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4315" />
                    <RANKING order="2" place="2" resultid="4277" />
                    <RANKING order="3" place="3" resultid="4572" />
                    <RANKING order="4" place="4" resultid="2746" />
                    <RANKING order="5" place="5" resultid="1998" />
                    <RANKING order="6" place="-1" resultid="4439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1395" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4579" />
                    <RANKING order="2" place="2" resultid="5972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1396" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2664" />
                    <RANKING order="2" place="2" resultid="2362" />
                    <RANKING order="3" place="3" resultid="4495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1398" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7881" daytime="16:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7882" daytime="16:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7883" daytime="16:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7884" daytime="16:47" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7885" daytime="16:49" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7886" daytime="16:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7887" daytime="16:54" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7888" daytime="16:57" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7889" daytime="16:59" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7890" daytime="17:01" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7891" daytime="17:03" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7892" daytime="17:05" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7893" daytime="17:07" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7894" daytime="17:09" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7895" daytime="17:12" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7896" daytime="17:13" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1399" daytime="17:16" gender="F" number="22" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1400" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1971" />
                    <RANKING order="2" place="2" resultid="2064" />
                    <RANKING order="3" place="3" resultid="3780" />
                    <RANKING order="4" place="4" resultid="2997" />
                    <RANKING order="5" place="5" resultid="3031" />
                    <RANKING order="6" place="6" resultid="5841" />
                    <RANKING order="7" place="7" resultid="2217" />
                    <RANKING order="8" place="8" resultid="3952" />
                    <RANKING order="9" place="9" resultid="6256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1401" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5570" />
                    <RANKING order="2" place="2" resultid="6023" />
                    <RANKING order="3" place="3" resultid="3543" />
                    <RANKING order="4" place="4" resultid="5236" />
                    <RANKING order="5" place="5" resultid="4796" />
                    <RANKING order="6" place="6" resultid="3963" />
                    <RANKING order="7" place="7" resultid="2648" />
                    <RANKING order="8" place="8" resultid="3075" />
                    <RANKING order="9" place="9" resultid="2585" />
                    <RANKING order="10" place="10" resultid="5311" />
                    <RANKING order="11" place="11" resultid="6297" />
                    <RANKING order="12" place="12" resultid="3080" />
                    <RANKING order="13" place="13" resultid="5362" />
                    <RANKING order="14" place="-1" resultid="5367" />
                    <RANKING order="15" place="-1" resultid="5794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1402" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5444" />
                    <RANKING order="2" place="2" resultid="4044" />
                    <RANKING order="3" place="3" resultid="5875" />
                    <RANKING order="4" place="4" resultid="4742" />
                    <RANKING order="5" place="5" resultid="6034" />
                    <RANKING order="6" place="6" resultid="6015" />
                    <RANKING order="7" place="7" resultid="6464" />
                    <RANKING order="8" place="8" resultid="3684" />
                    <RANKING order="9" place="9" resultid="3754" />
                    <RANKING order="10" place="-1" resultid="4099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1403" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5411" />
                    <RANKING order="2" place="2" resultid="3385" />
                    <RANKING order="3" place="3" resultid="2937" />
                    <RANKING order="4" place="4" resultid="2944" />
                    <RANKING order="5" place="5" resultid="5901" />
                    <RANKING order="6" place="-1" resultid="3696" />
                    <RANKING order="7" place="-1" resultid="5765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1404" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4549" />
                    <RANKING order="2" place="2" resultid="5038" />
                    <RANKING order="3" place="3" resultid="3891" />
                    <RANKING order="4" place="4" resultid="3749" />
                    <RANKING order="5" place="5" resultid="6219" />
                    <RANKING order="6" place="6" resultid="6307" />
                    <RANKING order="7" place="7" resultid="6129" />
                    <RANKING order="8" place="-1" resultid="6103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1405" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5173" />
                    <RANKING order="2" place="2" resultid="4369" />
                    <RANKING order="3" place="3" resultid="3881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1406" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4988" />
                    <RANKING order="2" place="2" resultid="4996" />
                    <RANKING order="3" place="3" resultid="5179" />
                    <RANKING order="4" place="4" resultid="3937" />
                    <RANKING order="5" place="5" resultid="4621" />
                    <RANKING order="6" place="6" resultid="3323" />
                    <RANKING order="7" place="7" resultid="5939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1407" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2130" />
                    <RANKING order="2" place="2" resultid="3732" />
                    <RANKING order="3" place="3" resultid="3928" />
                    <RANKING order="4" place="-1" resultid="4605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1408" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4343" />
                    <RANKING order="2" place="2" resultid="5502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1409" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4357" />
                    <RANKING order="2" place="2" resultid="3824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1412" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1413" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1414" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7897" daytime="17:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7898" daytime="17:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7899" daytime="17:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7900" daytime="17:21" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7901" daytime="17:23" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7902" daytime="17:24" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7903" daytime="17:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7904" daytime="17:27" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7905" daytime="17:28" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1415" daytime="17:30" gender="M" number="23" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1416" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3565" />
                    <RANKING order="2" place="2" resultid="6394" />
                    <RANKING order="3" place="3" resultid="6408" />
                    <RANKING order="4" place="4" resultid="2595" />
                    <RANKING order="5" place="5" resultid="2581" />
                    <RANKING order="6" place="6" resultid="5751" />
                    <RANKING order="7" place="7" resultid="6214" />
                    <RANKING order="8" place="8" resultid="6267" />
                    <RANKING order="9" place="9" resultid="2563" />
                    <RANKING order="10" place="-1" resultid="2225" />
                    <RANKING order="11" place="-1" resultid="2290" />
                    <RANKING order="12" place="-1" resultid="3536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1417" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5956" />
                    <RANKING order="2" place="2" resultid="6329" />
                    <RANKING order="3" place="3" resultid="6278" />
                    <RANKING order="4" place="4" resultid="5137" />
                    <RANKING order="5" place="5" resultid="4075" />
                    <RANKING order="6" place="6" resultid="3521" />
                    <RANKING order="7" place="7" resultid="5383" />
                    <RANKING order="8" place="8" resultid="3898" />
                    <RANKING order="9" place="9" resultid="5354" />
                    <RANKING order="10" place="10" resultid="5433" />
                    <RANKING order="11" place="11" resultid="5117" />
                    <RANKING order="12" place="12" resultid="2058" />
                    <RANKING order="13" place="-1" resultid="3690" />
                    <RANKING order="14" place="-1" resultid="2318" />
                    <RANKING order="15" place="-1" resultid="2636" />
                    <RANKING order="16" place="-1" resultid="4066" />
                    <RANKING order="17" place="-1" resultid="5734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1418" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1873" />
                    <RANKING order="2" place="2" resultid="4771" />
                    <RANKING order="3" place="3" resultid="1908" />
                    <RANKING order="4" place="4" resultid="5966" />
                    <RANKING order="5" place="5" resultid="4229" />
                    <RANKING order="6" place="6" resultid="3247" />
                    <RANKING order="7" place="7" resultid="4071" />
                    <RANKING order="8" place="8" resultid="2070" />
                    <RANKING order="9" place="9" resultid="4192" />
                    <RANKING order="10" place="10" resultid="4111" />
                    <RANKING order="11" place="11" resultid="3059" />
                    <RANKING order="12" place="12" resultid="4081" />
                    <RANKING order="13" place="12" resultid="6271" />
                    <RANKING order="14" place="14" resultid="4182" />
                    <RANKING order="15" place="15" resultid="2391" />
                    <RANKING order="16" place="16" resultid="4718" />
                    <RANKING order="17" place="17" resultid="4177" />
                    <RANKING order="18" place="18" resultid="5590" />
                    <RANKING order="19" place="19" resultid="3528" />
                    <RANKING order="20" place="20" resultid="5244" />
                    <RANKING order="21" place="-1" resultid="2035" />
                    <RANKING order="22" place="-1" resultid="3498" />
                    <RANKING order="23" place="-1" resultid="5563" />
                    <RANKING order="24" place="-1" resultid="5778" />
                    <RANKING order="25" place="-1" resultid="6263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5556" />
                    <RANKING order="2" place="2" resultid="6052" />
                    <RANKING order="3" place="3" resultid="2355" />
                    <RANKING order="4" place="4" resultid="6067" />
                    <RANKING order="5" place="5" resultid="4707" />
                    <RANKING order="6" place="6" resultid="2917" />
                    <RANKING order="7" place="7" resultid="5399" />
                    <RANKING order="8" place="8" resultid="1928" />
                    <RANKING order="9" place="9" resultid="4209" />
                    <RANKING order="10" place="10" resultid="2967" />
                    <RANKING order="11" place="11" resultid="2398" />
                    <RANKING order="12" place="12" resultid="5203" />
                    <RANKING order="13" place="13" resultid="2302" />
                    <RANKING order="14" place="14" resultid="4104" />
                    <RANKING order="15" place="15" resultid="4202" />
                    <RANKING order="16" place="16" resultid="5304" />
                    <RANKING order="17" place="17" resultid="1949" />
                    <RANKING order="18" place="18" resultid="5696" />
                    <RANKING order="19" place="-1" resultid="2644" />
                    <RANKING order="20" place="-1" resultid="3703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1420" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3330" />
                    <RANKING order="2" place="2" resultid="2795" />
                    <RANKING order="3" place="3" resultid="5418" />
                    <RANKING order="4" place="4" resultid="4332" />
                    <RANKING order="5" place="5" resultid="3944" />
                    <RANKING order="6" place="6" resultid="6300" />
                    <RANKING order="7" place="7" resultid="2092" />
                    <RANKING order="8" place="8" resultid="2716" />
                    <RANKING order="9" place="9" resultid="6115" />
                    <RANKING order="10" place="10" resultid="5482" />
                    <RANKING order="11" place="11" resultid="5191" />
                    <RANKING order="12" place="12" resultid="4321" />
                    <RANKING order="13" place="13" resultid="5219" />
                    <RANKING order="14" place="14" resultid="6177" />
                    <RANKING order="15" place="15" resultid="4431" />
                    <RANKING order="16" place="16" resultid="5744" />
                    <RANKING order="17" place="17" resultid="4702" />
                    <RANKING order="18" place="18" resultid="2962" />
                    <RANKING order="19" place="19" resultid="2117" />
                    <RANKING order="20" place="20" resultid="6360" />
                    <RANKING order="21" place="21" resultid="3468" />
                    <RANKING order="22" place="22" resultid="6029" />
                    <RANKING order="23" place="23" resultid="5702" />
                    <RANKING order="24" place="-1" resultid="3606" />
                    <RANKING order="25" place="-1" resultid="4592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1421" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4375" />
                    <RANKING order="2" place="2" resultid="2856" />
                    <RANKING order="3" place="3" resultid="3869" />
                    <RANKING order="4" place="4" resultid="2170" />
                    <RANKING order="5" place="5" resultid="3096" />
                    <RANKING order="6" place="6" resultid="5275" />
                    <RANKING order="7" place="7" resultid="5715" />
                    <RANKING order="8" place="-1" resultid="2186" />
                    <RANKING order="9" place="-1" resultid="3267" />
                    <RANKING order="10" place="-1" resultid="6401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1422" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4472" />
                    <RANKING order="2" place="2" resultid="2546" />
                    <RANKING order="3" place="3" resultid="3832" />
                    <RANKING order="4" place="4" resultid="2691" />
                    <RANKING order="5" place="5" resultid="3346" />
                    <RANKING order="6" place="6" resultid="2603" />
                    <RANKING order="7" place="7" resultid="1888" />
                    <RANKING order="8" place="8" resultid="4726" />
                    <RANKING order="9" place="9" resultid="5268" />
                    <RANKING order="10" place="-1" resultid="3183" />
                    <RANKING order="11" place="-1" resultid="2164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1423" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5185" />
                    <RANKING order="2" place="2" resultid="6008" />
                    <RANKING order="3" place="3" resultid="2538" />
                    <RANKING order="4" place="4" resultid="5949" />
                    <RANKING order="5" place="5" resultid="4465" />
                    <RANKING order="6" place="6" resultid="4487" />
                    <RANKING order="7" place="7" resultid="3315" />
                    <RANKING order="8" place="8" resultid="3175" />
                    <RANKING order="9" place="9" resultid="3198" />
                    <RANKING order="10" place="-1" resultid="4093" />
                    <RANKING order="11" place="-1" resultid="5045" />
                    <RANKING order="12" place="-1" resultid="6287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1424" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3514" />
                    <RANKING order="2" place="2" resultid="5868" />
                    <RANKING order="3" place="3" resultid="4302" />
                    <RANKING order="4" place="4" resultid="5650" />
                    <RANKING order="5" place="5" resultid="2147" />
                    <RANKING order="6" place="6" resultid="5537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2241" />
                    <RANKING order="2" place="2" resultid="2681" />
                    <RANKING order="3" place="3" resultid="6224" />
                    <RANKING order="4" place="4" resultid="5026" />
                    <RANKING order="5" place="5" resultid="6446" />
                    <RANKING order="6" place="6" resultid="4509" />
                    <RANKING order="7" place="7" resultid="4361" />
                    <RANKING order="8" place="8" resultid="4505" />
                    <RANKING order="9" place="9" resultid="1894" />
                    <RANKING order="10" place="-1" resultid="3802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6253" />
                    <RANKING order="2" place="2" resultid="4297" />
                    <RANKING order="3" place="3" resultid="4278" />
                    <RANKING order="4" place="4" resultid="3555" />
                    <RANKING order="5" place="5" resultid="4573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1879" />
                    <RANKING order="2" place="2" resultid="4456" />
                    <RANKING order="3" place="3" resultid="5252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3311" />
                    <RANKING order="2" place="2" resultid="2617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1430" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7906" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7907" daytime="17:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7908" daytime="17:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7909" daytime="17:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7910" daytime="17:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7911" daytime="17:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7912" daytime="17:39" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7913" daytime="17:40" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7914" daytime="17:42" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7915" daytime="17:43" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7916" daytime="17:44" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7917" daytime="17:46" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7918" daytime="17:47" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7919" daytime="17:48" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7920" daytime="17:49" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7921" daytime="17:51" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7922" daytime="17:52" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7923" daytime="17:53" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7924" daytime="17:54" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7925" daytime="17:56" number="20" order="20" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1431" daytime="17:57" gender="F" number="24" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1432" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6200" />
                    <RANKING order="2" place="2" resultid="3905" />
                    <RANKING order="3" place="3" resultid="2630" />
                    <RANKING order="4" place="4" resultid="3032" />
                    <RANKING order="5" place="5" resultid="5842" />
                    <RANKING order="6" place="6" resultid="1989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6352" />
                    <RANKING order="2" place="2" resultid="3845" />
                    <RANKING order="3" place="3" resultid="4733" />
                    <RANKING order="4" place="4" resultid="2923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5585" />
                    <RANKING order="2" place="2" resultid="5942" />
                    <RANKING order="3" place="3" resultid="6035" />
                    <RANKING order="4" place="4" resultid="5932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1435" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2930" />
                    <RANKING order="2" place="2" resultid="6204" />
                    <RANKING order="3" place="3" resultid="5282" />
                    <RANKING order="4" place="4" resultid="4022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1436" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5032" />
                    <RANKING order="2" place="2" resultid="5485" />
                    <RANKING order="3" place="3" resultid="3643" />
                    <RANKING order="4" place="4" resultid="2949" />
                    <RANKING order="5" place="5" resultid="6385" />
                    <RANKING order="6" place="6" resultid="6460" />
                    <RANKING order="7" place="-1" resultid="3750" />
                    <RANKING order="8" place="-1" resultid="3875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1437" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4370" />
                    <RANKING order="2" place="2" resultid="4653" />
                    <RANKING order="3" place="3" resultid="3219" />
                    <RANKING order="4" place="-1" resultid="4415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1438" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2139" />
                    <RANKING order="2" place="2" resultid="3040" />
                    <RANKING order="3" place="3" resultid="4989" />
                    <RANKING order="4" place="4" resultid="3599" />
                    <RANKING order="5" place="-1" resultid="4557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1439" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3399" />
                    <RANKING order="2" place="2" resultid="1981" />
                    <RANKING order="3" place="3" resultid="2009" />
                    <RANKING order="4" place="-1" resultid="2533" />
                    <RANKING order="5" place="-1" resultid="3144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1440" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4344" />
                    <RANKING order="2" place="2" resultid="6317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1441" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4056" />
                    <RANKING order="2" place="2" resultid="4674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5261" />
                    <RANKING order="2" place="-1" resultid="6347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1444" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1446" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7926" daytime="17:57" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7927" daytime="18:01" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7928" daytime="18:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7929" daytime="18:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7930" daytime="18:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7931" daytime="18:10" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1447" daytime="18:13" gender="M" number="25" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1448" agemax="24" agemin="20" name="Kategoria 0" />
                <AGEGROUP agegroupid="1449" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6140" />
                    <RANKING order="2" place="2" resultid="6330" />
                    <RANKING order="3" place="3" resultid="6279" />
                    <RANKING order="4" place="4" resultid="5143" />
                    <RANKING order="5" place="5" resultid="2589" />
                    <RANKING order="6" place="6" resultid="2076" />
                    <RANKING order="7" place="7" resultid="5118" />
                    <RANKING order="8" place="-1" resultid="2278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5603" />
                    <RANKING order="2" place="2" resultid="3239" />
                    <RANKING order="3" place="3" resultid="4061" />
                    <RANKING order="4" place="4" resultid="5632" />
                    <RANKING order="5" place="-1" resultid="3742" />
                    <RANKING order="6" place="-1" resultid="4217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1451" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1902" />
                    <RANKING order="2" place="2" resultid="2786" />
                    <RANKING order="3" place="3" resultid="6334" />
                    <RANKING order="4" place="4" resultid="1916" />
                    <RANKING order="5" place="5" resultid="3760" />
                    <RANKING order="6" place="6" resultid="5920" />
                    <RANKING order="7" place="7" resultid="2989" />
                    <RANKING order="8" place="8" resultid="5305" />
                    <RANKING order="9" place="9" resultid="4766" />
                    <RANKING order="10" place="10" resultid="3852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1452" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4333" />
                    <RANKING order="2" place="2" resultid="4668" />
                    <RANKING order="3" place="3" resultid="3579" />
                    <RANKING order="4" place="4" resultid="5212" />
                    <RANKING order="5" place="5" resultid="2777" />
                    <RANKING order="6" place="6" resultid="6372" />
                    <RANKING order="7" place="7" resultid="2118" />
                    <RANKING order="8" place="-1" resultid="3364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1453" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4376" />
                    <RANKING order="2" place="2" resultid="5347" />
                    <RANKING order="3" place="3" resultid="6339" />
                    <RANKING order="4" place="4" resultid="5887" />
                    <RANKING order="5" place="5" resultid="3234" />
                    <RANKING order="6" place="6" resultid="6060" />
                    <RANKING order="7" place="7" resultid="5710" />
                    <RANKING order="8" place="-1" resultid="2177" />
                    <RANKING order="9" place="-1" resultid="2857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1454" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4038" />
                    <RANKING order="2" place="2" resultid="4473" />
                    <RANKING order="3" place="3" resultid="3347" />
                    <RANKING order="4" place="4" resultid="4662" />
                    <RANKING order="5" place="5" resultid="2358" />
                    <RANKING order="6" place="6" resultid="5478" />
                    <RANKING order="7" place="7" resultid="2252" />
                    <RANKING order="8" place="8" resultid="3228" />
                    <RANKING order="9" place="9" resultid="4337" />
                    <RANKING order="10" place="10" resultid="5320" />
                    <RANKING order="11" place="-1" resultid="3833" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1455" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6009" />
                    <RANKING order="2" place="2" resultid="2539" />
                    <RANKING order="3" place="3" resultid="3319" />
                    <RANKING order="4" place="4" resultid="2625" />
                    <RANKING order="5" place="5" resultid="5523" />
                    <RANKING order="6" place="6" resultid="5427" />
                    <RANKING order="7" place="7" resultid="3205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1456" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2654" />
                    <RANKING order="2" place="2" resultid="4980" />
                    <RANKING order="3" place="3" resultid="2812" />
                    <RANKING order="4" place="4" resultid="3410" />
                    <RANKING order="5" place="5" resultid="5516" />
                    <RANKING order="6" place="6" resultid="4449" />
                    <RANKING order="7" place="7" resultid="5611" />
                    <RANKING order="8" place="-1" resultid="2672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1457" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3440" />
                    <RANKING order="2" place="2" resultid="4282" />
                    <RANKING order="3" place="3" resultid="5510" />
                    <RANKING order="4" place="4" resultid="3294" />
                    <RANKING order="5" place="5" resultid="3414" />
                    <RANKING order="6" place="6" resultid="3153" />
                    <RANKING order="7" place="-1" resultid="5618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1458" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3556" />
                    <RANKING order="2" place="2" resultid="6236" />
                    <RANKING order="3" place="3" resultid="2747" />
                    <RANKING order="4" place="-1" resultid="3795" />
                    <RANKING order="5" place="-1" resultid="5625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1460" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2665" />
                    <RANKING order="2" place="2" resultid="2015" />
                    <RANKING order="3" place="3" resultid="1958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1461" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1462" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7932" daytime="18:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7933" daytime="18:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7934" daytime="18:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7935" daytime="18:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7936" daytime="18:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7937" daytime="18:27" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7938" daytime="18:29" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7939" daytime="18:32" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7940" daytime="18:34" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7941" daytime="18:36" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7942" daytime="18:37" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1463" daytime="18:40" gender="F" number="26" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1464" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2573" />
                    <RANKING order="2" place="2" resultid="5152" />
                    <RANKING order="3" place="3" resultid="3910" />
                    <RANKING order="4" place="4" resultid="2609" />
                    <RANKING order="5" place="5" resultid="3781" />
                    <RANKING order="6" place="6" resultid="1972" />
                    <RANKING order="7" place="7" resultid="6257" />
                    <RANKING order="8" place="8" resultid="5579" />
                    <RANKING order="9" place="9" resultid="5111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4050" />
                    <RANKING order="2" place="2" resultid="6353" />
                    <RANKING order="3" place="3" resultid="4678" />
                    <RANKING order="4" place="4" resultid="6024" />
                    <RANKING order="5" place="5" resultid="4412" />
                    <RANKING order="6" place="6" resultid="5237" />
                    <RANKING order="7" place="7" resultid="3128" />
                    <RANKING order="8" place="8" resultid="5363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1466" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2274" />
                    <RANKING order="2" place="2" resultid="5876" />
                    <RANKING order="3" place="3" resultid="4790" />
                    <RANKING order="4" place="4" resultid="4743" />
                    <RANKING order="5" place="5" resultid="5943" />
                    <RANKING order="6" place="6" resultid="4030" />
                    <RANKING order="7" place="7" resultid="6016" />
                    <RANKING order="8" place="8" resultid="3685" />
                    <RANKING order="9" place="-1" resultid="5784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1941" />
                    <RANKING order="2" place="2" resultid="3697" />
                    <RANKING order="3" place="3" resultid="2958" />
                    <RANKING order="4" place="4" resultid="5283" />
                    <RANKING order="5" place="5" resultid="5902" />
                    <RANKING order="6" place="6" resultid="4023" />
                    <RANKING order="7" place="7" resultid="3861" />
                    <RANKING order="8" place="-1" resultid="3490" />
                    <RANKING order="9" place="-1" resultid="5766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1468" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4308" />
                    <RANKING order="2" place="2" resultid="6220" />
                    <RANKING order="3" place="3" resultid="6130" />
                    <RANKING order="4" place="-1" resultid="4755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1469" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3106" />
                    <RANKING order="2" place="2" resultid="6322" />
                    <RANKING order="3" place="3" resultid="4148" />
                    <RANKING order="4" place="4" resultid="6073" />
                    <RANKING order="5" place="5" resultid="3220" />
                    <RANKING order="6" place="6" resultid="4654" />
                    <RANKING order="7" place="7" resultid="2373" />
                    <RANKING order="8" place="8" resultid="4416" />
                    <RANKING order="9" place="-1" resultid="5373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1470" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5180" />
                    <RANKING order="2" place="2" resultid="3938" />
                    <RANKING order="3" place="3" resultid="6366" />
                    <RANKING order="4" place="4" resultid="2267" />
                    <RANKING order="5" place="5" resultid="4565" />
                    <RANKING order="6" place="6" resultid="3135" />
                    <RANKING order="7" place="7" resultid="2764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1471" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2131" />
                    <RANKING order="2" place="2" resultid="2258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1472" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5503" />
                    <RANKING order="2" place="2" resultid="4287" />
                    <RANKING order="3" place="3" resultid="5390" />
                    <RANKING order="4" place="-1" resultid="5008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1473" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5395" />
                    <RANKING order="2" place="2" resultid="3825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1474" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1475" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1476" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1477" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1478" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7943" daytime="18:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7944" daytime="18:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7945" daytime="18:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7946" daytime="18:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7947" daytime="19:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7948" daytime="19:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7949" daytime="19:08" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7950" daytime="19:12" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7951" daytime="19:15" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1479" daytime="19:19" gender="M" number="27" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1480" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3566" />
                    <RANKING order="2" place="2" resultid="6215" />
                    <RANKING order="3" place="3" resultid="4760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5138" />
                    <RANKING order="2" place="2" resultid="5957" />
                    <RANKING order="3" place="3" resultid="5827" />
                    <RANKING order="4" place="4" resultid="4076" />
                    <RANKING order="5" place="5" resultid="3839" />
                    <RANKING order="6" place="6" resultid="3899" />
                    <RANKING order="7" place="7" resultid="5434" />
                    <RANKING order="8" place="8" resultid="3691" />
                    <RANKING order="9" place="-1" resultid="5404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2071" />
                    <RANKING order="2" place="2" resultid="3242" />
                    <RANKING order="3" place="3" resultid="5821" />
                    <RANKING order="4" place="4" resultid="3584" />
                    <RANKING order="5" place="5" resultid="4157" />
                    <RANKING order="6" place="6" resultid="5633" />
                    <RANKING order="7" place="7" resultid="4193" />
                    <RANKING order="8" place="8" resultid="2392" />
                    <RANKING order="9" place="9" resultid="5245" />
                    <RANKING order="10" place="10" resultid="5299" />
                    <RANKING order="11" place="-1" resultid="1994" />
                    <RANKING order="12" place="-1" resultid="3743" />
                    <RANKING order="13" place="-1" resultid="4082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2311" />
                    <RANKING order="2" place="2" resultid="6053" />
                    <RANKING order="3" place="3" resultid="5557" />
                    <RANKING order="4" place="4" resultid="3112" />
                    <RANKING order="5" place="5" resultid="2881" />
                    <RANKING order="6" place="6" resultid="5400" />
                    <RANKING order="7" place="7" resultid="2399" />
                    <RANKING order="8" place="8" resultid="2968" />
                    <RANKING order="9" place="9" resultid="3761" />
                    <RANKING order="10" place="10" resultid="5146" />
                    <RANKING order="11" place="11" resultid="5542" />
                    <RANKING order="12" place="12" resultid="2976" />
                    <RANKING order="13" place="13" resultid="1950" />
                    <RANKING order="14" place="14" resultid="3056" />
                    <RANKING order="15" place="15" resultid="4203" />
                    <RANKING order="16" place="16" resultid="5982" />
                    <RANKING order="17" place="17" resultid="2303" />
                    <RANKING order="18" place="18" resultid="3167" />
                    <RANKING order="19" place="19" resultid="5438" />
                    <RANKING order="20" place="20" resultid="3122" />
                    <RANKING order="21" place="21" resultid="5697" />
                    <RANKING order="22" place="22" resultid="4767" />
                    <RANKING order="23" place="23" resultid="3672" />
                    <RANKING order="24" place="-1" resultid="2918" />
                    <RANKING order="25" place="-1" resultid="3704" />
                    <RANKING order="26" place="-1" resultid="3949" />
                    <RANKING order="27" place="-1" resultid="4708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1484" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5419" />
                    <RANKING order="2" place="2" resultid="6178" />
                    <RANKING order="3" place="3" resultid="3331" />
                    <RANKING order="4" place="4" resultid="5192" />
                    <RANKING order="5" place="5" resultid="2778" />
                    <RANKING order="6" place="6" resultid="6301" />
                    <RANKING order="7" place="7" resultid="6188" />
                    <RANKING order="8" place="8" resultid="4432" />
                    <RANKING order="9" place="9" resultid="6380" />
                    <RANKING order="10" place="10" resultid="6208" />
                    <RANKING order="11" place="11" resultid="3469" />
                    <RANKING order="12" place="12" resultid="4750" />
                    <RANKING order="13" place="13" resultid="3475" />
                    <RANKING order="14" place="14" resultid="5703" />
                    <RANKING order="15" place="-1" resultid="3547" />
                    <RANKING order="16" place="-1" resultid="2598" />
                    <RANKING order="17" place="-1" resultid="5738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1485" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6195" />
                    <RANKING order="2" place="2" resultid="3637" />
                    <RANKING order="3" place="3" resultid="2181" />
                    <RANKING order="4" place="4" resultid="5888" />
                    <RANKING order="5" place="5" resultid="2348" />
                    <RANKING order="6" place="6" resultid="5531" />
                    <RANKING order="7" place="7" resultid="2695" />
                    <RANKING order="8" place="8" resultid="2041" />
                    <RANKING order="9" place="9" resultid="3920" />
                    <RANKING order="10" place="10" resultid="6229" />
                    <RANKING order="11" place="11" resultid="5716" />
                    <RANKING order="12" place="-1" resultid="3482" />
                    <RANKING order="13" place="-1" resultid="5126" />
                    <RANKING order="14" place="-1" resultid="6061" />
                    <RANKING order="15" place="-1" resultid="2368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1486" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3256" />
                    <RANKING order="2" place="2" resultid="1922" />
                    <RANKING order="3" place="3" resultid="3650" />
                    <RANKING order="4" place="4" resultid="6040" />
                    <RANKING order="5" place="5" resultid="3212" />
                    <RANKING order="6" place="6" resultid="3171" />
                    <RANKING order="7" place="7" resultid="4727" />
                    <RANKING order="8" place="8" resultid="5269" />
                    <RANKING order="9" place="9" resultid="5289" />
                    <RANKING order="10" place="-1" resultid="2547" />
                    <RANKING order="11" place="-1" resultid="2830" />
                    <RANKING order="12" place="-1" resultid="5294" />
                    <RANKING order="13" place="-1" resultid="5895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1487" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5046" />
                    <RANKING order="2" place="2" resultid="3610" />
                    <RANKING order="3" place="3" resultid="4466" />
                    <RANKING order="4" place="4" resultid="6288" />
                    <RANKING order="5" place="5" resultid="4488" />
                    <RANKING order="6" place="6" resultid="6121" />
                    <RANKING order="7" place="7" resultid="5198" />
                    <RANKING order="8" place="8" resultid="2754" />
                    <RANKING order="9" place="-1" resultid="1867" />
                    <RANKING order="10" place="-1" resultid="3049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1488" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3515" />
                    <RANKING order="2" place="2" resultid="4613" />
                    <RANKING order="3" place="3" resultid="3450" />
                    <RANKING order="4" place="4" resultid="5869" />
                    <RANKING order="5" place="5" resultid="4691" />
                    <RANKING order="6" place="-1" resultid="2673" />
                    <RANKING order="7" place="-1" resultid="4543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1489" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2707" />
                    <RANKING order="2" place="2" resultid="3815" />
                    <RANKING order="3" place="3" resultid="3441" />
                    <RANKING order="4" place="4" resultid="5027" />
                    <RANKING order="5" place="5" resultid="2407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1490" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4316" />
                    <RANKING order="2" place="2" resultid="3796" />
                    <RANKING order="3" place="-1" resultid="4440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1491" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1492" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2016" />
                    <RANKING order="2" place="2" resultid="5166" />
                    <RANKING order="3" place="3" resultid="1959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1494" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7952" daytime="19:19" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7953" daytime="19:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7954" daytime="19:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7955" daytime="19:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7956" daytime="19:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7957" daytime="19:42" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7958" daytime="19:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7959" daytime="19:49" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7960" daytime="19:52" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7961" daytime="19:56" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7962" daytime="19:59" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7963" daytime="20:02" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7964" daytime="20:05" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7965" daytime="20:08" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7966" daytime="20:11" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7967" daytime="20:14" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1495" daytime="20:18" gender="F" number="28" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1559" agemax="96" agemin="80" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="1560" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1561" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3002" />
                    <RANKING order="2" place="2" resultid="6077" />
                    <RANKING order="3" place="3" resultid="3972" />
                    <RANKING order="4" place="4" resultid="5986" />
                    <RANKING order="5" place="5" resultid="6454" />
                    <RANKING order="6" place="6" resultid="3089" />
                    <RANKING order="7" place="-1" resultid="4117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1562" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5053" />
                    <RANKING order="2" place="-1" resultid="5798" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1563" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3986" />
                    <RANKING order="2" place="2" resultid="4635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1564" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1565" agemax="400" agemin="280" name="Kategoria F" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7968" daytime="20:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7969" daytime="20:21" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1511" daytime="20:25" gender="M" number="29" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1566" agemax="96" agemin="80" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="1567" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6448" />
                    <RANKING order="2" place="-1" resultid="6410" />
                    <RANKING order="3" place="-1" resultid="8772" />
                    <RANKING order="4" place="-1" resultid="2078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1568" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5753" />
                    <RANKING order="2" place="2" resultid="4119" />
                    <RANKING order="3" place="3" resultid="3270" />
                    <RANKING order="4" place="4" resultid="4813" />
                    <RANKING order="5" place="5" resultid="3981" />
                    <RANKING order="6" place="6" resultid="4243" />
                    <RANKING order="7" place="7" resultid="4244" />
                    <RANKING order="8" place="8" resultid="6455" />
                    <RANKING order="9" place="9" resultid="4246" />
                    <RANKING order="10" place="-1" resultid="2337" />
                    <RANKING order="11" place="-1" resultid="3087" />
                    <RANKING order="12" place="-1" resultid="3708" />
                    <RANKING order="13" place="-1" resultid="4121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1569" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5985" />
                    <RANKING order="2" place="2" resultid="2887" />
                    <RANKING order="3" place="3" resultid="3983" />
                    <RANKING order="4" place="4" resultid="2097" />
                    <RANKING order="5" place="5" resultid="5223" />
                    <RANKING order="6" place="6" resultid="3003" />
                    <RANKING order="7" place="7" resultid="3272" />
                    <RANKING order="8" place="8" resultid="6082" />
                    <RANKING order="9" place="9" resultid="4815" />
                    <RANKING order="10" place="10" resultid="5718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2190" />
                    <RANKING order="2" place="2" resultid="5545" />
                    <RANKING order="3" place="3" resultid="4517" />
                    <RANKING order="4" place="4" resultid="3984" />
                    <RANKING order="5" place="-1" resultid="2378" />
                    <RANKING order="6" place="-1" resultid="3500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1571" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5055" />
                    <RANKING order="2" place="2" resultid="4385" />
                    <RANKING order="3" place="3" resultid="4515" />
                    <RANKING order="4" place="-1" resultid="4634" />
                    <RANKING order="5" place="-1" resultid="5664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1572" agemax="400" agemin="280" name="Kategoria F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4384" />
                    <RANKING order="2" place="-1" resultid="5666" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7970" daytime="20:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7971" daytime="20:29" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7972" daytime="20:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7973" daytime="20:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7974" daytime="20:37" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1527" daytime="20:40" gender="F" number="30" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1528" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1529" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3846" />
                    <RANKING order="2" place="2" resultid="3808" />
                    <RANKING order="3" place="3" resultid="5312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1530" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5103" />
                    <RANKING order="2" place="2" resultid="4031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1531" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1943" />
                    <RANKING order="2" place="2" resultid="3386" />
                    <RANKING order="3" place="-1" resultid="3619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1532" agemax="44" agemin="40" name="Kategoria D" />
                <AGEGROUP agegroupid="1533" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5174" />
                    <RANKING order="2" place="2" resultid="6074" />
                    <RANKING order="3" place="3" resultid="4149" />
                    <RANKING order="4" place="-1" resultid="2849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1534" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3041" />
                    <RANKING order="2" place="2" resultid="4558" />
                    <RANKING order="3" place="3" resultid="3136" />
                    <RANKING order="4" place="-1" resultid="4628" />
                    <RANKING order="5" place="-1" resultid="4685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1535" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3929" />
                    <RANKING order="2" place="2" resultid="2534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1536" agemax="64" agemin="60" name="Kategoria H" />
                <AGEGROUP agegroupid="1537" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="1538" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="1539" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1540" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1541" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1542" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8802" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8803" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8804" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1543" daytime="21:09" gender="M" number="31" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1544" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5160" />
                    <RANKING order="2" place="2" resultid="3661" />
                    <RANKING order="3" place="-1" resultid="2582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1545" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2053" />
                    <RANKING order="2" place="2" resultid="2279" />
                    <RANKING order="3" place="3" resultid="4778" />
                    <RANKING order="4" place="4" resultid="2030" />
                    <RANKING order="5" place="-1" resultid="2590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1546" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5604" />
                    <RANKING order="2" place="2" resultid="1909" />
                    <RANKING order="3" place="3" resultid="6045" />
                    <RANKING order="4" place="4" resultid="4230" />
                    <RANKING order="5" place="5" resultid="5591" />
                    <RANKING order="6" place="-1" resultid="4158" />
                    <RANKING order="7" place="-1" resultid="4804" />
                    <RANKING order="8" place="-1" resultid="5779" />
                    <RANKING order="9" place="-1" resultid="4167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1547" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2312" />
                    <RANKING order="2" place="2" resultid="5921" />
                    <RANKING order="3" place="3" resultid="5204" />
                    <RANKING order="4" place="4" resultid="2840" />
                    <RANKING order="5" place="-1" resultid="1917" />
                    <RANKING order="6" place="-1" resultid="2865" />
                    <RANKING order="7" place="-1" resultid="2873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1548" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3856" />
                    <RANKING order="2" place="2" resultid="6373" />
                    <RANKING order="3" place="3" resultid="5220" />
                    <RANKING order="4" place="4" resultid="2732" />
                    <RANKING order="5" place="-1" resultid="3666" />
                    <RANKING order="6" place="-1" resultid="5745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1549" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3656" />
                    <RANKING order="2" place="2" resultid="3018" />
                    <RANKING order="3" place="-1" resultid="6196" />
                    <RANKING order="4" place="-1" resultid="6402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1550" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2604" />
                    <RANKING order="2" place="2" resultid="5019" />
                    <RANKING order="3" place="3" resultid="3184" />
                    <RANKING order="4" place="-1" resultid="2831" />
                    <RANKING order="5" place="-1" resultid="5321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1551" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2556" />
                    <RANKING order="2" place="2" resultid="5524" />
                    <RANKING order="3" place="3" resultid="4137" />
                    <RANKING order="4" place="4" resultid="3176" />
                    <RANKING order="5" place="-1" resultid="3050" />
                    <RANKING order="6" place="-1" resultid="6122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1552" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4424" />
                    <RANKING order="2" place="2" resultid="4479" />
                    <RANKING order="3" place="3" resultid="2813" />
                    <RANKING order="4" place="4" resultid="3451" />
                    <RANKING order="5" place="5" resultid="2655" />
                    <RANKING order="6" place="6" resultid="5651" />
                    <RANKING order="7" place="7" resultid="5658" />
                    <RANKING order="8" place="8" resultid="3191" />
                    <RANKING order="9" place="9" resultid="3460" />
                    <RANKING order="10" place="-1" resultid="4981" />
                    <RANKING order="11" place="-1" resultid="4586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1553" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2242" />
                    <RANKING order="2" place="2" resultid="3816" />
                    <RANKING order="3" place="3" resultid="3295" />
                    <RANKING order="4" place="4" resultid="3305" />
                    <RANKING order="5" place="-1" resultid="2739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1554" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1555" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1556" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1557" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1558" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8806" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8807" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8808" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8809" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8810" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8811" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8812" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="8925" />
            <JUDGE officialid="8910" />
            <JUDGE officialid="8924" />
            <JUDGE officialid="8926" />
            <JUDGE officialid="8906" />
            <JUDGE officialid="8919" />
            <JUDGE officialid="8923" />
            <JUDGE officialid="8909" />
            <JUDGE officialid="8921" />
            <JUDGE officialid="8914" />
            <JUDGE officialid="8915" />
            <JUDGE officialid="8918" />
            <JUDGE officialid="8922" />
            <JUDGE officialid="8917" />
            <JUDGE officialid="8920" />
            <JUDGE officialid="8928" />
            <JUDGE officialid="8912" />
            <JUDGE officialid="8916" />
            <JUDGE officialid="8916" />
            <JUDGE officialid="8908" />
            <JUDGE officialid="8908" />
            <JUDGE officialid="8911" />
            <JUDGE officialid="8911" />
            <JUDGE officialid="8913" />
            <JUDGE officialid="8927" />
            <JUDGE officialid="8905" />
            <JUDGE officialid="8904" />
            <JUDGE officialid="8903" />
            <JUDGE officialid="8907" />
            <JUDGE officialid="8941" />
            <JUDGE officialid="8901" />
            <JUDGE officialid="8902" />
          </JUDGES>
        </SESSION>
        <SESSION date="2013-11-17" daytime="09:00" name="MP Masters BLOK IV" number="4" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1574" daytime="09:00" gender="F" number="32" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1576" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3033" />
                    <RANKING order="2" place="2" resultid="2218" />
                    <RANKING order="3" place="3" resultid="3953" />
                    <RANKING order="4" place="4" resultid="3912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1577" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6025" />
                    <RANKING order="2" place="2" resultid="5571" />
                    <RANKING order="3" place="3" resultid="5238" />
                    <RANKING order="4" place="4" resultid="5313" />
                    <RANKING order="5" place="-1" resultid="3964" />
                    <RANKING order="6" place="-1" resultid="4797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1578" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5445" />
                    <RANKING order="2" place="2" resultid="5877" />
                    <RANKING order="3" place="3" resultid="4744" />
                    <RANKING order="4" place="4" resultid="5104" />
                    <RANKING order="5" place="5" resultid="6017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1579" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2938" />
                    <RANKING order="2" place="2" resultid="3387" />
                    <RANKING order="3" place="-1" resultid="5767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1580" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5039" />
                    <RANKING order="2" place="2" resultid="4309" />
                    <RANKING order="3" place="-1" resultid="6104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1581" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5175" />
                    <RANKING order="2" place="2" resultid="2850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1582" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4990" />
                    <RANKING order="2" place="2" resultid="3939" />
                    <RANKING order="3" place="3" resultid="4622" />
                    <RANKING order="4" place="4" resultid="3137" />
                    <RANKING order="5" place="-1" resultid="4629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2132" />
                    <RANKING order="2" place="2" resultid="3930" />
                    <RANKING order="3" place="3" resultid="4606" />
                    <RANKING order="4" place="4" resultid="2259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1584" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="1586" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1587" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1588" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1589" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1590" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7987" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7988" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7989" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7990" daytime="09:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7991" daytime="09:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1591" daytime="09:12" gender="M" number="33" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1592" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3567" />
                    <RANKING order="2" place="2" resultid="2583" />
                    <RANKING order="3" place="3" resultid="6395" />
                    <RANKING order="4" place="4" resultid="5752" />
                    <RANKING order="5" place="5" resultid="2564" />
                    <RANKING order="6" place="-1" resultid="2226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1593" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5729" />
                    <RANKING order="2" place="2" resultid="5958" />
                    <RANKING order="3" place="3" resultid="5139" />
                    <RANKING order="4" place="4" resultid="6280" />
                    <RANKING order="5" place="5" resultid="4077" />
                    <RANKING order="6" place="6" resultid="4514" />
                    <RANKING order="7" place="-1" resultid="2637" />
                    <RANKING order="8" place="-1" resultid="4067" />
                    <RANKING order="9" place="-1" resultid="5748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1594" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1874" />
                    <RANKING order="2" place="2" resultid="1910" />
                    <RANKING order="3" place="3" resultid="3248" />
                    <RANKING order="4" place="4" resultid="4231" />
                    <RANKING order="5" place="5" resultid="4194" />
                    <RANKING order="6" place="6" resultid="4083" />
                    <RANKING order="7" place="7" resultid="5822" />
                    <RANKING order="8" place="8" resultid="2393" />
                    <RANKING order="9" place="9" resultid="4719" />
                    <RANKING order="10" place="10" resultid="5592" />
                    <RANKING order="11" place="-1" resultid="4183" />
                    <RANKING order="12" place="-1" resultid="5780" />
                    <RANKING order="13" place="-1" resultid="3499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1595" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5558" />
                    <RANKING order="2" place="2" resultid="2313" />
                    <RANKING order="3" place="3" resultid="6054" />
                    <RANKING order="4" place="4" resultid="2919" />
                    <RANKING order="5" place="5" resultid="6068" />
                    <RANKING order="6" place="6" resultid="5205" />
                    <RANKING order="7" place="7" resultid="5922" />
                    <RANKING order="8" place="8" resultid="2972" />
                    <RANKING order="9" place="9" resultid="2400" />
                    <RANKING order="10" place="10" resultid="2304" />
                    <RANKING order="11" place="11" resultid="2874" />
                    <RANKING order="12" place="-1" resultid="1929" />
                    <RANKING order="13" place="-1" resultid="3673" />
                    <RANKING order="14" place="-1" resultid="4210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1596" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2796" />
                    <RANKING order="2" place="2" resultid="5420" />
                    <RANKING order="3" place="3" resultid="3332" />
                    <RANKING order="4" place="4" resultid="6302" />
                    <RANKING order="5" place="5" resultid="3857" />
                    <RANKING order="6" place="6" resultid="4322" />
                    <RANKING order="7" place="7" resultid="2779" />
                    <RANKING order="8" place="8" resultid="4433" />
                    <RANKING order="9" place="9" resultid="6030" />
                    <RANKING order="10" place="-1" resultid="2733" />
                    <RANKING order="11" place="-1" resultid="5221" />
                    <RANKING order="12" place="-1" resultid="5746" />
                    <RANKING order="13" place="-1" resultid="6179" />
                    <RANKING order="14" place="-1" resultid="4593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1597" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5532" />
                    <RANKING order="2" place="2" resultid="2858" />
                    <RANKING order="3" place="3" resultid="5276" />
                    <RANKING order="4" place="-1" resultid="3097" />
                    <RANKING order="5" place="-1" resultid="6403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1923" />
                    <RANKING order="2" place="2" resultid="2548" />
                    <RANKING order="3" place="3" resultid="3834" />
                    <RANKING order="4" place="4" resultid="2832" />
                    <RANKING order="5" place="5" resultid="3213" />
                    <RANKING order="6" place="6" resultid="5020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6010" />
                    <RANKING order="2" place="2" resultid="5950" />
                    <RANKING order="3" place="3" resultid="4467" />
                    <RANKING order="4" place="4" resultid="2557" />
                    <RANKING order="5" place="5" resultid="2755" />
                    <RANKING order="6" place="6" resultid="3199" />
                    <RANKING order="7" place="-1" resultid="3051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5652" />
                    <RANKING order="2" place="2" resultid="4480" />
                    <RANKING order="3" place="3" resultid="4425" />
                    <RANKING order="4" place="4" resultid="5659" />
                    <RANKING order="5" place="5" resultid="4587" />
                    <RANKING order="6" place="6" resultid="3192" />
                    <RANKING order="7" place="-1" resultid="5870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6225" />
                    <RANKING order="2" place="2" resultid="2682" />
                    <RANKING order="3" place="3" resultid="2243" />
                    <RANKING order="4" place="4" resultid="5028" />
                    <RANKING order="5" place="5" resultid="3817" />
                    <RANKING order="6" place="6" resultid="2740" />
                    <RANKING order="7" place="7" resultid="1896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6254" />
                    <RANKING order="2" place="2" resultid="2748" />
                    <RANKING order="3" place="3" resultid="4574" />
                    <RANKING order="4" place="4" resultid="3557" />
                    <RANKING order="5" place="-1" resultid="6238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1881" />
                    <RANKING order="2" place="2" resultid="5254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1606" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7992" daytime="09:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7993" daytime="09:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7994" daytime="09:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7995" daytime="09:21" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7996" daytime="09:23" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7997" daytime="09:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7998" daytime="09:28" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7999" daytime="09:30" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8000" daytime="09:32" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8001" daytime="09:34" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="8002" daytime="09:36" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="8003" daytime="09:37" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1607" daytime="09:40" gender="F" number="34" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1608" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2631" />
                    <RANKING order="2" place="2" resultid="3957" />
                    <RANKING order="3" place="3" resultid="1973" />
                    <RANKING order="4" place="4" resultid="5580" />
                    <RANKING order="5" place="5" resultid="1990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1609" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4734" />
                    <RANKING order="2" place="2" resultid="3847" />
                    <RANKING order="3" place="3" resultid="6354" />
                    <RANKING order="4" place="4" resultid="2924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1610" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5586" />
                    <RANKING order="2" place="2" resultid="3593" />
                    <RANKING order="3" place="3" resultid="5944" />
                    <RANKING order="4" place="4" resultid="6036" />
                    <RANKING order="5" place="5" resultid="4032" />
                    <RANKING order="6" place="6" resultid="5933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1611" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2931" />
                    <RANKING order="2" place="2" resultid="5284" />
                    <RANKING order="3" place="-1" resultid="4024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1612" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5033" />
                    <RANKING order="2" place="2" resultid="3644" />
                    <RANKING order="3" place="3" resultid="2950" />
                    <RANKING order="4" place="4" resultid="3751" />
                    <RANKING order="5" place="5" resultid="3876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1613" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4371" />
                    <RANKING order="2" place="2" resultid="3107" />
                    <RANKING order="3" place="3" resultid="4150" />
                    <RANKING order="4" place="4" resultid="4655" />
                    <RANKING order="5" place="5" resultid="3221" />
                    <RANKING order="6" place="6" resultid="6075" />
                    <RANKING order="7" place="7" resultid="4417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1614" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3042" />
                    <RANKING order="2" place="2" resultid="2268" />
                    <RANKING order="3" place="-1" resultid="2140" />
                    <RANKING order="4" place="-1" resultid="3600" />
                    <RANKING order="5" place="-1" resultid="4559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1615" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1982" />
                    <RANKING order="2" place="2" resultid="2010" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1616" agemax="64" agemin="60" name="Kategoria H" />
                <AGEGROUP agegroupid="1617" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5396" />
                    <RANKING order="2" place="2" resultid="4675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4293" />
                    <RANKING order="2" place="2" resultid="5262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1620" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1621" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1622" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8004" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8005" daytime="09:47" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8006" daytime="09:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8007" daytime="09:57" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8008" daytime="10:01" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8009" daytime="10:04" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1623" daytime="10:08" gender="M" number="35" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1624" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1625" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6331" />
                    <RANKING order="2" place="2" resultid="2591" />
                    <RANKING order="3" place="3" resultid="2280" />
                    <RANKING order="4" place="4" resultid="2031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1626" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5605" />
                    <RANKING order="2" place="2" resultid="4062" />
                    <RANKING order="3" place="3" resultid="5634" />
                    <RANKING order="4" place="4" resultid="4232" />
                    <RANKING order="5" place="5" resultid="4168" />
                    <RANKING order="6" place="-1" resultid="4159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1627" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1903" />
                    <RANKING order="2" place="2" resultid="2787" />
                    <RANKING order="3" place="3" resultid="6335" />
                    <RANKING order="4" place="4" resultid="2866" />
                    <RANKING order="5" place="5" resultid="4709" />
                    <RANKING order="6" place="6" resultid="5923" />
                    <RANKING order="7" place="7" resultid="1918" />
                    <RANKING order="8" place="8" resultid="4768" />
                    <RANKING order="9" place="-1" resultid="2841" />
                    <RANKING order="10" place="-1" resultid="3113" />
                    <RANKING order="11" place="-1" resultid="4204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1628" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4334" />
                    <RANKING order="2" place="2" resultid="4669" />
                    <RANKING order="3" place="3" resultid="3580" />
                    <RANKING order="4" place="4" resultid="5213" />
                    <RANKING order="5" place="5" resultid="6374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1629" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4377" />
                    <RANKING order="2" place="2" resultid="5348" />
                    <RANKING order="3" place="3" resultid="6340" />
                    <RANKING order="4" place="4" resultid="5889" />
                    <RANKING order="5" place="5" resultid="2349" />
                    <RANKING order="6" place="6" resultid="3235" />
                    <RANKING order="7" place="7" resultid="2859" />
                    <RANKING order="8" place="-1" resultid="2178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1630" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4039" />
                    <RANKING order="2" place="2" resultid="4474" />
                    <RANKING order="3" place="3" resultid="2549" />
                    <RANKING order="4" place="4" resultid="2833" />
                    <RANKING order="5" place="5" resultid="5479" />
                    <RANKING order="6" place="6" resultid="4338" />
                    <RANKING order="7" place="7" resultid="3185" />
                    <RANKING order="8" place="8" resultid="3214" />
                    <RANKING order="9" place="-1" resultid="3651" />
                    <RANKING order="10" place="-1" resultid="4663" />
                    <RANKING order="11" place="-1" resultid="5322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1631" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3320" />
                    <RANKING order="2" place="2" resultid="5047" />
                    <RANKING order="3" place="3" resultid="2626" />
                    <RANKING order="4" place="4" resultid="5525" />
                    <RANKING order="5" place="5" resultid="4489" />
                    <RANKING order="6" place="6" resultid="2641" />
                    <RANKING order="7" place="7" resultid="3177" />
                    <RANKING order="8" place="8" resultid="3206" />
                    <RANKING order="9" place="9" resultid="5428" />
                    <RANKING order="10" place="-1" resultid="4138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1632" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3452" />
                    <RANKING order="2" place="2" resultid="2814" />
                    <RANKING order="3" place="3" resultid="2656" />
                    <RANKING order="4" place="4" resultid="4982" />
                    <RANKING order="5" place="5" resultid="4450" />
                    <RANKING order="6" place="6" resultid="5612" />
                    <RANKING order="7" place="-1" resultid="3411" />
                    <RANKING order="8" place="-1" resultid="2767" />
                    <RANKING order="9" place="-1" resultid="5517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2708" />
                    <RANKING order="2" place="2" resultid="3442" />
                    <RANKING order="3" place="3" resultid="5511" />
                    <RANKING order="4" place="4" resultid="4283" />
                    <RANKING order="5" place="5" resultid="3296" />
                    <RANKING order="6" place="6" resultid="3415" />
                    <RANKING order="7" place="7" resultid="3306" />
                    <RANKING order="8" place="8" resultid="3154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3558" />
                    <RANKING order="2" place="2" resultid="6239" />
                    <RANKING order="3" place="-1" resultid="5626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4458" />
                    <RANKING order="2" place="-1" resultid="5255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2017" />
                    <RANKING order="2" place="2" resultid="1960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1638" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8010" daytime="10:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8011" daytime="10:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8012" daytime="10:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8013" daytime="10:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8014" daytime="10:29" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8015" daytime="10:33" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8016" daytime="10:37" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8017" daytime="10:41" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8018" daytime="10:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8019" daytime="10:48" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1639" daytime="10:51" gender="F" number="36" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1640" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2574" />
                    <RANKING order="2" place="2" resultid="1974" />
                    <RANKING order="3" place="3" resultid="2219" />
                    <RANKING order="4" place="4" resultid="3782" />
                    <RANKING order="5" place="5" resultid="5112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1641" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5572" />
                    <RANKING order="2" place="2" resultid="3544" />
                    <RANKING order="3" place="3" resultid="3965" />
                    <RANKING order="4" place="4" resultid="3809" />
                    <RANKING order="5" place="5" resultid="6295" />
                    <RANKING order="6" place="-1" resultid="5368" />
                    <RANKING order="7" place="-1" resultid="5795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1642" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4045" />
                    <RANKING order="2" place="2" resultid="6165" />
                    <RANKING order="3" place="3" resultid="4745" />
                    <RANKING order="4" place="4" resultid="4100" />
                    <RANKING order="5" place="5" resultid="5934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1643" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5412" />
                    <RANKING order="2" place="2" resultid="2932" />
                    <RANKING order="3" place="3" resultid="2939" />
                    <RANKING order="4" place="4" resultid="5132" />
                    <RANKING order="5" place="5" resultid="5903" />
                    <RANKING order="6" place="6" resultid="3491" />
                    <RANKING order="7" place="-1" resultid="5768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1644" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4550" />
                    <RANKING order="2" place="2" resultid="2679" />
                    <RANKING order="3" place="3" resultid="2954" />
                    <RANKING order="4" place="4" resultid="4698" />
                    <RANKING order="5" place="5" resultid="3070" />
                    <RANKING order="6" place="6" resultid="2142" />
                    <RANKING order="7" place="7" resultid="3877" />
                    <RANKING order="8" place="-1" resultid="4756" />
                    <RANKING order="9" place="-1" resultid="6105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1645" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3714" />
                    <RANKING order="2" place="2" resultid="5374" />
                    <RANKING order="3" place="3" resultid="2851" />
                    <RANKING order="4" place="4" resultid="5490" />
                    <RANKING order="5" place="5" resultid="6323" />
                    <RANKING order="6" place="6" resultid="6782" />
                    <RANKING order="7" place="7" resultid="6468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1646" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4997" />
                    <RANKING order="2" place="2" resultid="3886" />
                    <RANKING order="3" place="3" resultid="4623" />
                    <RANKING order="4" place="4" resultid="6367" />
                    <RANKING order="5" place="5" resultid="5940" />
                    <RANKING order="6" place="6" resultid="2269" />
                    <RANKING order="7" place="7" resultid="2765" />
                    <RANKING order="8" place="-1" resultid="3419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1647" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2260" />
                    <RANKING order="2" place="2" resultid="3341" />
                    <RANKING order="3" place="3" resultid="3401" />
                    <RANKING order="4" place="4" resultid="3145" />
                    <RANKING order="5" place="-1" resultid="4607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1648" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4345" />
                    <RANKING order="2" place="2" resultid="5504" />
                    <RANKING order="3" place="3" resultid="3789" />
                    <RANKING order="4" place="4" resultid="3357" />
                    <RANKING order="5" place="5" resultid="5010" />
                    <RANKING order="6" place="6" resultid="3159" />
                    <RANKING order="7" place="-1" resultid="4598" />
                    <RANKING order="8" place="-1" resultid="6170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1649" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4327" />
                    <RANKING order="2" place="2" resultid="3826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4274" />
                    <RANKING order="2" place="2" resultid="5263" />
                    <RANKING order="3" place="-1" resultid="6346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3118" />
                    <RANKING order="2" place="2" resultid="2125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1653" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1654" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8020" daytime="10:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8021" daytime="10:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8022" daytime="10:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8023" daytime="10:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8024" daytime="11:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8025" daytime="11:01" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8026" daytime="11:03" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8027" daytime="11:04" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8028" daytime="11:06" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1655" daytime="11:08" gender="M" number="37" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1656" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5161" />
                    <RANKING order="2" place="2" resultid="2284" />
                    <RANKING order="3" place="2" resultid="6244" />
                    <RANKING order="4" place="4" resultid="3568" />
                    <RANKING order="5" place="5" resultid="2210" />
                    <RANKING order="6" place="6" resultid="2565" />
                    <RANKING order="7" place="7" resultid="2291" />
                    <RANKING order="8" place="-1" resultid="3538" />
                    <RANKING order="9" place="-1" resultid="5691" />
                    <RANKING order="10" place="-1" resultid="6216" />
                    <RANKING order="11" place="-1" resultid="6324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1657" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5359" />
                    <RANKING order="2" place="2" resultid="5818" />
                    <RANKING order="3" place="3" resultid="5384" />
                    <RANKING order="4" place="4" resultid="2025" />
                    <RANKING order="5" place="5" resultid="5811" />
                    <RANKING order="6" place="6" resultid="3252" />
                    <RANKING order="7" place="6" resultid="5814" />
                    <RANKING order="8" place="8" resultid="6281" />
                    <RANKING order="9" place="9" resultid="2592" />
                    <RANKING order="10" place="10" resultid="5355" />
                    <RANKING order="11" place="11" resultid="3736" />
                    <RANKING order="12" place="-1" resultid="2059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1658" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4772" />
                    <RANKING order="2" place="2" resultid="5967" />
                    <RANKING order="3" place="3" resultid="4088" />
                    <RANKING order="4" place="4" resultid="6046" />
                    <RANKING order="5" place="5" resultid="4188" />
                    <RANKING order="6" place="6" resultid="3679" />
                    <RANKING order="7" place="7" resultid="3060" />
                    <RANKING order="8" place="8" resultid="4720" />
                    <RANKING order="9" place="9" resultid="2332" />
                    <RANKING order="10" place="10" resultid="4169" />
                    <RANKING order="11" place="11" resultid="4173" />
                    <RANKING order="12" place="12" resultid="4218" />
                    <RANKING order="13" place="13" resultid="2759" />
                    <RANKING order="14" place="-1" resultid="2036" />
                    <RANKING order="15" place="-1" resultid="3530" />
                    <RANKING order="16" place="-1" resultid="4112" />
                    <RANKING order="17" place="-1" resultid="4198" />
                    <RANKING order="18" place="-1" resultid="5246" />
                    <RANKING order="19" place="-1" resultid="5597" />
                    <RANKING order="20" place="-1" resultid="4233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1659" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2867" />
                    <RANKING order="2" place="2" resultid="3339" />
                    <RANKING order="3" place="3" resultid="2882" />
                    <RANKING order="4" place="4" resultid="3351" />
                    <RANKING order="5" place="5" resultid="5543" />
                    <RANKING order="6" place="6" resultid="5790" />
                    <RANKING order="7" place="7" resultid="2986" />
                    <RANKING order="8" place="8" resultid="2788" />
                    <RANKING order="9" place="9" resultid="2323" />
                    <RANKING order="10" place="10" resultid="2875" />
                    <RANKING order="11" place="11" resultid="4105" />
                    <RANKING order="12" place="12" resultid="4205" />
                    <RANKING order="13" place="13" resultid="1951" />
                    <RANKING order="14" place="14" resultid="3705" />
                    <RANKING order="15" place="15" resultid="5914" />
                    <RANKING order="16" place="16" resultid="4769" />
                    <RANKING order="17" place="17" resultid="5439" />
                    <RANKING order="18" place="18" resultid="4785" />
                    <RANKING order="19" place="-1" resultid="2203" />
                    <RANKING order="20" place="-1" resultid="2842" />
                    <RANKING order="21" place="-1" resultid="6137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1660" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2797" />
                    <RANKING order="2" place="2" resultid="2717" />
                    <RANKING order="3" place="3" resultid="3667" />
                    <RANKING order="4" place="4" resultid="2992" />
                    <RANKING order="5" place="5" resultid="5214" />
                    <RANKING order="6" place="6" resultid="6361" />
                    <RANKING order="7" place="7" resultid="2734" />
                    <RANKING order="8" place="-1" resultid="3365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1661" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5127" />
                    <RANKING order="2" place="2" resultid="3870" />
                    <RANKING order="3" place="3" resultid="3019" />
                    <RANKING order="4" place="4" resultid="5533" />
                    <RANKING order="5" place="5" resultid="2171" />
                    <RANKING order="6" place="6" resultid="5379" />
                    <RANKING order="7" place="7" resultid="5711" />
                    <RANKING order="8" place="8" resultid="3390" />
                    <RANKING order="9" place="9" resultid="2633" />
                    <RANKING order="10" place="10" resultid="3394" />
                    <RANKING order="11" place="11" resultid="5277" />
                    <RANKING order="12" place="12" resultid="3766" />
                    <RANKING order="13" place="-1" resultid="2187" />
                    <RANKING order="14" place="-1" resultid="3098" />
                    <RANKING order="15" place="-1" resultid="3268" />
                    <RANKING order="16" place="-1" resultid="3638" />
                    <RANKING order="17" place="-1" resultid="3921" />
                    <RANKING order="18" place="-1" resultid="6062" />
                    <RANKING order="19" place="-1" resultid="3483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1662" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1924" />
                    <RANKING order="2" place="2" resultid="5295" />
                    <RANKING order="3" place="3" resultid="4664" />
                    <RANKING order="4" place="4" resultid="3229" />
                    <RANKING order="5" place="5" resultid="2692" />
                    <RANKING order="6" place="6" resultid="3835" />
                    <RANKING order="7" place="7" resultid="2159" />
                    <RANKING order="8" place="8" resultid="1889" />
                    <RANKING order="9" place="9" resultid="3326" />
                    <RANKING order="10" place="10" resultid="5014" />
                    <RANKING order="11" place="11" resultid="2165" />
                    <RANKING order="12" place="12" resultid="3772" />
                    <RANKING order="13" place="13" resultid="3262" />
                    <RANKING order="14" place="-1" resultid="5896" />
                    <RANKING order="15" place="-1" resultid="2712" />
                    <RANKING order="16" place="-1" resultid="4539" />
                    <RANKING order="17" place="-1" resultid="5323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1663" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3335" />
                    <RANKING order="2" place="2" resultid="2558" />
                    <RANKING order="3" place="3" resultid="3623" />
                    <RANKING order="4" place="4" resultid="2154" />
                    <RANKING order="5" place="5" resultid="5640" />
                    <RANKING order="6" place="6" resultid="4500" />
                    <RANKING order="7" place="7" resultid="4960" />
                    <RANKING order="8" place="8" resultid="5526" />
                    <RANKING order="9" place="9" resultid="3207" />
                    <RANKING order="10" place="10" resultid="6123" />
                    <RANKING order="11" place="-1" resultid="3628" />
                    <RANKING order="12" place="-1" resultid="4094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1664" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4426" />
                    <RANKING order="2" place="2" resultid="6185" />
                    <RANKING order="3" place="3" resultid="4692" />
                    <RANKING order="4" place="4" resultid="2049" />
                    <RANKING order="5" place="5" resultid="4481" />
                    <RANKING order="6" place="6" resultid="5644" />
                    <RANKING order="7" place="7" resultid="3193" />
                    <RANKING order="8" place="8" resultid="4588" />
                    <RANKING order="9" place="9" resultid="5660" />
                    <RANKING order="10" place="10" resultid="3461" />
                    <RANKING order="11" place="-1" resultid="2148" />
                    <RANKING order="12" place="-1" resultid="4614" />
                    <RANKING order="13" place="-1" resultid="3633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1665" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5001" />
                    <RANKING order="2" place="2" resultid="2687" />
                    <RANKING order="3" place="3" resultid="2725" />
                    <RANKING order="4" place="4" resultid="4510" />
                    <RANKING order="5" place="5" resultid="5512" />
                    <RANKING order="6" place="6" resultid="3307" />
                    <RANKING order="7" place="7" resultid="3155" />
                    <RANKING order="8" place="8" resultid="1897" />
                    <RANKING order="9" place="9" resultid="3971" />
                    <RANKING order="10" place="10" resultid="6447" />
                    <RANKING order="11" place="-1" resultid="2741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1666" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4317" />
                    <RANKING order="2" place="2" resultid="4279" />
                    <RANKING order="3" place="3" resultid="4575" />
                    <RANKING order="4" place="4" resultid="2749" />
                    <RANKING order="5" place="5" resultid="4441" />
                    <RANKING order="6" place="6" resultid="1999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1667" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4580" />
                    <RANKING order="2" place="2" resultid="4459" />
                    <RANKING order="3" place="3" resultid="5973" />
                    <RANKING order="4" place="-1" resultid="5621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1668" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2666" />
                    <RANKING order="2" place="2" resultid="2619" />
                    <RANKING order="3" place="3" resultid="2363" />
                    <RANKING order="4" place="4" resultid="4496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1670" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8029" daytime="11:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8030" daytime="11:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8031" daytime="11:13" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8032" daytime="11:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8033" daytime="11:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8034" daytime="11:17" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8035" daytime="11:19" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8036" daytime="11:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8037" daytime="11:22" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8038" daytime="11:23" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="8039" daytime="11:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="8040" daytime="11:26" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="8041" daytime="11:27" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="8042" daytime="11:29" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="8043" daytime="11:30" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="8044" daytime="11:31" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="8045" daytime="11:33" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="8046" daytime="11:34" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="8047" daytime="11:35" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="8048" daytime="11:37" number="20" order="20" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1671" daytime="11:38" gender="X" number="38" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1719" agemax="96" agemin="80" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="1720" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4113" />
                    <RANKING order="2" place="2" resultid="4809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1721" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5984" />
                    <RANKING order="2" place="2" resultid="5662" />
                    <RANKING order="3" place="3" resultid="4807" />
                    <RANKING order="4" place="4" resultid="6078" />
                    <RANKING order="5" place="5" resultid="3000" />
                    <RANKING order="6" place="6" resultid="3977" />
                    <RANKING order="7" place="7" resultid="3085" />
                    <RANKING order="8" place="8" resultid="3707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1722" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3974" />
                    <RANKING order="2" place="2" resultid="6456" />
                    <RANKING order="3" place="3" resultid="6080" />
                    <RANKING order="4" place="4" resultid="5491" />
                    <RANKING order="5" place="5" resultid="4712" />
                    <RANKING order="6" place="-1" resultid="4116" />
                    <RANKING order="7" place="-1" resultid="5796" />
                    <RANKING order="8" place="-1" resultid="3082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1723" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5056" />
                    <RANKING order="2" place="2" resultid="4388" />
                    <RANKING order="3" place="3" resultid="3979" />
                    <RANKING order="4" place="4" resultid="5057" />
                    <RANKING order="5" place="-1" resultid="2191" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1724" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4387" />
                    <RANKING order="2" place="-1" resultid="4630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1725" agemax="400" agemin="280" name="Kategoria F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4386" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8049" daytime="11:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8050" daytime="11:43" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8051" daytime="11:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8052" daytime="11:50" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1687" daytime="11:53" gender="F" number="39" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1688" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2575" />
                    <RANKING order="2" place="2" resultid="3913" />
                    <RANKING order="3" place="3" resultid="2610" />
                    <RANKING order="4" place="4" resultid="3958" />
                    <RANKING order="5" place="5" resultid="3783" />
                    <RANKING order="6" place="6" resultid="6258" />
                    <RANKING order="7" place="-1" resultid="5581" />
                    <RANKING order="8" place="-1" resultid="5843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1689" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6355" />
                    <RANKING order="2" place="2" resultid="4051" />
                    <RANKING order="3" place="3" resultid="4679" />
                    <RANKING order="4" place="4" resultid="3848" />
                    <RANKING order="5" place="5" resultid="4798" />
                    <RANKING order="6" place="6" resultid="5239" />
                    <RANKING order="7" place="7" resultid="3076" />
                    <RANKING order="8" place="8" resultid="4413" />
                    <RANKING order="9" place="9" resultid="3081" />
                    <RANKING order="10" place="10" resultid="5314" />
                    <RANKING order="11" place="11" resultid="3129" />
                    <RANKING order="12" place="-1" resultid="5364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1690" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2275" />
                    <RANKING order="2" place="2" resultid="4791" />
                    <RANKING order="3" place="3" resultid="5105" />
                    <RANKING order="4" place="4" resultid="5945" />
                    <RANKING order="5" place="5" resultid="4033" />
                    <RANKING order="6" place="6" resultid="6018" />
                    <RANKING order="7" place="7" resultid="6465" />
                    <RANKING order="8" place="8" resultid="3755" />
                    <RANKING order="9" place="-1" resultid="5785" />
                    <RANKING order="10" place="-1" resultid="5878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1691" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3698" />
                    <RANKING order="2" place="2" resultid="2231" />
                    <RANKING order="3" place="3" resultid="4025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1692" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4310" />
                    <RANKING order="2" place="2" resultid="5486" />
                    <RANKING order="3" place="3" resultid="3645" />
                    <RANKING order="4" place="4" resultid="6461" />
                    <RANKING order="5" place="5" resultid="6131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1693" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3108" />
                    <RANKING order="2" place="2" resultid="6076" />
                    <RANKING order="3" place="3" resultid="3222" />
                    <RANKING order="4" place="4" resultid="4418" />
                    <RANKING order="5" place="-1" resultid="2374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1694" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3043" />
                    <RANKING order="2" place="2" resultid="3940" />
                    <RANKING order="3" place="3" resultid="4686" />
                    <RANKING order="4" place="4" resultid="6368" />
                    <RANKING order="5" place="5" resultid="4566" />
                    <RANKING order="6" place="6" resultid="3138" />
                    <RANKING order="7" place="7" resultid="2766" />
                    <RANKING order="8" place="-1" resultid="4560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1695" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3931" />
                    <RANKING order="2" place="-1" resultid="2133" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1696" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5391" />
                    <RANKING order="2" place="-1" resultid="6318" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1697" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1698" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1699" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="1700" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1701" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1702" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9047" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9048" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9049" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9050" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9051" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9052" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9053" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1703" daytime="12:59" gender="M" number="40" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1704" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5162" />
                    <RANKING order="2" place="2" resultid="3662" />
                    <RANKING order="3" place="3" resultid="2211" />
                    <RANKING order="4" place="4" resultid="4761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1705" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5959" />
                    <RANKING order="2" place="2" resultid="2026" />
                    <RANKING order="3" place="3" resultid="2054" />
                    <RANKING order="4" place="4" resultid="3840" />
                    <RANKING order="5" place="5" resultid="5405" />
                    <RANKING order="6" place="6" resultid="3900" />
                    <RANKING order="7" place="7" resultid="5385" />
                    <RANKING order="8" place="8" resultid="5435" />
                    <RANKING order="9" place="9" resultid="5119" />
                    <RANKING order="10" place="-1" resultid="4779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1706" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5606" />
                    <RANKING order="2" place="2" resultid="3243" />
                    <RANKING order="3" place="3" resultid="2072" />
                    <RANKING order="4" place="4" resultid="3065" />
                    <RANKING order="5" place="5" resultid="4805" />
                    <RANKING order="6" place="6" resultid="4160" />
                    <RANKING order="7" place="7" resultid="3585" />
                    <RANKING order="8" place="8" resultid="2394" />
                    <RANKING order="9" place="9" resultid="5247" />
                    <RANKING order="10" place="10" resultid="5593" />
                    <RANKING order="11" place="11" resultid="5300" />
                    <RANKING order="12" place="12" resultid="3524" />
                    <RANKING order="13" place="-1" resultid="1995" />
                    <RANKING order="14" place="-1" resultid="3744" />
                    <RANKING order="15" place="-1" resultid="5635" />
                    <RANKING order="16" place="-1" resultid="5968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1707" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2314" />
                    <RANKING order="2" place="2" resultid="5559" />
                    <RANKING order="3" place="3" resultid="6055" />
                    <RANKING order="4" place="4" resultid="3114" />
                    <RANKING order="5" place="5" resultid="3762" />
                    <RANKING order="6" place="6" resultid="2401" />
                    <RANKING order="7" place="7" resultid="4211" />
                    <RANKING order="8" place="8" resultid="5147" />
                    <RANKING order="9" place="9" resultid="3057" />
                    <RANKING order="10" place="10" resultid="2977" />
                    <RANKING order="11" place="11" resultid="1952" />
                    <RANKING order="12" place="12" resultid="5983" />
                    <RANKING order="13" place="13" resultid="5440" />
                    <RANKING order="14" place="-1" resultid="4710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1708" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6180" />
                    <RANKING order="2" place="2" resultid="2780" />
                    <RANKING order="3" place="3" resultid="5193" />
                    <RANKING order="4" place="4" resultid="6375" />
                    <RANKING order="5" place="5" resultid="6189" />
                    <RANKING order="6" place="6" resultid="5222" />
                    <RANKING order="7" place="7" resultid="4434" />
                    <RANKING order="8" place="8" resultid="6379" />
                    <RANKING order="9" place="9" resultid="5096" />
                    <RANKING order="10" place="10" resultid="2981" />
                    <RANKING order="11" place="11" resultid="4751" />
                    <RANKING order="12" place="-1" resultid="2599" />
                    <RANKING order="13" place="-1" resultid="5421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1709" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3657" />
                    <RANKING order="2" place="2" resultid="6197" />
                    <RANKING order="3" place="3" resultid="2182" />
                    <RANKING order="4" place="4" resultid="5890" />
                    <RANKING order="5" place="5" resultid="2042" />
                    <RANKING order="6" place="6" resultid="2696" />
                    <RANKING order="7" place="7" resultid="3020" />
                    <RANKING order="8" place="8" resultid="6063" />
                    <RANKING order="9" place="9" resultid="3727" />
                    <RANKING order="10" place="10" resultid="3922" />
                    <RANKING order="11" place="-1" resultid="3484" />
                    <RANKING order="12" place="-1" resultid="5712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1710" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3257" />
                    <RANKING order="2" place="2" resultid="3652" />
                    <RANKING order="3" place="3" resultid="6041" />
                    <RANKING order="4" place="4" resultid="3773" />
                    <RANKING order="5" place="5" resultid="4728" />
                    <RANKING order="6" place="6" resultid="5270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1711" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6011" />
                    <RANKING order="2" place="2" resultid="3611" />
                    <RANKING order="3" place="3" resultid="2642" />
                    <RANKING order="4" place="4" resultid="6289" />
                    <RANKING order="5" place="5" resultid="5429" />
                    <RANKING order="6" place="6" resultid="5199" />
                    <RANKING order="7" place="-1" resultid="1868" />
                    <RANKING order="8" place="-1" resultid="2756" />
                    <RANKING order="9" place="-1" resultid="6124" />
                    <RANKING order="10" place="-1" resultid="3052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1712" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4615" />
                    <RANKING order="2" place="2" resultid="2815" />
                    <RANKING order="3" place="3" resultid="3453" />
                    <RANKING order="4" place="4" resultid="2657" />
                    <RANKING order="5" place="5" resultid="2674" />
                    <RANKING order="6" place="6" resultid="3462" />
                    <RANKING order="7" place="-1" resultid="4544" />
                    <RANKING order="8" place="-1" resultid="5518" />
                    <RANKING order="9" place="-1" resultid="4983" />
                    <RANKING order="10" place="-1" resultid="5613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1713" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2244" />
                    <RANKING order="2" place="2" resultid="3818" />
                    <RANKING order="3" place="3" resultid="2408" />
                    <RANKING order="4" place="4" resultid="3297" />
                    <RANKING order="5" place="-1" resultid="3443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1714" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4298" />
                    <RANKING order="2" place="2" resultid="3797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1715" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1716" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2620" />
                    <RANKING order="2" place="2" resultid="2018" />
                    <RANKING order="3" place="3" resultid="5167" />
                    <RANKING order="4" place="-1" resultid="1961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1717" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1718" agemax="94" agemin="90" name="Kategoria  N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9059" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9060" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9061" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9062" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9063" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9064" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9065" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9066" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9067" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9068" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9069" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="9070" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="8925" />
            <JUDGE officialid="8910" />
            <JUDGE officialid="8924" />
            <JUDGE officialid="8926" />
            <JUDGE officialid="8906" />
            <JUDGE officialid="8919" />
            <JUDGE officialid="8923" />
            <JUDGE officialid="8909" />
            <JUDGE officialid="8921" />
            <JUDGE officialid="8914" />
            <JUDGE officialid="8915" />
            <JUDGE officialid="8918" />
            <JUDGE officialid="8922" />
            <JUDGE officialid="8917" />
            <JUDGE officialid="8920" />
            <JUDGE officialid="8928" />
            <JUDGE officialid="8912" />
            <JUDGE officialid="8916" />
            <JUDGE officialid="8916" />
            <JUDGE officialid="8908" />
            <JUDGE officialid="8908" />
            <JUDGE officialid="8911" />
            <JUDGE officialid="8911" />
            <JUDGE officialid="8913" />
            <JUDGE officialid="8927" />
            <JUDGE officialid="8905" />
            <JUDGE officialid="8904" />
            <JUDGE officialid="8903" />
            <JUDGE officialid="8907" />
            <JUDGE officialid="8941" />
            <JUDGE officialid="8901" />
            <JUDGE officialid="8902" />
          </JUDGES>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="00611" nation="POL" region="11" clubid="5153" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1991-09-13" firstname="Tomasz" gender="M" lastname="Czermak" nation="POL" license="100611200197" athleteid="5154">
              <RESULTS>
                <RESULT eventid="1108" points="800" reactiontime="+74" swimtime="00:02:16.77" resultid="5155" heatid="7733" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="100" swimtime="00:01:06.36" />
                    <SPLIT distance="150" swimtime="00:01:44.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="726" reactiontime="+76" swimtime="00:17:46.83" resultid="5156" heatid="8717" lane="6" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="150" swimtime="00:01:40.35" />
                    <SPLIT distance="200" swimtime="00:02:15.48" />
                    <SPLIT distance="250" swimtime="00:02:50.61" />
                    <SPLIT distance="300" swimtime="00:03:26.35" />
                    <SPLIT distance="350" swimtime="00:04:02.10" />
                    <SPLIT distance="400" swimtime="00:04:37.57" />
                    <SPLIT distance="450" swimtime="00:05:13.43" />
                    <SPLIT distance="500" swimtime="00:05:49.27" />
                    <SPLIT distance="550" swimtime="00:06:25.22" />
                    <SPLIT distance="600" swimtime="00:07:01.07" />
                    <SPLIT distance="650" swimtime="00:07:37.41" />
                    <SPLIT distance="700" swimtime="00:08:13.54" />
                    <SPLIT distance="750" swimtime="00:08:49.50" />
                    <SPLIT distance="800" swimtime="00:09:25.14" />
                    <SPLIT distance="850" swimtime="00:10:00.93" />
                    <SPLIT distance="900" swimtime="00:10:36.74" />
                    <SPLIT distance="950" swimtime="00:11:12.96" />
                    <SPLIT distance="1000" swimtime="00:11:49.29" />
                    <SPLIT distance="1050" swimtime="00:12:25.34" />
                    <SPLIT distance="1100" swimtime="00:13:01.50" />
                    <SPLIT distance="1150" swimtime="00:13:37.28" />
                    <SPLIT distance="1200" swimtime="00:14:13.35" />
                    <SPLIT distance="1250" swimtime="00:14:49.66" />
                    <SPLIT distance="1300" swimtime="00:15:26.05" />
                    <SPLIT distance="1350" swimtime="00:16:02.25" />
                    <SPLIT distance="1400" swimtime="00:16:37.85" />
                    <SPLIT distance="1450" swimtime="00:17:13.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="786" reactiontime="+73" swimtime="00:02:31.15" resultid="5157" heatid="7795" lane="4" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                    <SPLIT distance="150" swimtime="00:01:52.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="607" reactiontime="+75" swimtime="00:02:27.40" resultid="5158" heatid="7865" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                    <SPLIT distance="150" swimtime="00:01:48.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="744" reactiontime="+74" swimtime="00:01:08.16" resultid="5159" heatid="7896" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="696" reactiontime="+72" swimtime="00:05:02.77" resultid="5160" heatid="8806" lane="4" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:10.78" />
                    <SPLIT distance="150" swimtime="00:01:50.94" />
                    <SPLIT distance="200" swimtime="00:02:30.75" />
                    <SPLIT distance="250" swimtime="00:03:11.49" />
                    <SPLIT distance="300" swimtime="00:03:53.59" />
                    <SPLIT distance="350" swimtime="00:04:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="771" reactiontime="+70" swimtime="00:00:30.81" resultid="5161" heatid="8048" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1703" points="772" reactiontime="+71" swimtime="00:04:27.49" resultid="5162" heatid="9059" lane="4" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="100" swimtime="00:01:02.98" />
                    <SPLIT distance="150" swimtime="00:01:36.64" />
                    <SPLIT distance="200" swimtime="00:02:10.77" />
                    <SPLIT distance="250" swimtime="00:02:45.12" />
                    <SPLIT distance="300" swimtime="00:03:20.25" />
                    <SPLIT distance="350" swimtime="00:03:55.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1931-04-27" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" athleteid="5163">
              <RESULTS>
                <RESULT eventid="1156" points="296" swimtime="00:44:50.33" resultid="5164" heatid="8725" lane="5" entrytime="00:45:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.47" />
                    <SPLIT distance="100" swimtime="00:02:44.04" />
                    <SPLIT distance="200" swimtime="00:05:43.87" />
                    <SPLIT distance="300" swimtime="00:08:43.74" />
                    <SPLIT distance="400" swimtime="00:11:42.22" />
                    <SPLIT distance="500" swimtime="00:14:44.26" />
                    <SPLIT distance="600" swimtime="00:17:47.70" />
                    <SPLIT distance="700" swimtime="00:20:52.97" />
                    <SPLIT distance="800" swimtime="00:23:54.77" />
                    <SPLIT distance="900" swimtime="00:26:57.93" />
                    <SPLIT distance="1000" swimtime="00:30:00.11" />
                    <SPLIT distance="1100" swimtime="00:33:00.42" />
                    <SPLIT distance="1200" swimtime="00:35:59.83" />
                    <SPLIT distance="1300" swimtime="00:39:00.11" />
                    <SPLIT distance="1400" swimtime="00:41:57.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="318" reactiontime="+106" swimtime="00:05:23.08" resultid="5165" heatid="7785" lane="7" entrytime="00:05:22.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.84" />
                    <SPLIT distance="100" swimtime="00:02:33.78" />
                    <SPLIT distance="150" swimtime="00:04:00.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="209" reactiontime="+123" swimtime="00:05:03.23" resultid="5166" heatid="7952" lane="3" entrytime="00:05:09.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.32" />
                    <SPLIT distance="100" swimtime="00:02:24.40" />
                    <SPLIT distance="150" swimtime="00:03:46.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="219" reactiontime="+93" swimtime="00:10:46.77" resultid="5167" heatid="9070" lane="6" entrytime="00:10:50.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.73" />
                    <SPLIT distance="100" swimtime="00:02:33.96" />
                    <SPLIT distance="150" swimtime="00:03:58.09" />
                    <SPLIT distance="200" swimtime="00:05:20.75" />
                    <SPLIT distance="250" swimtime="00:06:43.52" />
                    <SPLIT distance="300" swimtime="00:08:06.56" />
                    <SPLIT distance="350" swimtime="00:09:30.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZRAC" nation="POL" region="11" clubid="2550" name="AZS PWSZ Racibórz">
          <CONTACT city="Racibórz" email="m,kunicki@" name="Kunicki" phone="504 233 267" state="ŚLĄSK" street="Słowackiego55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-04-11" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="2551">
              <RESULTS>
                <RESULT eventid="1108" points="593" reactiontime="+92" swimtime="00:02:56.36" resultid="2552" heatid="7726" lane="5" entrytime="00:02:56.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:23.00" />
                    <SPLIT distance="150" swimtime="00:02:15.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="525" reactiontime="+97" swimtime="00:03:21.48" resultid="2553" heatid="7791" lane="2" entrytime="00:03:13.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                    <SPLIT distance="100" swimtime="00:01:35.37" />
                    <SPLIT distance="150" swimtime="00:02:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="485" reactiontime="+100" swimtime="00:03:07.85" resultid="2554" heatid="7863" lane="1" entrytime="00:03:05.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                    <SPLIT distance="150" swimtime="00:02:19.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="495" reactiontime="+91" swimtime="00:01:26.11" resultid="2555" heatid="7890" lane="6" entrytime="00:01:24.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="603" reactiontime="+114" swimtime="00:06:23.61" resultid="2556" heatid="8809" lane="6" entrytime="00:06:25.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                    <SPLIT distance="100" swimtime="00:01:35.97" />
                    <SPLIT distance="150" swimtime="00:02:25.49" />
                    <SPLIT distance="200" swimtime="00:03:13.65" />
                    <SPLIT distance="250" swimtime="00:04:08.06" />
                    <SPLIT distance="300" swimtime="00:05:01.18" />
                    <SPLIT distance="350" swimtime="00:05:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="455" reactiontime="+92" swimtime="00:01:24.18" resultid="2557" heatid="7996" lane="4" entrytime="00:01:21.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="519" reactiontime="+85" swimtime="00:00:37.94" resultid="2558" heatid="8040" lane="7" entrytime="00:00:37.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01113" nation="POL" region="13" clubid="5989" name="AZS UWM Masters Olsztyn">
          <CONTACT city="Łupstych" email="gozdzik@uwm.edu.pl" name="Goździejewska Anna" state="WARM-" street="Leśna 1" zip="11-041" />
          <ATHLETES>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="6004">
              <RESULTS>
                <RESULT eventid="1108" points="892" reactiontime="+84" swimtime="00:02:33.92" resultid="6005" heatid="7730" lane="5" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:11.46" />
                    <SPLIT distance="150" swimtime="00:01:57.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="956" reactiontime="+84" swimtime="00:01:10.22" resultid="6006" heatid="7840" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="6007" heatid="7865" lane="8" entrytime="00:02:42.00" />
                <RESULT eventid="1415" points="821" reactiontime="+85" swimtime="00:00:30.45" resultid="6008" heatid="7908" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1447" points="803" reactiontime="+85" swimtime="00:01:13.84" resultid="6009" heatid="7940" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="826" reactiontime="+82" swimtime="00:01:09.02" resultid="6010" heatid="8001" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="869" reactiontime="+94" swimtime="00:05:02.78" resultid="6011" heatid="9063" lane="7" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:12.12" />
                    <SPLIT distance="150" swimtime="00:01:50.45" />
                    <SPLIT distance="200" swimtime="00:02:29.20" />
                    <SPLIT distance="250" swimtime="00:03:08.10" />
                    <SPLIT distance="300" swimtime="00:03:46.89" />
                    <SPLIT distance="350" swimtime="00:04:25.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-26" firstname="Aleksandra" gender="F" lastname="Przybysz" nation="POL" athleteid="6012">
              <RESULTS>
                <RESULT eventid="1140" points="453" swimtime="00:12:32.78" resultid="6013" heatid="8713" lane="7" entrytime="00:12:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:01:26.09" />
                    <SPLIT distance="200" swimtime="00:02:58.79" />
                    <SPLIT distance="300" swimtime="00:04:33.34" />
                    <SPLIT distance="400" swimtime="00:06:08.03" />
                    <SPLIT distance="500" swimtime="00:07:42.53" />
                    <SPLIT distance="600" swimtime="00:09:18.29" />
                    <SPLIT distance="700" swimtime="00:10:55.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="433" reactiontime="+96" swimtime="00:01:15.96" resultid="6014" heatid="7801" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="380" reactiontime="+95" swimtime="00:00:40.09" resultid="6015" heatid="7900" lane="8" entrytime="00:00:41.00" />
                <RESULT eventid="1463" points="400" reactiontime="+90" swimtime="00:02:50.90" resultid="6016" heatid="7948" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:22.13" />
                    <SPLIT distance="150" swimtime="00:02:06.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="321" reactiontime="+91" swimtime="00:01:33.09" resultid="6017" heatid="7989" lane="7" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="417" reactiontime="+93" swimtime="00:06:06.02" resultid="6018" heatid="9050" lane="3" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:24.00" />
                    <SPLIT distance="150" swimtime="00:02:10.39" />
                    <SPLIT distance="200" swimtime="00:02:57.07" />
                    <SPLIT distance="250" swimtime="00:03:44.94" />
                    <SPLIT distance="300" swimtime="00:04:32.95" />
                    <SPLIT distance="350" swimtime="00:05:20.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="Piekut" nation="POL" athleteid="6019">
              <RESULTS>
                <RESULT eventid="1092" points="557" reactiontime="+84" swimtime="00:02:53.98" resultid="6020" heatid="7717" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:17.83" />
                    <SPLIT distance="150" swimtime="00:02:10.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="605" reactiontime="+74" swimtime="00:00:36.49" resultid="6021" heatid="7760" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1302" points="578" reactiontime="+90" swimtime="00:02:49.05" resultid="6022" heatid="7858" lane="4" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:20.66" />
                    <SPLIT distance="150" swimtime="00:02:05.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="637" reactiontime="+86" swimtime="00:00:33.78" resultid="6023" heatid="7903" lane="4" entrytime="00:00:34.25" />
                <RESULT eventid="1463" points="530" reactiontime="+88" swimtime="00:02:35.70" resultid="6024" heatid="7950" lane="1" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:14.78" />
                    <SPLIT distance="150" swimtime="00:01:56.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="618" reactiontime="+84" swimtime="00:01:15.09" resultid="6025" heatid="7991" lane="1" entrytime="00:01:16.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-01" firstname="Grzegorz" gender="M" lastname="Mówiński" nation="POL" athleteid="6026">
              <RESULTS>
                <RESULT eventid="1076" points="388" reactiontime="+87" swimtime="00:00:32.55" resultid="6027" heatid="7691" lane="7" entrytime="00:00:33.14" />
                <RESULT eventid="1286" points="320" reactiontime="+99" swimtime="00:01:27.37" resultid="6028" heatid="7842" lane="4" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="323" reactiontime="+81" swimtime="00:00:36.60" resultid="6029" heatid="7911" lane="1" entrytime="00:00:37.52" />
                <RESULT eventid="1591" points="265" reactiontime="+91" swimtime="00:01:28.08" resultid="6030" heatid="7995" lane="8" entrytime="00:01:37.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="6031">
              <RESULTS>
                <RESULT eventid="1173" points="531" reactiontime="+76" swimtime="00:00:37.47" resultid="6032" heatid="7759" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1270" points="530" reactiontime="+93" swimtime="00:01:20.44" resultid="6033" heatid="7834" lane="3" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="572" reactiontime="+95" swimtime="00:00:34.99" resultid="6034" heatid="7903" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1431" points="538" reactiontime="+77" swimtime="00:01:21.81" resultid="6035" heatid="7930" lane="1" entrytime="00:01:23.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="524" reactiontime="+79" swimtime="00:02:55.60" resultid="6036" heatid="8007" lane="5" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:26.86" />
                    <SPLIT distance="150" swimtime="00:02:12.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-09" firstname="Marek" gender="M" lastname="Koźlikowski" nation="POL" athleteid="6037">
              <RESULTS>
                <RESULT eventid="1254" points="507" reactiontime="+100" swimtime="00:01:10.74" resultid="6038" heatid="7807" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="482" reactiontime="+101" swimtime="00:01:23.52" resultid="6039" heatid="7845" lane="4" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="439" reactiontime="+106" swimtime="00:02:45.44" resultid="6040" heatid="7959" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:02:02.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="403" reactiontime="+104" swimtime="00:06:00.43" resultid="6041" heatid="9065" lane="6" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:11.36" />
                    <SPLIT distance="200" swimtime="00:02:57.73" />
                    <SPLIT distance="250" swimtime="00:03:45.11" />
                    <SPLIT distance="300" swimtime="00:04:31.52" />
                    <SPLIT distance="350" swimtime="00:05:18.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-13" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="6042">
              <RESULTS>
                <RESULT eventid="1222" points="656" reactiontime="+72" swimtime="00:02:41.68" resultid="6043" heatid="7794" lane="4" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="150" swimtime="00:01:57.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="584" reactiontime="+70" swimtime="00:01:13.35" resultid="6044" heatid="7894" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="501" reactiontime="+73" swimtime="00:05:36.12" resultid="6045" heatid="8806" lane="2" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:01.93" />
                    <SPLIT distance="200" swimtime="00:02:43.41" />
                    <SPLIT distance="250" swimtime="00:03:28.87" />
                    <SPLIT distance="300" swimtime="00:04:14.84" />
                    <SPLIT distance="350" swimtime="00:04:56.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="594" reactiontime="+68" swimtime="00:00:33.08" resultid="6046" heatid="8045" lane="3" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="6047">
              <RESULTS>
                <RESULT eventid="1076" points="762" reactiontime="+76" swimtime="00:00:25.96" resultid="6048" heatid="7708" lane="3" entrytime="00:00:26.64" />
                <RESULT eventid="1108" points="626" reactiontime="+82" swimtime="00:02:28.78" resultid="6049" heatid="7730" lane="7" entrytime="00:02:36.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:11.49" />
                    <SPLIT distance="150" swimtime="00:01:53.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="774" reactiontime="+80" swimtime="00:00:56.01" resultid="6050" heatid="7807" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="695" reactiontime="+78" swimtime="00:01:06.65" resultid="6051" heatid="7852" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="727" reactiontime="+80" swimtime="00:00:28.53" resultid="6052" heatid="7922" lane="7" entrytime="00:00:28.60" />
                <RESULT eventid="1479" points="671" reactiontime="+82" swimtime="00:02:07.27" resultid="6053" heatid="7965" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                    <SPLIT distance="100" swimtime="00:01:00.41" />
                    <SPLIT distance="150" swimtime="00:01:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="676" reactiontime="+83" swimtime="00:01:04.77" resultid="6054" heatid="8000" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="644" reactiontime="+95" swimtime="00:04:40.60" resultid="6055" heatid="9059" lane="8" entrytime="00:04:44.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:06.66" />
                    <SPLIT distance="150" swimtime="00:01:41.56" />
                    <SPLIT distance="200" swimtime="00:02:17.25" />
                    <SPLIT distance="250" swimtime="00:02:52.82" />
                    <SPLIT distance="300" swimtime="00:03:28.96" />
                    <SPLIT distance="350" swimtime="00:04:05.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-25" firstname="Piotr" gender="M" lastname="Markowicz" nation="POL" athleteid="6056">
              <RESULTS>
                <RESULT eventid="1108" points="579" reactiontime="+88" swimtime="00:02:43.88" resultid="6057" heatid="7728" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                    <SPLIT distance="150" swimtime="00:02:02.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="430" swimtime="00:21:49.79" resultid="6058" heatid="8721" lane="5" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:20.19" />
                    <SPLIT distance="200" swimtime="00:02:44.37" />
                    <SPLIT distance="300" swimtime="00:04:10.61" />
                    <SPLIT distance="400" swimtime="00:05:37.19" />
                    <SPLIT distance="500" swimtime="00:07:04.62" />
                    <SPLIT distance="600" swimtime="00:08:31.53" />
                    <SPLIT distance="700" swimtime="00:09:57.87" />
                    <SPLIT distance="800" swimtime="00:11:26.11" />
                    <SPLIT distance="900" swimtime="00:12:52.78" />
                    <SPLIT distance="1000" swimtime="00:14:20.61" />
                    <SPLIT distance="1100" swimtime="00:15:48.59" />
                    <SPLIT distance="1200" swimtime="00:17:18.36" />
                    <SPLIT distance="1300" swimtime="00:18:48.77" />
                    <SPLIT distance="1400" swimtime="00:20:20.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="522" reactiontime="+90" swimtime="00:01:15.11" resultid="6059" heatid="7849" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="556" reactiontime="+77" swimtime="00:01:15.56" resultid="6060" heatid="7938" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="6061" heatid="7960" lane="1" entrytime="00:02:35.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="6062" heatid="8039" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1703" points="441" reactiontime="+97" swimtime="00:05:22.93" resultid="6063" heatid="9062" lane="8" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:57.15" />
                    <SPLIT distance="200" swimtime="00:02:37.94" />
                    <SPLIT distance="250" swimtime="00:03:18.29" />
                    <SPLIT distance="300" swimtime="00:03:58.78" />
                    <SPLIT distance="350" swimtime="00:04:40.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-02" firstname="Piotr" gender="M" lastname="Suchecki" nation="POL" athleteid="6064">
              <RESULTS>
                <RESULT eventid="1190" points="677" reactiontime="+79" swimtime="00:00:30.90" resultid="6065" heatid="7777" lane="8" entrytime="00:00:29.92" />
                <RESULT eventid="1286" points="633" reactiontime="+79" swimtime="00:01:08.76" resultid="6066" heatid="7853" lane="4" entrytime="00:01:07.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="698" reactiontime="+83" swimtime="00:00:28.92" resultid="6067" heatid="7924" lane="1" entrytime="00:00:27.42" />
                <RESULT eventid="1591" points="550" reactiontime="+85" swimtime="00:01:09.37" resultid="6068" heatid="8002" lane="1" entrytime="00:01:03.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="6069">
              <RESULTS>
                <RESULT eventid="1140" points="519" swimtime="00:11:56.35" resultid="6070" heatid="8713" lane="4" entrytime="00:12:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:25.96" />
                    <SPLIT distance="200" swimtime="00:02:56.59" />
                    <SPLIT distance="300" swimtime="00:04:28.12" />
                    <SPLIT distance="400" swimtime="00:05:58.54" />
                    <SPLIT distance="500" swimtime="00:07:28.18" />
                    <SPLIT distance="600" swimtime="00:08:58.79" />
                    <SPLIT distance="700" swimtime="00:10:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="581" reactiontime="+89" swimtime="00:03:24.13" resultid="6071" heatid="7781" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                    <SPLIT distance="100" swimtime="00:01:39.16" />
                    <SPLIT distance="150" swimtime="00:02:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="534" reactiontime="+86" swimtime="00:01:26.95" resultid="6072" heatid="7832" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="538" reactiontime="+86" swimtime="00:02:44.38" resultid="6073" heatid="7945" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="150" swimtime="00:02:00.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="562" reactiontime="+93" swimtime="00:06:36.88" resultid="6074" heatid="8802" lane="1" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                    <SPLIT distance="100" swimtime="00:01:40.05" />
                    <SPLIT distance="150" swimtime="00:02:30.37" />
                    <SPLIT distance="200" swimtime="00:03:18.82" />
                    <SPLIT distance="250" swimtime="00:04:12.13" />
                    <SPLIT distance="300" swimtime="00:05:06.67" />
                    <SPLIT distance="350" swimtime="00:05:52.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="469" reactiontime="+80" swimtime="00:03:17.79" resultid="6075" heatid="8005" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:36.68" />
                    <SPLIT distance="150" swimtime="00:02:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="557" reactiontime="+87" swimtime="00:05:44.85" resultid="6076" heatid="9049" lane="4" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                    <SPLIT distance="150" swimtime="00:02:04.54" />
                    <SPLIT distance="200" swimtime="00:02:49.29" />
                    <SPLIT distance="250" swimtime="00:03:34.34" />
                    <SPLIT distance="300" swimtime="00:04:19.14" />
                    <SPLIT distance="350" swimtime="00:05:03.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="AZS UWM Masters Olsztyn C" number="1">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+80" swimtime="00:02:00.93" resultid="6081" heatid="7871" lane="5" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:04.52" />
                    <SPLIT distance="150" swimtime="00:01:33.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6064" number="1" />
                    <RELAYPOSITION athleteid="6042" number="2" />
                    <RELAYPOSITION athleteid="6026" number="3" />
                    <RELAYPOSITION athleteid="6004" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" reactiontime="+92" swimtime="00:02:00.83" resultid="6082" heatid="7972" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:01:00.64" />
                    <SPLIT distance="150" swimtime="00:01:32.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6056" number="1" />
                    <RELAYPOSITION athleteid="6037" number="2" />
                    <RELAYPOSITION athleteid="6026" number="3" />
                    <RELAYPOSITION athleteid="6064" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="AZS UWM Masters Olsztyn B" number="1">
              <RESULTS>
                <RESULT eventid="1495" reactiontime="+87" swimtime="00:02:12.04" resultid="6077" heatid="7969" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:05.48" />
                    <SPLIT distance="150" swimtime="00:01:38.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6031" number="1" />
                    <RELAYPOSITION athleteid="6069" number="2" />
                    <RELAYPOSITION athleteid="6019" number="3" />
                    <RELAYPOSITION athleteid="6012" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" reactiontime="+77" swimtime="00:02:28.60" resultid="6079" heatid="7866" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="100" swimtime="00:01:22.03" />
                    <SPLIT distance="150" swimtime="00:01:55.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6031" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="6069" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="6019" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="6012" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="AZS UWM Masters Olsztyn B" number="1">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+82" swimtime="00:02:09.61" resultid="6078" heatid="8051" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:04.34" />
                    <SPLIT distance="150" swimtime="00:01:38.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6064" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="6042" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="6019" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="6031" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="AZS UWM Masters Olsztyn C" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+85" swimtime="00:02:09.55" resultid="6083" heatid="7736" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="150" swimtime="00:01:40.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6069" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="6019" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="6026" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="6004" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="AZS UWM Masters Olsztyn C" number="2">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+82" swimtime="00:02:22.22" resultid="6080" heatid="8051" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:19.33" />
                    <SPLIT distance="150" swimtime="00:01:48.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6056" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="6069" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="6047" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="6012" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AZDAB" nation="POL" region="11" clubid="6290" name="AZS WSB Dabrowa Grn.">
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="6209">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="6210" heatid="7710" lane="5" entrytime="00:00:26.00" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="6211" heatid="7732" lane="3" entrytime="00:02:24.00" />
                <RESULT eventid="1254" points="636" reactiontime="+70" swimtime="00:00:59.21" resultid="6212" heatid="7824" lane="5" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="6213" heatid="7851" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1415" points="653" reactiontime="+71" swimtime="00:00:28.80" resultid="6214" heatid="7924" lane="8" entrytime="00:00:27.50" />
                <RESULT eventid="1479" points="526" reactiontime="+68" swimtime="00:02:16.28" resultid="6215" heatid="7966" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="100" swimtime="00:01:02.49" />
                    <SPLIT distance="150" swimtime="00:01:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="6216" heatid="8047" lane="7" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZSUM" nation="POL" region="11" clubid="5668" name="AZS Śląski Uniwersytet Medyczny" shortname="AZS Śląski UM">
          <CONTACT name="Pałka Karol" />
          <ATHLETES>
            <ATHLETE birthdate="1990-03-18" firstname="Karol" gender="M" lastname="Pałka" nation="POL" athleteid="5686">
              <RESULTS>
                <RESULT eventid="1190" points="332" reactiontime="+69" swimtime="00:00:37.40" resultid="5687" heatid="7773" lane="5" entrytime="00:00:33.87" />
                <RESULT eventid="1222" points="430" reactiontime="+77" swimtime="00:03:04.83" resultid="5688" heatid="7794" lane="6" entrytime="00:02:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:26.10" />
                    <SPLIT distance="150" swimtime="00:02:14.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="5689" heatid="7847" lane="6" entrytime="00:01:16.00" entrycourse="SCM" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="5690" heatid="7893" lane="2" entrytime="00:01:19.00" entrycourse="SCM" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="5691" heatid="8044" lane="6" entrytime="00:00:34.67" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ARWAR" nation="POL" region="14" clubid="3668" name="Akademia Ruchu AG Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1977-02-11" firstname="Marcin" gender="M" lastname="Siwonia" nation="POL" athleteid="3669">
              <RESULTS>
                <RESULT eventid="1254" points="202" reactiontime="+89" swimtime="00:01:27.51" resultid="3670" heatid="7807" lane="3" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="130" reactiontime="+99" swimtime="00:02:06.27" resultid="3671" heatid="7882" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="173" reactiontime="+108" swimtime="00:03:19.90" resultid="3672" heatid="7954" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                    <SPLIT distance="100" swimtime="00:01:36.74" />
                    <SPLIT distance="150" swimtime="00:02:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="3673" heatid="7993" lane="8" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-22" firstname="Andrzej" gender="M" lastname="Gadaś" nation="POL" athleteid="3674">
              <RESULTS>
                <RESULT eventid="1076" points="457" reactiontime="+86" swimtime="00:00:28.72" resultid="3675" heatid="7701" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1254" points="409" reactiontime="+82" swimtime="00:01:06.04" resultid="3676" heatid="7814" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="389" reactiontime="+82" swimtime="00:01:15.33" resultid="3677" heatid="7846" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="429" reactiontime="+76" swimtime="00:01:21.27" resultid="3678" heatid="7893" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="450" reactiontime="+80" swimtime="00:00:36.29" resultid="3679" heatid="8041" lane="7" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-13" firstname="Izabela" gender="F" lastname="Chmielewska" nation="POL" athleteid="3680">
              <RESULTS>
                <RESULT eventid="1059" points="227" reactiontime="+86" swimtime="00:00:42.79" resultid="3681" heatid="7674" lane="3" entrytime="00:00:41.90" />
                <RESULT eventid="1173" status="DNS" swimtime="00:00:00.00" resultid="3682" heatid="7755" lane="2" entrytime="00:00:52.00" />
                <RESULT eventid="1238" points="198" reactiontime="+98" swimtime="00:01:38.45" resultid="3683" heatid="7798" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="195" reactiontime="+83" swimtime="00:00:50.04" resultid="3684" heatid="7898" lane="2" entrytime="00:00:52.00" />
                <RESULT eventid="1463" points="175" reactiontime="+90" swimtime="00:03:45.01" resultid="3685" heatid="7946" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                    <SPLIT distance="100" swimtime="00:01:42.85" />
                    <SPLIT distance="150" swimtime="00:02:43.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-07" firstname="Rafał" gender="M" lastname="Kowalczyk" nation="POL" athleteid="3686">
              <RESULTS>
                <RESULT eventid="1076" points="376" reactiontime="+76" swimtime="00:00:31.63" resultid="3687" heatid="7692" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="1190" points="196" reactiontime="+81" swimtime="00:00:43.08" resultid="3688" heatid="7766" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="1254" points="304" reactiontime="+89" swimtime="00:01:12.24" resultid="3689" heatid="7809" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M9 - Naprzemienna lub nierównoczesna praca nóg" eventid="1415" reactiontime="+92" status="DSQ" swimtime="00:00:38.17" resultid="3690" heatid="7909" lane="8" entrytime="00:00:41.50" />
                <RESULT eventid="1479" points="273" reactiontime="+91" swimtime="00:02:53.35" resultid="3691" heatid="7955" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:21.90" />
                    <SPLIT distance="150" swimtime="00:02:07.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-29" firstname="Marta" gender="F" lastname="Maryl" nation="POL" athleteid="3692">
              <RESULTS>
                <RESULT eventid="1140" points="485" swimtime="00:12:00.37" resultid="3693" heatid="8714" lane="8" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:01:24.22" />
                    <SPLIT distance="200" swimtime="00:02:55.55" />
                    <SPLIT distance="300" swimtime="00:04:27.93" />
                    <SPLIT distance="400" swimtime="00:05:54.71" />
                    <SPLIT distance="500" swimtime="00:07:31.67" />
                    <SPLIT distance="600" swimtime="00:09:02.96" />
                    <SPLIT distance="700" swimtime="00:10:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="500" reactiontime="+91" swimtime="00:01:12.77" resultid="3694" heatid="7802" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="541" reactiontime="+93" swimtime="00:01:23.33" resultid="3695" heatid="7834" lane="8" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" status="DNS" swimtime="00:00:00.00" resultid="3696" heatid="7903" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1463" points="507" reactiontime="+91" swimtime="00:02:40.66" resultid="3697" heatid="7949" lane="1" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:17.66" />
                    <SPLIT distance="150" swimtime="00:01:59.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="484" reactiontime="+94" swimtime="00:05:47.68" resultid="3698" heatid="9048" lane="1" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:21.25" />
                    <SPLIT distance="150" swimtime="00:02:06.20" />
                    <SPLIT distance="200" swimtime="00:02:51.47" />
                    <SPLIT distance="250" swimtime="00:03:36.23" />
                    <SPLIT distance="300" swimtime="00:04:21.07" />
                    <SPLIT distance="350" swimtime="00:05:05.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-20" firstname="Robert" gender="M" lastname="Budek" nation="POL" athleteid="3699">
              <RESULTS>
                <RESULT eventid="1076" points="397" reactiontime="+78" swimtime="00:00:32.25" resultid="3700" heatid="7693" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1254" points="303" reactiontime="+95" swimtime="00:01:16.55" resultid="3701" heatid="7812" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="251" reactiontime="+90" swimtime="00:01:33.53" resultid="3702" heatid="7843" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="3703" heatid="7911" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="3704" heatid="7957" lane="1" entrytime="00:02:50.00" />
                <RESULT eventid="1655" points="356" reactiontime="+85" swimtime="00:00:40.73" resultid="3705" heatid="8033" lane="6" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Akademia Ruchu AG B" number="1">
              <RESULTS>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="3708" heatid="7971" lane="7" entrytime="00:02:12.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3674" number="1" />
                    <RELAYPOSITION athleteid="3699" number="2" />
                    <RELAYPOSITION athleteid="3686" number="3" />
                    <RELAYPOSITION athleteid="3669" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start), na trzeciej zmianie" eventid="1357" reactiontime="+81" status="DSQ" swimtime="00:02:34.30" resultid="3709" heatid="7870" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:26.23" />
                    <SPLIT distance="150" swimtime="00:02:01.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3674" number="1" reactiontime="+81" status="DSQ" />
                    <RELAYPOSITION athleteid="3669" number="2" reactiontime="+55" status="DSQ" />
                    <RELAYPOSITION athleteid="3686" number="3" reactiontime="+9" status="DSQ" />
                    <RELAYPOSITION athleteid="3699" number="4" reactiontime="-12" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Akademia Ruchu AG B" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+81" swimtime="00:02:21.34" resultid="3706" heatid="7735" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="150" swimtime="00:01:38.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3686" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3699" number="2" reactiontime="-3" />
                    <RELAYPOSITION athleteid="3692" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3680" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" reactiontime="+84" swimtime="00:02:34.02" resultid="3707" heatid="8050" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:52.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3686" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3669" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="3692" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3680" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ALLST" nation="RUS" clubid="2005" name="All Stars Moscow">
          <ATHLETES>
            <ATHLETE birthdate="1955-04-20" firstname="Ludmila" gender="F" lastname="Lukashova" nation="RUS" athleteid="2006">
              <RESULTS>
                <RESULT eventid="1173" points="289" reactiontime="+78" swimtime="00:00:55.04" resultid="2007" heatid="7754" lane="4" entrytime="00:00:55.00" />
                <RESULT eventid="1270" points="294" reactiontime="+102" swimtime="00:01:56.52" resultid="2008" heatid="7827" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="251" reactiontime="+89" swimtime="00:02:06.35" resultid="2009" heatid="7927" lane="8" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="257" reactiontime="+77" swimtime="00:04:30.82" resultid="2010" heatid="8005" lane="2" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.23" />
                    <SPLIT distance="100" swimtime="00:02:08.99" />
                    <SPLIT distance="150" swimtime="00:03:20.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQLVI" nation="UKR" clubid="4519" name="Aqua Masters SC Kyiv" shortname="Aqua Masters Kyiv">
          <CONTACT city="Kyiv" email="vikup@cyfra.net" name="VIIUK Iurii" phone="+38 050 3314460" street="Mateyuka str. 13, ap. 114" zip="02156" />
          <ATHLETES>
            <ATHLETE birthdate="1959-11-17" firstname="Iurii" gender="M" lastname="Viiuk" nation="UKR" athleteid="4535">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4536" heatid="7699" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="4537" heatid="7817" lane="3" entrytime="00:01:05.00" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="4538" heatid="7890" lane="2" entrytime="00:01:25.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="4539" heatid="8041" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-08-14" firstname="Fedir" gender="M" lastname="Pshenychnyy" nation="UKR" athleteid="4540">
              <RESULTS>
                <RESULT eventid="1076" points="439" reactiontime="+109" swimtime="00:00:35.51" resultid="4541" heatid="7689" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1254" points="370" reactiontime="+119" swimtime="00:01:23.36" resultid="4542" heatid="7809" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="4543" heatid="7955" lane="5" entrytime="00:03:00.00" />
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="4544" heatid="9069" lane="2" entrytime="00:07:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQWRO" nation="POL" region="01" clubid="5800" name="Aquapark Wrocław">
          <CONTACT name="Stasiaczek" phone="792883772" />
          <ATHLETES>
            <ATHLETE birthdate="1984-11-17" firstname="Michał" gender="M" lastname="Stasiaczek" nation="POL" athleteid="5806">
              <RESULTS>
                <RESULT eventid="1108" points="494" reactiontime="+74" swimtime="00:02:32.44" resultid="5807" heatid="7732" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:11.05" />
                    <SPLIT distance="150" swimtime="00:01:53.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="577" reactiontime="+75" swimtime="00:02:46.22" resultid="5808" heatid="7795" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                    <SPLIT distance="100" swimtime="00:01:17.02" />
                    <SPLIT distance="150" swimtime="00:02:00.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="536" reactiontime="+78" swimtime="00:01:07.93" resultid="5809" heatid="7855" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="570" reactiontime="+85" swimtime="00:01:14.77" resultid="5810" heatid="7895" lane="3" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="641" reactiontime="+74" swimtime="00:00:32.77" resultid="5811" heatid="8047" lane="6" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-10-01" firstname="Tomasz" gender="M" lastname="Cimicki" nation="POL" athleteid="5812">
              <RESULTS>
                <RESULT eventid="1383" points="565" reactiontime="+89" swimtime="00:01:14.99" resultid="5813" heatid="7894" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="633" reactiontime="+81" swimtime="00:00:32.91" resultid="5814" heatid="8046" lane="3" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-21" firstname="Mateusz" gender="M" lastname="Dudek" nation="POL" athleteid="5815">
              <RESULTS>
                <RESULT eventid="1222" points="721" reactiontime="+76" swimtime="00:02:34.36" resultid="5816" heatid="7795" lane="5" entrytime="00:02:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                    <SPLIT distance="150" swimtime="00:01:53.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="713" reactiontime="+78" swimtime="00:01:09.41" resultid="5817" heatid="7895" lane="5" entrytime="00:01:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="734" reactiontime="+75" swimtime="00:00:31.32" resultid="5818" heatid="8047" lane="4" entrytime="00:00:30.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-01" firstname="Szymon" gender="M" lastname="Kujat" nation="POL" athleteid="5819">
              <RESULTS>
                <RESULT eventid="1318" points="399" reactiontime="+91" swimtime="00:02:48.40" resultid="5820" heatid="7865" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:12.49" />
                    <SPLIT distance="150" swimtime="00:02:02.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="493" reactiontime="+95" swimtime="00:02:14.80" resultid="5821" heatid="7966" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:04.70" />
                    <SPLIT distance="150" swimtime="00:01:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="413" reactiontime="+88" swimtime="00:01:10.63" resultid="5822" heatid="8001" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-26" firstname="Mateusz" gender="M" lastname="Stawiany" nation="POL" athleteid="5823">
              <RESULTS>
                <RESULT eventid="1108" points="600" reactiontime="+73" swimtime="00:02:22.90" resultid="5824" heatid="7733" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                    <SPLIT distance="100" swimtime="00:01:05.36" />
                    <SPLIT distance="150" swimtime="00:01:46.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="636" reactiontime="+75" swimtime="00:00:56.48" resultid="5825" heatid="7825" lane="1" entrytime="00:00:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="689" reactiontime="+77" swimtime="00:01:02.47" resultid="5826" heatid="7855" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="744" reactiontime="+78" swimtime="00:02:04.17" resultid="5827" heatid="7967" lane="5" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                    <SPLIT distance="100" swimtime="00:00:58.45" />
                    <SPLIT distance="150" swimtime="00:01:30.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-03-09" firstname="Piotr" gender="M" lastname="Rzeczkowski" nation="POL" athleteid="6405">
              <RESULTS>
                <RESULT eventid="1108" points="734" reactiontime="+86" swimtime="00:02:20.76" resultid="6406" heatid="7733" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="100" swimtime="00:01:04.20" />
                    <SPLIT distance="150" swimtime="00:01:47.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="788" reactiontime="+83" swimtime="00:01:02.17" resultid="6407" heatid="7856" lane="2" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="851" reactiontime="+76" swimtime="00:00:26.37" resultid="6408" heatid="7924" lane="5" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="Aquapark Wrocław A" number="1">
              <RESULTS>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="6409" heatid="7872" lane="3" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5819" number="1" />
                    <RELAYPOSITION athleteid="5806" number="2" />
                    <RELAYPOSITION athleteid="5815" number="3" />
                    <RELAYPOSITION athleteid="5823" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="Aquapark Wrocław A" number="2">
              <RESULTS>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="6410" heatid="7973" lane="2" entrytime="00:01:52.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5823" number="1" />
                    <RELAYPOSITION athleteid="5815" number="2" />
                    <RELAYPOSITION athleteid="5819" number="3" />
                    <RELAYPOSITION athleteid="5806" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="CMKRA" nation="POL" region="06" clubid="2079" name="Collegium Medicum UJ Masters Kraków" shortname="CM UJ Masters Kraków">
          <CONTACT city="Kraków" email="MariuszBaranik@gmail.com" name="Mariusz Baranik" phone="698128222" state="MAŁOP" street="Białoprądnicka 32c/3" zip="31-221" />
          <ATHLETES>
            <ATHLETE birthdate="1969-08-22" firstname="Mirosław" gender="M" lastname="Woźniak" nation="POL" athleteid="2087">
              <RESULTS>
                <RESULT eventid="1108" points="464" reactiontime="+79" swimtime="00:02:45.18" resultid="2088" heatid="7727" lane="4" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:16.12" />
                    <SPLIT distance="150" swimtime="00:02:05.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="533" reactiontime="+80" swimtime="00:01:13.75" resultid="2089" heatid="7849" lane="5" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-29" firstname="Mariusz" gender="M" lastname="Baranik" nation="POL" athleteid="2090">
              <RESULTS>
                <RESULT eventid="1076" points="673" reactiontime="+81" swimtime="00:00:27.10" resultid="2091" heatid="7706" lane="3" entrytime="00:00:27.20" entrycourse="SCM" />
                <RESULT eventid="1415" points="623" reactiontime="+85" swimtime="00:00:29.42" resultid="2092" heatid="7920" lane="3" entrytime="00:00:29.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-17" firstname="Wojciech" gender="M" lastname="Liszkowski" nation="POL" athleteid="2093">
              <RESULTS>
                <RESULT eventid="1190" points="626" reactiontime="+75" swimtime="00:00:31.73" resultid="2094" heatid="7772" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-11" firstname="Marcin" gender="M" lastname="Szczurek" nation="POL" athleteid="2095" />
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="2566">
              <RESULTS>
                <RESULT eventid="1059" points="818" reactiontime="+85" swimtime="00:00:28.31" resultid="2567" heatid="7683" lane="4" entrytime="00:00:27.95" />
                <RESULT eventid="1092" points="874" reactiontime="+85" swimtime="00:02:29.57" resultid="2568" heatid="7718" lane="4" entrytime="00:02:30.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:10.83" />
                    <SPLIT distance="150" swimtime="00:01:54.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="865" reactiontime="+85" swimtime="00:01:00.72" resultid="2570" heatid="7805" lane="5" entrytime="00:01:01.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="840" reactiontime="+81" swimtime="00:01:09.00" resultid="2571" heatid="7837" lane="3" entrytime="00:01:08.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="741" reactiontime="+85" swimtime="00:01:19.05" resultid="2572" heatid="7880" lane="5" entrytime="00:01:18.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="805" reactiontime="+85" swimtime="00:02:12.37" resultid="2573" heatid="7951" lane="4" entrytime="00:02:14.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:02.79" />
                    <SPLIT distance="150" swimtime="00:01:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="744" reactiontime="+85" swimtime="00:00:36.23" resultid="2574" heatid="8028" lane="5" entrytime="00:00:35.51" />
                <RESULT eventid="1687" points="722" reactiontime="+86" swimtime="00:04:48.24" resultid="2575" heatid="9047" lane="4" entrytime="00:04:49.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="150" swimtime="00:01:41.38" />
                    <SPLIT distance="200" swimtime="00:02:18.64" />
                    <SPLIT distance="250" swimtime="00:02:56.41" />
                    <SPLIT distance="300" swimtime="00:03:34.54" />
                    <SPLIT distance="350" swimtime="00:04:12.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="CM UJ Ktraków C" number="1">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+75" swimtime="00:02:11.08" resultid="2096" heatid="7871" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="150" swimtime="00:01:43.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2093" number="1" />
                    <RELAYPOSITION athleteid="2095" number="2" />
                    <RELAYPOSITION athleteid="2090" number="3" />
                    <RELAYPOSITION athleteid="2087" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" reactiontime="+86" swimtime="00:01:53.95" resultid="2097" heatid="7973" lane="7" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                    <SPLIT distance="100" swimtime="00:00:59.58" />
                    <SPLIT distance="150" swimtime="00:01:27.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2095" number="1" />
                    <RELAYPOSITION athleteid="2087" number="2" />
                    <RELAYPOSITION athleteid="2093" number="3" />
                    <RELAYPOSITION athleteid="2090" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="FLGDY" nation="POL" region="10" clubid="2044" name="Flota Masters Gdynia">
          <CONTACT city="Gdynia" email="ajot@life.pl" name="JACASZEK Andrzej" phone="697 055 044" state="POM" street="Starowiejska 3/1A" zip="81-356" />
          <ATHLETES>
            <ATHLETE birthdate="1953-01-24" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="2045">
              <RESULTS>
                <RESULT eventid="1076" points="473" reactiontime="+101" swimtime="00:00:34.64" resultid="2046" heatid="7690" lane="8" entrytime="00:00:34.80" entrycourse="SCM" />
                <RESULT eventid="1286" points="433" reactiontime="+98" swimtime="00:01:35.71" resultid="2047" heatid="7841" lane="6" entrytime="00:01:35.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="612" reactiontime="+106" swimtime="00:01:32.02" resultid="2048" heatid="7885" lane="6" entrytime="00:01:38.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="563" reactiontime="+102" swimtime="00:00:40.93" resultid="2049" heatid="8034" lane="5" entrytime="00:00:42.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01610" nation="POL" region="10" clubid="4551" name="GP Gdynia Masters" shortname="Gdynia Masters">
          <CONTACT email="k.mysiak@wpit.am.gdynia.pl" name="mysiak katarzyna" />
          <ATHLETES>
            <ATHLETE birthdate="1959-01-01" firstname="Renata" gender="F" lastname="Polańczyk" nation="POL" athleteid="4552">
              <RESULTS>
                <RESULT eventid="1092" points="322" reactiontime="+103" swimtime="00:03:46.65" resultid="4553" heatid="7715" lane="1" entrytime="00:03:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                    <SPLIT distance="100" swimtime="00:01:41.46" />
                    <SPLIT distance="150" swimtime="00:02:56.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="323" swimtime="00:14:12.43" resultid="4554" heatid="8714" lane="6" entrytime="00:13:38.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:32.96" />
                    <SPLIT distance="200" swimtime="00:03:15.46" />
                    <SPLIT distance="300" swimtime="00:05:01.84" />
                    <SPLIT distance="400" swimtime="00:06:50.12" />
                    <SPLIT distance="500" swimtime="00:08:42.74" />
                    <SPLIT distance="600" swimtime="01:03:31.18" />
                    <SPLIT distance="700" swimtime="00:12:22.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" status="DNS" swimtime="00:00:00.00" resultid="4555" heatid="7756" lane="6" entrytime="00:00:44.02" />
                <RESULT eventid="1302" points="313" reactiontime="+115" swimtime="00:04:10.53" resultid="4556" heatid="7858" lane="7" entrytime="00:03:57.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.41" />
                    <SPLIT distance="100" swimtime="00:01:58.76" />
                    <SPLIT distance="150" swimtime="00:03:04.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" status="DNS" swimtime="00:00:00.00" resultid="4557" heatid="7927" lane="5" entrytime="00:01:35.46" />
                <RESULT eventid="1527" points="340" reactiontime="+109" swimtime="00:08:01.16" resultid="4558" heatid="8803" lane="1" entrytime="00:08:02.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.59" />
                    <SPLIT distance="100" swimtime="00:01:56.92" />
                    <SPLIT distance="150" swimtime="00:02:52.43" />
                    <SPLIT distance="200" swimtime="00:03:45.76" />
                    <SPLIT distance="250" swimtime="00:05:01.05" />
                    <SPLIT distance="300" swimtime="00:06:17.48" />
                    <SPLIT distance="350" swimtime="00:07:11.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" status="DNS" swimtime="00:00:00.00" resultid="4559" heatid="8006" lane="1" entrytime="00:03:25.36" />
                <RESULT eventid="1687" status="DNS" swimtime="00:00:00.00" resultid="4560" heatid="9052" lane="4" entrytime="00:06:42.18" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Katarzyna" gender="F" lastname="Mysiak" nation="POL" athleteid="4561">
              <RESULTS>
                <RESULT eventid="1140" points="307" swimtime="00:14:27.10" resultid="4562" heatid="8714" lane="2" entrytime="00:13:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:33.48" />
                    <SPLIT distance="200" swimtime="00:03:18.44" />
                    <SPLIT distance="300" swimtime="00:05:08.05" />
                    <SPLIT distance="400" swimtime="00:07:00.30" />
                    <SPLIT distance="500" swimtime="00:08:53.03" />
                    <SPLIT distance="600" swimtime="00:10:46.04" />
                    <SPLIT distance="700" swimtime="00:12:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="362" reactiontime="+78" swimtime="00:00:46.58" resultid="4563" heatid="7756" lane="5" entrytime="00:00:44.00" />
                <RESULT eventid="1238" points="338" reactiontime="+102" swimtime="00:01:28.89" resultid="4564" heatid="7799" lane="6" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="304" reactiontime="+107" swimtime="00:03:20.54" resultid="4565" heatid="7947" lane="1" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                    <SPLIT distance="100" swimtime="00:01:34.36" />
                    <SPLIT distance="150" swimtime="00:02:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="328" reactiontime="+101" swimtime="00:06:54.92" resultid="4566" heatid="9051" lane="1" entrytime="00:06:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                    <SPLIT distance="100" swimtime="00:01:34.54" />
                    <SPLIT distance="150" swimtime="00:02:26.63" />
                    <SPLIT distance="200" swimtime="00:03:19.72" />
                    <SPLIT distance="250" swimtime="00:04:13.63" />
                    <SPLIT distance="300" swimtime="00:05:08.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="4567">
              <RESULTS>
                <RESULT eventid="1076" points="443" reactiontime="+104" swimtime="00:00:38.03" resultid="4568" heatid="7687" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1108" points="470" reactiontime="+108" swimtime="00:03:48.57" resultid="4569" heatid="7721" lane="7" entrytime="00:03:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.86" />
                    <SPLIT distance="100" swimtime="00:01:50.10" />
                    <SPLIT distance="150" swimtime="00:02:53.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="385" reactiontime="+86" swimtime="00:00:47.64" resultid="4570" heatid="7766" lane="6" entrytime="00:00:46.00" />
                <RESULT eventid="1222" points="454" reactiontime="+106" swimtime="00:04:00.92" resultid="4571" heatid="7787" lane="1" entrytime="00:03:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.25" />
                    <SPLIT distance="100" swimtime="00:01:52.99" />
                    <SPLIT distance="150" swimtime="00:02:57.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="536" reactiontime="+99" swimtime="00:01:43.03" resultid="4572" heatid="7884" lane="1" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="378" reactiontime="+108" swimtime="00:00:45.23" resultid="4573" heatid="7908" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1591" points="383" reactiontime="+99" swimtime="00:01:51.57" resultid="4574" heatid="7994" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="592" reactiontime="+106" swimtime="00:00:44.57" resultid="4575" heatid="8034" lane="7" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="4576">
              <RESULTS>
                <RESULT eventid="1190" points="544" reactiontime="+81" swimtime="00:00:48.86" resultid="4577" heatid="7766" lane="7" entrytime="00:00:47.10" />
                <RESULT eventid="1222" points="474" reactiontime="+107" swimtime="00:04:10.70" resultid="4578" heatid="7787" lane="6" entrytime="00:03:46.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.62" />
                    <SPLIT distance="100" swimtime="00:02:02.38" />
                    <SPLIT distance="150" swimtime="00:03:08.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="477" reactiontime="+103" swimtime="00:01:50.99" resultid="4579" heatid="7883" lane="5" entrytime="00:01:44.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="519" reactiontime="+111" swimtime="00:00:48.76" resultid="4580" heatid="8032" lane="7" entrytime="00:00:46.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="Mikołajczyk" nation="POL" athleteid="4581">
              <RESULTS>
                <RESULT eventid="1108" points="481" reactiontime="+97" swimtime="00:03:29.58" resultid="4582" heatid="7722" lane="1" entrytime="00:03:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.12" />
                    <SPLIT distance="100" swimtime="00:01:45.15" />
                    <SPLIT distance="150" swimtime="00:02:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="516" reactiontime="+97" swimtime="00:03:38.09" resultid="4583" heatid="7788" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.27" />
                    <SPLIT distance="100" swimtime="00:01:44.97" />
                    <SPLIT distance="150" swimtime="00:02:41.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="339" reactiontime="+99" swimtime="00:03:48.96" resultid="4584" heatid="7861" lane="6" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:49.31" />
                    <SPLIT distance="150" swimtime="00:02:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="477" reactiontime="+100" swimtime="00:01:39.99" resultid="4585" heatid="7885" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="WDR" swimtime="00:00:00.00" resultid="4586" entrytime="00:07:36.00" />
                <RESULT eventid="1591" points="277" reactiontime="+102" swimtime="00:01:44.77" resultid="4587" heatid="7993" lane="5" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="428" reactiontime="+96" swimtime="00:00:44.83" resultid="4588" heatid="8033" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Piotr" gender="M" lastname="Stasiuk" nation="POL" athleteid="4589">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="4590" heatid="7727" lane="2" entrytime="00:02:52.00" />
                <RESULT eventid="1286" status="WDR" swimtime="00:00:00.00" resultid="4591" heatid="7848" lane="5" entrytime="00:01:15.00" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="4592" heatid="7915" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1591" status="WDR" swimtime="00:00:00.00" resultid="4593" heatid="7998" lane="5" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Grażyna" gender="F" lastname="Heisler" nation="POL" athleteid="4594">
              <RESULTS>
                <RESULT eventid="1059" points="337" reactiontime="+110" swimtime="00:00:46.16" resultid="4595" heatid="7673" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1270" points="303" reactiontime="+91" swimtime="00:01:57.71" resultid="4596" heatid="7827" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="298" reactiontime="+96" swimtime="00:02:09.29" resultid="4597" heatid="7874" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" status="DNS" swimtime="00:00:00.00" resultid="4598" heatid="8023" lane="5" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Hanka" gender="F" lastname="Kania" nation="POL" athleteid="4599">
              <RESULTS>
                <RESULT eventid="1059" status="WDR" swimtime="00:00:00.00" resultid="4600" heatid="7675" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1092" points="453" reactiontime="+107" swimtime="00:03:42.64" resultid="4601" heatid="7714" lane="3" entrytime="00:04:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.14" />
                    <SPLIT distance="100" swimtime="00:01:48.71" />
                    <SPLIT distance="150" swimtime="00:02:51.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="493" reactiontime="+107" swimtime="00:03:54.45" resultid="4602" heatid="7780" lane="4" entrytime="00:03:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.22" />
                    <SPLIT distance="100" swimtime="00:01:51.84" />
                    <SPLIT distance="150" swimtime="00:02:53.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" status="WDR" swimtime="00:00:00.00" resultid="4603" heatid="7829" lane="8" entrytime="00:01:42.00" />
                <RESULT eventid="1366" points="407" reactiontime="+108" swimtime="00:01:52.87" resultid="4604" heatid="7875" lane="4" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" status="DNS" swimtime="00:00:00.00" resultid="4605" heatid="7898" lane="3" entrytime="00:00:48.00" />
                <RESULT eventid="1574" points="358" reactiontime="+110" swimtime="00:01:50.78" resultid="4606" heatid="7988" lane="1" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" status="WDR" swimtime="00:00:00.00" resultid="4607" heatid="8022" lane="3" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Leszek" gender="M" lastname="Kubicki" nation="POL" athleteid="4608">
              <RESULTS>
                <RESULT eventid="1076" points="605" reactiontime="+94" swimtime="00:00:31.92" resultid="4609" heatid="7691" lane="2" entrytime="00:00:33.03" />
                <RESULT eventid="1156" points="829" swimtime="00:22:45.01" resultid="4610" heatid="8720" lane="3" entrytime="00:22:19.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:01:20.80" />
                    <SPLIT distance="200" swimtime="00:02:51.34" />
                    <SPLIT distance="300" swimtime="00:04:22.38" />
                    <SPLIT distance="400" swimtime="00:05:53.34" />
                    <SPLIT distance="500" swimtime="00:07:24.11" />
                    <SPLIT distance="600" swimtime="00:08:54.80" />
                    <SPLIT distance="700" swimtime="00:10:25.01" />
                    <SPLIT distance="800" swimtime="00:11:56.82" />
                    <SPLIT distance="900" swimtime="00:13:28.55" />
                    <SPLIT distance="1000" swimtime="00:15:00.56" />
                    <SPLIT distance="1100" swimtime="00:16:33.75" />
                    <SPLIT distance="1200" swimtime="00:18:06.94" />
                    <SPLIT distance="1300" swimtime="00:19:40.50" />
                    <SPLIT distance="1400" swimtime="00:21:14.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="565" reactiontime="+98" swimtime="00:03:31.60" resultid="4611" heatid="7790" lane="7" entrytime="00:03:24.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                    <SPLIT distance="100" swimtime="00:01:39.48" />
                    <SPLIT distance="150" swimtime="00:02:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="550" reactiontime="+107" swimtime="00:01:28.40" resultid="4612" heatid="7843" lane="3" entrytime="00:01:25.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="602" reactiontime="+94" swimtime="00:02:43.22" resultid="4613" heatid="7958" lane="5" entrytime="00:02:41.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:16.29" />
                    <SPLIT distance="150" swimtime="00:02:00.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="4614" heatid="8029" lane="2" />
                <RESULT eventid="1703" points="559" reactiontime="+109" swimtime="00:06:05.20" resultid="4615" heatid="9065" lane="5" entrytime="00:05:34.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:20.85" />
                    <SPLIT distance="150" swimtime="00:02:12.46" />
                    <SPLIT distance="200" swimtime="00:02:57.92" />
                    <SPLIT distance="250" swimtime="00:03:44.72" />
                    <SPLIT distance="300" swimtime="00:04:31.93" />
                    <SPLIT distance="350" swimtime="00:05:19.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Katarzyna" gender="F" lastname="Mazurek" nation="POL" athleteid="4616">
              <RESULTS>
                <RESULT eventid="1059" points="481" reactiontime="+98" swimtime="00:00:36.37" resultid="4617" heatid="7678" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1238" points="418" reactiontime="+94" swimtime="00:01:22.81" resultid="4618" heatid="7800" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="483" reactiontime="+97" swimtime="00:01:32.53" resultid="4619" heatid="7832" lane="5" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="526" reactiontime="+96" swimtime="00:01:39.35" resultid="4620" heatid="7878" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="424" reactiontime="+98" swimtime="00:00:41.45" resultid="4621" heatid="7899" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1574" points="362" reactiontime="+96" swimtime="00:01:39.27" resultid="4622" heatid="7989" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="575" reactiontime="+97" swimtime="00:00:44.06" resultid="4623" heatid="8026" lane="4" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Danuta" gender="F" lastname="Radkowiak" nation="POL" athleteid="4624">
              <RESULTS>
                <RESULT eventid="1092" points="266" reactiontime="+100" swimtime="00:04:01.44" resultid="4625" heatid="7715" lane="8" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                    <SPLIT distance="100" swimtime="00:02:02.13" />
                    <SPLIT distance="150" swimtime="00:03:07.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="355" reactiontime="+108" swimtime="00:04:10.54" resultid="4626" heatid="7779" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.61" />
                    <SPLIT distance="100" swimtime="00:02:02.23" />
                    <SPLIT distance="150" swimtime="00:03:07.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="4627" heatid="7857" lane="5" entrytime="00:08:00.00" />
                <RESULT eventid="1527" status="DNS" swimtime="00:00:00.00" resultid="4628" heatid="8802" lane="5" entrytime="00:08:00.00" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="4629" heatid="7988" lane="2" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Masters Gdynia E" number="1">
              <RESULTS>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="4633" heatid="7868" lane="6" entrytime="00:03:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4567" number="1" />
                    <RELAYPOSITION athleteid="4576" number="2" />
                    <RELAYPOSITION athleteid="4581" number="3" />
                    <RELAYPOSITION athleteid="4589" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="4634" heatid="7970" lane="2" entrytime="00:03:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4576" number="1" />
                    <RELAYPOSITION athleteid="4608" number="2" />
                    <RELAYPOSITION athleteid="4567" number="3" />
                    <RELAYPOSITION athleteid="4589" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Masters Gdynia D" number="1">
              <RESULTS>
                <RESULT eventid="1334" reactiontime="+73" swimtime="00:02:56.06" resultid="4631" heatid="7866" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                    <SPLIT distance="100" swimtime="00:01:30.22" />
                    <SPLIT distance="150" swimtime="00:02:16.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4552" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4616" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4561" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4624" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1495" reactiontime="+114" swimtime="00:02:42.63" resultid="4635" heatid="7968" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:22.77" />
                    <SPLIT distance="150" swimtime="00:02:03.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4552" number="1" />
                    <RELAYPOSITION athleteid="4561" number="2" />
                    <RELAYPOSITION athleteid="4624" number="3" />
                    <RELAYPOSITION athleteid="4616" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Masters Gdynia D" number="1">
              <RESULTS>
                <RESULT eventid="1671" status="WDR" swimtime="00:00:00.00" resultid="4630" heatid="8049" lane="5" entrytime="00:03:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4561" number="1" />
                    <RELAYPOSITION athleteid="4567" number="2" />
                    <RELAYPOSITION athleteid="4581" number="3" />
                    <RELAYPOSITION athleteid="4616" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Masters Gdynia E" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+99" swimtime="00:02:24.85" resultid="4632" heatid="7734" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4608" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="4561" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="4567" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4616" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02210" nation="POL" region="10" clubid="5168" name="GP Sopot Masters" shortname="Sopot Masters">
          <CONTACT city="Sopot" email="puchalskaasia@wp.pl" name="Puchalska" phone="607035439" state="POM" street="Hallera 57" zip="81-715" />
          <ATHLETES>
            <ATHLETE birthdate="1964-08-04" firstname="Joanna" gender="F" lastname="Puchalska" nation="POL" athleteid="5169">
              <RESULTS>
                <RESULT eventid="1092" points="786" reactiontime="+85" swimtime="00:02:45.71" resultid="5170" heatid="7718" lane="8" entrytime="00:02:49.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="150" swimtime="00:02:06.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="830" reactiontime="+91" swimtime="00:03:01.33" resultid="5171" heatid="7783" lane="1" entrytime="00:03:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                    <SPLIT distance="100" swimtime="00:01:28.70" />
                    <SPLIT distance="150" swimtime="00:02:15.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="804" reactiontime="+85" swimtime="00:01:24.81" resultid="5172" heatid="7879" lane="5" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="710" reactiontime="+95" swimtime="00:00:33.65" resultid="5173" heatid="7904" lane="2" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1527" points="831" reactiontime="+93" swimtime="00:05:48.31" resultid="5174" heatid="8802" lane="4" entrytime="00:05:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:18.65" />
                    <SPLIT distance="150" swimtime="00:02:05.53" />
                    <SPLIT distance="200" swimtime="00:02:51.08" />
                    <SPLIT distance="250" swimtime="00:03:39.41" />
                    <SPLIT distance="300" swimtime="00:04:27.91" />
                    <SPLIT distance="350" swimtime="00:05:09.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="764" reactiontime="+84" swimtime="00:01:14.43" resultid="5175" heatid="7991" lane="3" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-08" firstname="Anna" gender="F" lastname="Maciejowska" nation="POL" athleteid="5176">
              <RESULTS>
                <RESULT eventid="1173" points="466" reactiontime="+81" swimtime="00:00:42.81" resultid="5177" heatid="7757" lane="5" entrytime="00:00:41.50" entrycourse="SCM" />
                <RESULT eventid="1238" points="459" reactiontime="+80" swimtime="00:01:20.31" resultid="5178" heatid="7800" lane="4" entrytime="00:01:21.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="480" reactiontime="+77" swimtime="00:00:39.76" resultid="5179" heatid="7900" lane="7" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1463" points="434" reactiontime="+86" swimtime="00:02:58.14" resultid="5180" heatid="7947" lane="4" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:24.52" />
                    <SPLIT distance="150" swimtime="00:02:11.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-12-28" firstname="Dariusz" gender="M" lastname="Gorbaczow" nation="POL" athleteid="5181">
              <RESULTS>
                <RESULT eventid="1076" points="743" reactiontime="+81" swimtime="00:00:28.79" resultid="5182" heatid="7697" lane="2" entrytime="00:00:30.10" entrycourse="SCM" />
                <RESULT eventid="1190" points="823" reactiontime="+81" swimtime="00:00:33.58" resultid="5183" heatid="7773" lane="3" entrytime="00:00:33.90" entrycourse="SCM" />
                <RESULT eventid="1286" points="847" reactiontime="+93" swimtime="00:01:13.10" resultid="5184" heatid="7849" lane="8" entrytime="00:01:14.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="825" reactiontime="+79" swimtime="00:00:30.40" resultid="5185" heatid="7916" lane="8" entrytime="00:00:32.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="HTKRA" nation="POL" region="06" clubid="6441" name="Happy TRI Friends Kraków">
          <ATHLETES>
            <ATHLETE birthdate="1973-04-13" firstname="Marcin" gender="M" lastname="Lewandowski" nation="POL" athleteid="6186">
              <RESULTS>
                <RESULT eventid="1156" points="416" swimtime="00:22:15.35" resultid="6187" heatid="8720" lane="6" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="100" swimtime="00:01:22.18" />
                    <SPLIT distance="200" swimtime="00:02:48.76" />
                    <SPLIT distance="300" swimtime="00:04:17.76" />
                    <SPLIT distance="400" swimtime="00:05:47.90" />
                    <SPLIT distance="500" swimtime="00:07:17.94" />
                    <SPLIT distance="600" swimtime="00:08:47.92" />
                    <SPLIT distance="700" swimtime="00:10:17.69" />
                    <SPLIT distance="800" swimtime="00:11:47.90" />
                    <SPLIT distance="900" swimtime="00:13:18.59" />
                    <SPLIT distance="1000" swimtime="00:14:48.83" />
                    <SPLIT distance="1100" swimtime="00:16:18.68" />
                    <SPLIT distance="1200" swimtime="00:17:49.36" />
                    <SPLIT distance="1300" swimtime="00:19:19.59" />
                    <SPLIT distance="1400" swimtime="00:20:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="416" reactiontime="+90" swimtime="00:02:31.34" resultid="6188" heatid="7957" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:53.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="408" reactiontime="+86" swimtime="00:05:24.44" resultid="6189" heatid="9066" lane="5" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="150" swimtime="00:01:57.60" />
                    <SPLIT distance="200" swimtime="00:02:39.16" />
                    <SPLIT distance="250" swimtime="00:03:21.41" />
                    <SPLIT distance="300" swimtime="00:04:03.85" />
                    <SPLIT distance="350" swimtime="00:04:45.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="IKKON" nation="POL" region="14" clubid="6132" name="IKS Konstancin">
          <CONTACT email="rafal@juchno.com" name="Juchno" phone="691-440-213" />
          <ATHLETES>
            <ATHLETE birthdate="1976-10-03" firstname="Rafał" gender="M" lastname="Juchno" nation="POL" athleteid="6133">
              <RESULTS>
                <RESULT eventid="1076" points="533" reactiontime="+101" swimtime="00:00:29.25" resultid="6134" heatid="7699" lane="5" entrytime="00:00:29.59" />
                <RESULT eventid="1254" points="448" reactiontime="+105" swimtime="00:01:07.19" resultid="6135" heatid="7815" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="372" reactiontime="+101" swimtime="00:01:28.96" resultid="6136" heatid="7888" lane="2" entrytime="00:01:29.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="6137" heatid="8038" lane="5" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="IGMLA" nation="POL" region="14" clubid="4545" name="Igan Mława">
          <CONTACT city="Mława" email="ewaszlagor@o2.pl" name="Szlagor" phone="609621127" state="MAZ" street="Żwirki 30" zip="06-500" />
          <ATHLETES>
            <ATHLETE birthdate="1971-12-24" firstname="Ewa" gender="F" lastname="Szlagor" nation="POL" athleteid="4546">
              <RESULTS>
                <RESULT eventid="1059" points="819" reactiontime="+80" swimtime="00:00:29.04" resultid="4547" heatid="7683" lane="1" entrytime="00:00:29.30" entrycourse="SCM" />
                <RESULT eventid="1270" status="DNS" swimtime="00:00:00.00" resultid="4548" heatid="7826" lane="6" />
                <RESULT eventid="1399" points="918" reactiontime="+81" swimtime="00:00:30.73" resultid="4549" heatid="7905" lane="5" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1639" points="899" reactiontime="+82" swimtime="00:00:35.58" resultid="4550" heatid="8020" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="JW2399" nation="POL" region="01" clubid="2305" name="JW 2399 Świętosżów">
          <CONTACT city="Świdnica" email="horbacz.marcin@wp.pl" name="Horbacz Marcin" phone="603672717" state="DOL" street="Buchałów" zip="66-008" />
          <ATHLETES>
            <ATHLETE birthdate="1974-06-16" firstname="Marcin" gender="M" lastname="Horbacz" nation="POL" athleteid="2306">
              <RESULTS>
                <RESULT eventid="1076" points="748" reactiontime="+79" swimtime="00:00:26.13" resultid="2307" heatid="7684" lane="6" entrytime="00:03:00.00" entrycourse="SCM" />
                <RESULT eventid="1108" points="799" reactiontime="+85" swimtime="00:02:17.17" resultid="2308" heatid="7733" lane="7" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:45.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="770" reactiontime="+77" swimtime="00:00:56.10" resultid="2309" heatid="7806" lane="3" entrytime="00:04:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="758" reactiontime="+76" swimtime="00:01:04.74" resultid="2310" heatid="7854" lane="1" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="794" reactiontime="+72" swimtime="00:02:00.34" resultid="2311" heatid="7952" lane="2" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                    <SPLIT distance="100" swimtime="00:00:59.42" />
                    <SPLIT distance="150" swimtime="00:01:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="818" reactiontime="+77" swimtime="00:04:51.80" resultid="2312" heatid="8806" lane="5" entrytime="00:05:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:04.55" />
                    <SPLIT distance="150" swimtime="00:01:44.45" />
                    <SPLIT distance="200" swimtime="00:02:23.47" />
                    <SPLIT distance="250" swimtime="00:03:04.20" />
                    <SPLIT distance="300" swimtime="00:03:45.32" />
                    <SPLIT distance="350" swimtime="00:04:19.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="709" reactiontime="+88" swimtime="00:01:03.74" resultid="2313" heatid="7992" lane="6" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="796" reactiontime="+81" swimtime="00:04:21.42" resultid="2314" heatid="9059" lane="7" entrytime="00:04:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:04.84" />
                    <SPLIT distance="150" swimtime="00:01:38.68" />
                    <SPLIT distance="200" swimtime="00:02:12.25" />
                    <SPLIT distance="250" swimtime="00:02:45.61" />
                    <SPLIT distance="300" swimtime="00:03:18.40" />
                    <SPLIT distance="350" swimtime="00:03:50.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-14" firstname="Jarosław" gender="M" lastname="Druciarek" nation="POL" athleteid="2315">
              <RESULTS>
                <RESULT eventid="1076" points="469" reactiontime="+90" swimtime="00:00:29.39" resultid="2316" heatid="7699" lane="7" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1254" points="370" reactiontime="+79" swimtime="00:01:07.61" resultid="2317" heatid="7807" lane="8" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="2318" heatid="7910" lane="7" entrytime="00:00:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-12-15" firstname="Oscar" gender="M" lastname="Bogucki" nation="POL" athleteid="2319">
              <RESULTS>
                <RESULT eventid="1076" points="400" reactiontime="+77" swimtime="00:00:32.17" resultid="2320" heatid="7693" lane="7" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1222" points="381" reactiontime="+87" swimtime="00:03:16.46" resultid="2321" heatid="7792" lane="1" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="150" swimtime="00:02:23.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="439" reactiontime="+89" swimtime="00:01:24.23" resultid="2322" heatid="7891" lane="6" entrytime="00:01:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="483" reactiontime="+83" swimtime="00:00:36.79" resultid="2323" heatid="8041" lane="4" entrytime="00:00:36.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-29" firstname="Radosław" gender="M" lastname="Stępień" nation="POL" athleteid="2324">
              <RESULTS>
                <RESULT eventid="1076" points="537" reactiontime="+67" swimtime="00:00:28.10" resultid="2325" heatid="7703" lane="6" entrytime="00:00:28.90" entrycourse="SCM" />
                <RESULT eventid="1254" points="415" reactiontime="+63" swimtime="00:01:05.12" resultid="2326" heatid="7816" lane="6" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="309" reactiontime="+71" swimtime="00:01:31.70" resultid="2327" heatid="7886" lane="1" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-11-04" firstname="Mariusz" gender="M" lastname="Janowski" nation="POL" athleteid="2328">
              <RESULTS>
                <RESULT eventid="1076" points="447" reactiontime="+80" swimtime="00:00:28.93" resultid="2329" heatid="7695" lane="4" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1222" points="379" reactiontime="+83" swimtime="00:03:14.13" resultid="2330" heatid="7791" lane="4" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:29.76" />
                    <SPLIT distance="150" swimtime="00:02:21.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="375" reactiontime="+87" swimtime="00:01:25.03" resultid="2331" heatid="7889" lane="5" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="412" reactiontime="+87" swimtime="00:00:37.35" resultid="2332" heatid="8041" lane="1" entrytime="00:00:37.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-27" firstname="Natalia" gender="F" lastname="Szczęsnowicz" nation="POL" athleteid="2333">
              <RESULTS>
                <RESULT eventid="1059" points="524" reactiontime="+79" swimtime="00:00:32.88" resultid="2334" heatid="7681" lane="1" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1238" points="414" reactiontime="+73" swimtime="00:01:18.30" resultid="2335" heatid="7801" lane="5" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="JW 2399 Świętoszów B" number="1">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+65" swimtime="00:02:13.29" resultid="2336" heatid="7870" lane="2" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="150" swimtime="00:01:43.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2306" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2319" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2324" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2315" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1511" reactiontime="+71" status="DSQ" swimtime="00:01:51.89" resultid="2337" heatid="7972" lane="3" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="100" swimtime="00:00:57.66" />
                    <SPLIT distance="150" swimtime="00:01:26.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2324" number="1" />
                    <RELAYPOSITION athleteid="2315" number="2" />
                    <RELAYPOSITION athleteid="2328" number="3" />
                    <RELAYPOSITION athleteid="2306" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="JW4408" nation="POL" region="04" clubid="6783" name="JW 4408 Sulechów">
          <ATHLETES>
            <ATHLETE birthdate="1987-07-18" firstname="Kamila" gender="F" lastname="Szymkowiak" nation="POL" athleteid="2920">
              <RESULTS>
                <RESULT eventid="1059" points="591" reactiontime="+88" swimtime="00:00:31.60" resultid="2921" heatid="7681" lane="6" entrytime="00:00:31.70" />
                <RESULT comment="G2 - Całkowite zanurzenie w trakcie wyścigu (za wyjątkiem 15 m po starcie lub nawrocie)  (Czas: 9:19)" eventid="1173" reactiontime="+72" status="DSQ" swimtime="00:00:35.87" resultid="2922" heatid="7759" lane="5" entrytime="00:00:36.50" />
                <RESULT eventid="1431" points="534" reactiontime="+84" swimtime="00:01:18.59" resultid="2923" heatid="7930" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="398" reactiontime="+82" swimtime="00:03:05.38" resultid="2924" heatid="8008" lane="3" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                    <SPLIT distance="150" swimtime="00:02:17.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="JELGA" nation="LAT" clubid="1891" name="Jelgava SPS">
          <ATHLETES>
            <ATHLETE birthdate="1974-10-14" firstname="Valerijs" gender="M" lastname="Minakovs" nation="LAT" athleteid="1898">
              <RESULTS>
                <RESULT eventid="1108" points="737" reactiontime="+76" swimtime="00:02:20.89" resultid="1899" heatid="7733" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                    <SPLIT distance="100" swimtime="00:01:03.81" />
                    <SPLIT distance="150" swimtime="00:01:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="891" reactiontime="+69" swimtime="00:00:28.20" resultid="1900" heatid="7777" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="1286" points="792" reactiontime="+79" swimtime="00:01:03.80" resultid="1901" heatid="7856" lane="8" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="927" reactiontime="+76" swimtime="00:01:00.63" resultid="1902" heatid="7942" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="930" reactiontime="+71" swimtime="00:02:13.16" resultid="1903" heatid="8019" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="100" swimtime="00:01:03.37" />
                    <SPLIT distance="150" swimtime="00:01:38.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-21" firstname="Jaroslavs" gender="M" lastname="Orbidans" nation="LAT" athleteid="1904">
              <RESULTS>
                <RESULT eventid="1076" points="707" reactiontime="+72" swimtime="00:00:24.84" resultid="1905" heatid="7712" lane="6" entrytime="00:00:24.98" />
                <RESULT eventid="1254" points="697" reactiontime="+70" swimtime="00:00:55.29" resultid="1906" heatid="7824" lane="3" entrytime="00:00:56.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="694" reactiontime="+73" swimtime="00:02:20.03" resultid="1907" heatid="7865" lane="5" entrytime="00:02:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:06.85" />
                    <SPLIT distance="150" swimtime="00:01:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="663" reactiontime="+73" swimtime="00:00:26.22" resultid="1908" heatid="7925" lane="7" entrytime="00:00:26.70" />
                <RESULT eventid="1543" points="670" reactiontime="+77" swimtime="00:05:05.07" resultid="1909" heatid="8806" lane="3" entrytime="00:05:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:08.01" />
                    <SPLIT distance="150" swimtime="00:01:46.65" />
                    <SPLIT distance="200" swimtime="00:02:25.78" />
                    <SPLIT distance="250" swimtime="00:03:09.60" />
                    <SPLIT distance="300" swimtime="00:03:55.20" />
                    <SPLIT distance="350" swimtime="00:04:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="701" reactiontime="+70" swimtime="00:00:59.24" resultid="1910" heatid="8003" lane="1" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01202" nation="POL" region="02" clubid="1875" name="KP Delfin Inowrocław" shortname="Delfin Inowrocław">
          <CONTACT city="Inowrocław" email="jarek.molenda@gmail.com" name="Molenda Jarosław" phone="660899358" state="KUJ" street="Wierzbińskiego 11" zip="88-100" />
          <ATHLETES>
            <ATHLETE birthdate="1937-09-19" firstname="Zygmunt" gender="M" lastname="Lewandowski" nation="POL" license="M01202200038" athleteid="1876">
              <RESULTS>
                <RESULT eventid="1156" points="585" swimtime="00:28:30.20" resultid="1877" heatid="8724" lane="2" entrytime="00:30:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.04" />
                    <SPLIT distance="100" swimtime="00:01:45.37" />
                    <SPLIT distance="200" swimtime="00:03:38.73" />
                    <SPLIT distance="300" swimtime="00:04:35.18" />
                    <SPLIT distance="400" swimtime="00:06:28.36" />
                    <SPLIT distance="500" swimtime="00:08:23.32" />
                    <SPLIT distance="600" swimtime="00:10:17.76" />
                    <SPLIT distance="700" swimtime="00:12:12.53" />
                    <SPLIT distance="800" swimtime="00:14:07.36" />
                    <SPLIT distance="900" swimtime="00:16:04.77" />
                    <SPLIT distance="1000" swimtime="00:18:00.35" />
                    <SPLIT distance="1100" swimtime="00:19:56.39" />
                    <SPLIT distance="1200" swimtime="00:21:52.84" />
                    <SPLIT distance="1300" swimtime="00:23:48.18" />
                    <SPLIT distance="1400" swimtime="00:25:43.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="457" reactiontime="+108" swimtime="00:01:48.39" resultid="1878" heatid="7840" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="400" reactiontime="+107" swimtime="00:00:50.43" resultid="1879" heatid="7907" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1479" points="472" reactiontime="+103" swimtime="00:03:24.16" resultid="1880" heatid="7953" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:39.36" />
                    <SPLIT distance="150" swimtime="00:02:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="455" reactiontime="+106" swimtime="00:01:59.67" resultid="1881" heatid="7992" lane="5" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="1882" entrytime="00:07:16.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-28" firstname="Krzysztof" gender="M" lastname="Derkowski" nation="POL" license="M01202200043" athleteid="1883">
              <RESULTS>
                <RESULT eventid="1076" points="453" reactiontime="+77" swimtime="00:00:33.07" resultid="1884" heatid="7690" lane="4" entrytime="00:00:33.40" />
                <RESULT eventid="1190" points="239" reactiontime="+75" swimtime="00:00:47.33" resultid="1885" heatid="7766" lane="2" entrytime="00:00:46.00" />
                <RESULT eventid="1286" points="399" reactiontime="+79" swimtime="00:01:28.92" resultid="1886" heatid="7842" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="400" reactiontime="+76" swimtime="00:01:34.36" resultid="1887" heatid="7887" lane="5" entrytime="00:01:31.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="419" reactiontime="+88" swimtime="00:00:36.81" resultid="1888" heatid="7912" lane="8" entrytime="00:00:36.40" />
                <RESULT eventid="1655" points="468" reactiontime="+80" swimtime="00:00:40.39" resultid="1889" heatid="8037" lane="1" entrytime="00:00:40.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KPKOZ" nation="POL" region="15" clubid="3034" name="KP Koziegłowy">
          <CONTACT city="Koziegłowy" email="ewaszala59@wp.pl" name="Ewa Szała" street="Osiedle Leśne 13/21" zip="62-028" />
          <ATHLETES>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="3035">
              <RESULTS>
                <RESULT eventid="1092" points="670" reactiontime="+95" swimtime="00:02:57.47" resultid="3036" heatid="7716" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:23.52" />
                    <SPLIT distance="150" swimtime="00:02:15.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="517" swimtime="00:12:08.88" resultid="3037" heatid="8713" lane="2" entrytime="00:12:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:24.15" />
                    <SPLIT distance="200" swimtime="00:02:55.34" />
                    <SPLIT distance="300" swimtime="00:04:27.07" />
                    <SPLIT distance="400" swimtime="00:05:58.71" />
                    <SPLIT distance="500" swimtime="00:07:30.13" />
                    <SPLIT distance="600" swimtime="00:09:02.67" />
                    <SPLIT distance="700" swimtime="00:10:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="689" reactiontime="+90" swimtime="00:01:22.21" resultid="3039" heatid="7833" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="616" reactiontime="+89" swimtime="00:01:24.87" resultid="3040" heatid="7930" lane="8" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="571" reactiontime="+95" swimtime="00:06:44.73" resultid="3041" heatid="8802" lane="2" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                    <SPLIT distance="100" swimtime="00:01:37.59" />
                    <SPLIT distance="150" swimtime="00:02:28.37" />
                    <SPLIT distance="200" swimtime="00:03:18.84" />
                    <SPLIT distance="250" swimtime="00:04:15.39" />
                    <SPLIT distance="300" swimtime="00:05:12.76" />
                    <SPLIT distance="350" swimtime="00:05:59.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="614" reactiontime="+88" swimtime="00:03:05.21" resultid="3042" heatid="8007" lane="4" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="519" reactiontime="+90" swimtime="00:05:56.22" resultid="3043" heatid="9049" lane="7" entrytime="00:05:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:22.90" />
                    <SPLIT distance="150" swimtime="00:02:08.19" />
                    <SPLIT distance="200" swimtime="00:02:54.94" />
                    <SPLIT distance="250" swimtime="00:03:40.32" />
                    <SPLIT distance="300" swimtime="00:04:26.21" />
                    <SPLIT distance="350" swimtime="00:05:12.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="568" reactiontime="+94" swimtime="00:01:14.81" resultid="6404" heatid="7802" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="3044">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="3045" heatid="7724" lane="4" entrytime="00:03:10.00" />
                <RESULT eventid="1156" status="WDR" swimtime="00:00:00.00" resultid="3046" entrytime="00:24:26.00" />
                <RESULT eventid="1254" status="WDR" swimtime="00:00:00.00" resultid="3047" heatid="7813" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1318" status="WDR" swimtime="00:00:00.00" resultid="3048" heatid="7862" lane="2" entrytime="00:03:20.00" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="3049" heatid="7958" lane="3" entrytime="00:02:42.00" />
                <RESULT eventid="1543" status="WDR" swimtime="00:00:00.00" resultid="3050" entrytime="00:06:45.00" />
                <RESULT eventid="1591" status="WDR" swimtime="00:00:00.00" resultid="3051" heatid="7996" lane="2" entrytime="00:01:25.00" />
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="3052" entrytime="00:05:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-08-24" firstname="Adam" gender="M" lastname="Witkowski" nation="POL" athleteid="3053">
              <RESULTS>
                <RESULT eventid="1156" points="437" swimtime="00:22:10.79" resultid="3054" heatid="8720" lane="2" entrytime="00:22:30.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:18.96" />
                    <SPLIT distance="200" swimtime="00:02:45.19" />
                    <SPLIT distance="300" swimtime="00:04:12.35" />
                    <SPLIT distance="400" swimtime="00:05:42.54" />
                    <SPLIT distance="500" swimtime="00:07:13.29" />
                    <SPLIT distance="600" swimtime="00:08:42.49" />
                    <SPLIT distance="700" swimtime="00:10:11.08" />
                    <SPLIT distance="800" swimtime="00:11:39.85" />
                    <SPLIT distance="900" swimtime="00:13:08.98" />
                    <SPLIT distance="1000" swimtime="00:14:38.51" />
                    <SPLIT distance="1100" swimtime="00:16:08.74" />
                    <SPLIT distance="1200" swimtime="00:17:39.22" />
                    <SPLIT distance="1300" swimtime="00:19:10.45" />
                    <SPLIT distance="1400" swimtime="00:20:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="327" reactiontime="+111" swimtime="00:03:26.69" resultid="3055" heatid="7790" lane="8" entrytime="00:03:25.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:36.72" />
                    <SPLIT distance="150" swimtime="00:02:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="353" reactiontime="+101" swimtime="00:02:37.65" resultid="3056" heatid="7961" lane="1" entrytime="00:02:31.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:13.17" />
                    <SPLIT distance="150" swimtime="00:01:55.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="391" reactiontime="+108" swimtime="00:05:31.42" resultid="3057" heatid="9065" lane="4" entrytime="00:05:32.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:17.16" />
                    <SPLIT distance="150" swimtime="00:01:59.74" />
                    <SPLIT distance="200" swimtime="00:02:42.92" />
                    <SPLIT distance="250" swimtime="00:03:25.95" />
                    <SPLIT distance="300" swimtime="00:04:09.07" />
                    <SPLIT distance="350" swimtime="00:04:51.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-02" firstname="Damian" gender="M" lastname="Jerszyński" nation="POL" athleteid="3058">
              <RESULTS>
                <RESULT eventid="1415" points="435" reactiontime="+79" swimtime="00:00:30.17" resultid="3059" heatid="7918" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1655" points="441" reactiontime="+79" swimtime="00:00:36.53" resultid="3060" heatid="8042" lane="2" entrytime="00:00:36.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-08-14" firstname="Przemysław" gender="M" lastname="Rydlewski" nation="POL" athleteid="3061">
              <RESULTS>
                <RESULT eventid="1108" points="405" reactiontime="+91" swimtime="00:02:39.60" resultid="3062" heatid="7731" lane="7" entrytime="00:02:30.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:11.98" />
                    <SPLIT distance="150" swimtime="00:02:01.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="484" reactiontime="+89" swimtime="00:01:10.05" resultid="3063" heatid="7851" lane="5" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="432" reactiontime="+93" swimtime="00:01:21.11" resultid="3064" heatid="7892" lane="2" entrytime="00:01:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="553" reactiontime="+93" swimtime="00:04:52.68" resultid="3065" heatid="9062" lane="4" entrytime="00:05:01.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                    <SPLIT distance="150" swimtime="00:01:44.24" />
                    <SPLIT distance="200" swimtime="00:02:21.60" />
                    <SPLIT distance="250" swimtime="00:02:59.12" />
                    <SPLIT distance="300" swimtime="00:03:37.41" />
                    <SPLIT distance="350" swimtime="00:04:16.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-26" firstname="Ewa" gender="F" lastname="Jakubowska" nation="POL" athleteid="3066">
              <RESULTS>
                <RESULT eventid="1059" points="288" reactiontime="+101" swimtime="00:00:41.12" resultid="3067" heatid="7674" lane="7" entrytime="00:00:43.20" />
                <RESULT eventid="1206" points="276" reactiontime="+98" swimtime="00:04:14.87" resultid="3068" heatid="7780" lane="2" entrytime="00:03:58.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.64" />
                    <SPLIT distance="100" swimtime="00:01:59.21" />
                    <SPLIT distance="150" swimtime="00:03:08.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="301" reactiontime="+94" swimtime="00:01:52.92" resultid="3069" heatid="7875" lane="2" entrytime="00:01:55.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="312" reactiontime="+103" swimtime="00:00:50.60" resultid="3070" heatid="8023" lane="8" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-12" firstname="Joanna" gender="F" lastname="Chomicz" nation="POL" athleteid="3071">
              <RESULTS>
                <RESULT eventid="1092" points="476" reactiontime="+87" swimtime="00:03:03.35" resultid="3072" heatid="7716" lane="2" entrytime="00:03:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:27.26" />
                    <SPLIT distance="150" swimtime="00:02:20.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="414" swimtime="00:12:26.26" resultid="3073" heatid="8714" lane="4" entrytime="00:13:15.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:01:28.89" />
                    <SPLIT distance="200" swimtime="00:03:00.28" />
                    <SPLIT distance="300" swimtime="00:04:34.28" />
                    <SPLIT distance="400" swimtime="00:06:09.79" />
                    <SPLIT distance="500" swimtime="01:07:46.92" />
                    <SPLIT distance="600" swimtime="00:09:21.50" />
                    <SPLIT distance="700" swimtime="00:10:56.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="452" reactiontime="+82" swimtime="00:01:25.20" resultid="3074" heatid="7833" lane="6" entrytime="00:01:24.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="436" reactiontime="+81" swimtime="00:00:38.33" resultid="3075" heatid="7901" lane="2" entrytime="00:00:38.20" />
                <RESULT eventid="1687" points="455" reactiontime="+82" swimtime="00:05:48.04" resultid="3076" heatid="9050" lane="2" entrytime="00:06:15.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                    <SPLIT distance="100" swimtime="00:01:21.89" />
                    <SPLIT distance="150" swimtime="00:02:05.53" />
                    <SPLIT distance="200" swimtime="00:02:50.22" />
                    <SPLIT distance="250" swimtime="00:03:35.25" />
                    <SPLIT distance="300" swimtime="00:04:21.34" />
                    <SPLIT distance="350" swimtime="00:05:06.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-24" firstname="Aneta" gender="F" lastname="Maduzia" nation="POL" athleteid="3077">
              <RESULTS>
                <RESULT eventid="1140" points="344" swimtime="00:13:13.82" resultid="3078" heatid="8714" lane="5" entrytime="00:13:26.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                    <SPLIT distance="100" swimtime="00:01:30.74" />
                    <SPLIT distance="200" swimtime="00:03:09.01" />
                    <SPLIT distance="300" swimtime="00:04:48.55" />
                    <SPLIT distance="400" swimtime="00:06:30.33" />
                    <SPLIT distance="500" swimtime="00:08:12.23" />
                    <SPLIT distance="600" swimtime="00:09:53.27" />
                    <SPLIT distance="700" swimtime="00:11:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="321" reactiontime="+96" swimtime="00:01:35.46" resultid="3079" heatid="7830" lane="6" entrytime="00:01:34.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="297" reactiontime="+87" swimtime="00:00:43.54" resultid="3080" heatid="7899" lane="2" entrytime="00:00:42.77" />
                <RESULT eventid="1687" points="375" reactiontime="+93" swimtime="00:06:11.23" resultid="3081" heatid="9050" lane="8" entrytime="00:06:21.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:22.83" />
                    <SPLIT distance="150" swimtime="00:02:09.91" />
                    <SPLIT distance="200" swimtime="00:02:57.94" />
                    <SPLIT distance="250" swimtime="00:03:46.71" />
                    <SPLIT distance="300" swimtime="00:04:34.98" />
                    <SPLIT distance="350" swimtime="00:05:23.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="KP Koziegłowy B" number="3">
              <RESULTS>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="3086" heatid="7868" lane="4" entrytime="00:02:33.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3044" number="1" />
                    <RELAYPOSITION athleteid="3053" number="2" />
                    <RELAYPOSITION athleteid="3058" number="3" />
                    <RELAYPOSITION athleteid="3061" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="3087" heatid="7971" lane="5" entrytime="00:02:04.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3044" number="1" />
                    <RELAYPOSITION athleteid="3053" number="2" />
                    <RELAYPOSITION athleteid="3058" number="3" />
                    <RELAYPOSITION athleteid="3061" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="KP Koziegłowy B" number="4">
              <RESULTS>
                <RESULT eventid="1334" reactiontime="+85" swimtime="00:02:47.40" resultid="3088" heatid="7867" lane="1" entrytime="00:02:35.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:30.88" />
                    <SPLIT distance="150" swimtime="00:02:14.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3035" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="3066" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3077" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3071" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1495" reactiontime="+88" swimtime="00:02:26.18" resultid="3089" heatid="7969" lane="8" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:53.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3035" number="1" />
                    <RELAYPOSITION athleteid="3077" number="2" />
                    <RELAYPOSITION athleteid="3066" number="3" />
                    <RELAYPOSITION athleteid="3071" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="KP Koziegłowy C" number="1">
              <RESULTS>
                <RESULT eventid="1671" status="WDR" swimtime="00:00:00.00" resultid="3082" heatid="8050" lane="4" entrytime="00:02:28.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3035" number="1" />
                    <RELAYPOSITION athleteid="3044" number="2" />
                    <RELAYPOSITION athleteid="3071" number="3" />
                    <RELAYPOSITION athleteid="3061" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1124" status="WDR" swimtime="00:00:00.00" resultid="3083" entrytime="00:02:08.44">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3044" number="1" />
                    <RELAYPOSITION athleteid="3035" number="2" />
                    <RELAYPOSITION athleteid="3071" number="3" />
                    <RELAYPOSITION athleteid="3061" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="KP Koziegłowy B" number="2">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+81" swimtime="00:02:03.14" resultid="3084" heatid="7735" lane="2" entrytime="00:02:20.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="150" swimtime="00:01:35.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3071" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3058" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="3035" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3061" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" reactiontime="+86" swimtime="00:02:18.03" resultid="3085" heatid="8050" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:15.51" />
                    <SPLIT distance="150" swimtime="00:01:45.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3035" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="3058" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3061" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="3071" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAKRO" nation="POL" region="08" clubid="5692" name="KP Masters Krosno" shortname="Masters Krosno">
          <CONTACT city="Krosno" email="maciejkoza@op.pl" internet="www.masters.krosoft.pl" name="Maciej Koza" phone="134201024" state="PDK" street="Żwirki i Wigury" street2="4B/19" zip="38-400" />
          <ATHLETES>
            <ATHLETE birthdate="1974-09-09" firstname="Maciej" gender="M" lastname="Koza" nation="POL" athleteid="5693">
              <RESULTS>
                <RESULT eventid="1254" points="260" reactiontime="+105" swimtime="00:01:20.53" resultid="5694" heatid="7809" lane="1" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="186" reactiontime="+108" swimtime="00:03:41.56" resultid="5695" heatid="7860" lane="3" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.33" />
                    <SPLIT distance="100" swimtime="00:01:41.63" />
                    <SPLIT distance="150" swimtime="00:02:41.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="263" reactiontime="+95" swimtime="00:00:40.04" resultid="5696" heatid="7910" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1479" points="223" reactiontime="+130" swimtime="00:03:03.56" resultid="5697" heatid="7953" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:15.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-19" firstname="Artur" gender="M" lastname="Kuryło" nation="POL" athleteid="5698">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5699" heatid="7695" lane="1" entrytime="00:00:31.25" />
                <RESULT eventid="1190" points="340" reactiontime="+85" swimtime="00:00:38.88" resultid="5700" heatid="7762" lane="4" />
                <RESULT eventid="1254" points="316" reactiontime="+87" swimtime="00:01:16.42" resultid="5701" heatid="7811" lane="2" entrytime="00:01:13.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="305" reactiontime="+90" swimtime="00:00:37.30" resultid="5702" heatid="7911" lane="5" entrytime="00:00:36.90" />
                <RESULT eventid="1479" points="268" reactiontime="+91" swimtime="00:02:55.16" resultid="5703" heatid="7954" lane="4" entrytime="00:03:09.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:24.61" />
                    <SPLIT distance="150" swimtime="00:02:12.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-10" firstname="Bogdan" gender="M" lastname="Żebracki" nation="POL" athleteid="5704">
              <RESULTS>
                <RESULT eventid="1076" points="539" reactiontime="+88" swimtime="00:00:29.71" resultid="5705" heatid="7699" lane="3" entrytime="00:00:29.60" />
                <RESULT eventid="1108" points="511" reactiontime="+98" swimtime="00:02:50.82" resultid="5706" heatid="7726" lane="3" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:22.73" />
                    <SPLIT distance="150" swimtime="00:02:12.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="536" reactiontime="+101" swimtime="00:00:35.28" resultid="5707" heatid="7773" lane="7" entrytime="00:00:34.19" />
                <RESULT eventid="1286" points="521" reactiontime="+99" swimtime="00:01:15.13" resultid="5708" heatid="7848" lane="4" entrytime="00:01:14.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="513" reactiontime="+93" swimtime="00:01:23.93" resultid="5709" heatid="7891" lane="2" entrytime="00:01:23.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="472" reactiontime="+92" swimtime="00:01:19.82" resultid="5710" heatid="7938" lane="6" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="544" reactiontime="+90" swimtime="00:00:37.58" resultid="5711" heatid="8040" lane="3" entrytime="00:00:37.10" />
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="5712" entrytime="00:05:40.52" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-08" firstname="Ryszard" gender="M" lastname="Majsiak" nation="POL" athleteid="5713">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)  (Czas: 12:00)" eventid="1254" reactiontime="+71" status="DSQ" swimtime="00:01:24.50" resultid="5714" heatid="7808" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="228" reactiontime="+90" swimtime="00:00:43.25" resultid="5715" heatid="7907" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1479" points="152" reactiontime="+109" swimtime="00:03:34.80" resultid="5716" heatid="7954" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                    <SPLIT distance="100" swimtime="00:01:38.74" />
                    <SPLIT distance="150" swimtime="00:02:37.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Masters Krosno C" number="1">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+87" swimtime="00:02:35.50" resultid="5717" heatid="7868" lane="5" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:24.35" />
                    <SPLIT distance="150" swimtime="00:02:03.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5704" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="5713" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="5693" number="3" reactiontime="+85" />
                    <RELAYPOSITION athleteid="5698" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" reactiontime="+94" swimtime="00:02:12.08" resultid="5718" heatid="7971" lane="2" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:05.42" />
                    <SPLIT distance="150" swimtime="00:01:39.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5704" number="1" />
                    <RELAYPOSITION athleteid="5713" number="2" />
                    <RELAYPOSITION athleteid="5693" number="3" />
                    <RELAYPOSITION athleteid="5698" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02203" nation="POL" region="03" clubid="2292" name="KS AZS AWF Biała Podl." shortname="AZS AWF Biała Podl.">
          <CONTACT city="Biała Podlaska" email="zielakko@gmail.com" name="KS AZS AWF Biała Podlaska" phone="781529483" state="LUBEL" street="Akademicka 2" zip="21-500" />
          <ATHLETES>
            <ATHLETE birthdate="1989-04-27" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" license="102203200002" athleteid="2293">
              <RESULTS>
                <RESULT eventid="1076" points="642" reactiontime="+74" swimtime="00:00:26.65" resultid="2294" heatid="7707" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1108" points="708" reactiontime="+76" swimtime="00:02:22.44" resultid="2295" heatid="7730" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="100" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:47.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEGDY" nation="POL" region="10" clubid="7642" name="KS Delfin Gdynia" shortname="Delfin Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Jakub" gender="M" lastname="Mańczak" nation="POL" athleteid="6298">
              <RESULTS>
                <RESULT eventid="1318" points="477" reactiontime="+73" swimtime="00:02:41.23" resultid="6299" heatid="7864" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:13.28" />
                    <SPLIT distance="150" swimtime="00:01:58.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="655" reactiontime="+75" swimtime="00:00:28.93" resultid="6300" heatid="7921" lane="2" entrytime="00:00:29.40" />
                <RESULT eventid="1479" points="530" reactiontime="+77" swimtime="00:02:19.67" resultid="6301" heatid="7963" lane="1" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:07.77" />
                    <SPLIT distance="150" swimtime="00:01:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="608" reactiontime="+71" swimtime="00:01:06.80" resultid="6302" heatid="8001" lane="8" entrytime="00:01:08.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04211" nation="POL" region="11" clubid="3147" name="KS Delfin Gliwice" shortname="Delfin Gliwice">
          <CONTACT city="Gliwice" email="ksdelfin@op,pl" name="Cupiał" phone="605065587" state="ŚLĄSK" street="Stwosza 8/3" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1944-11-23" firstname="Jerzy" gender="M" lastname="Marciniszko" nation="POL" athleteid="3148">
              <RESULTS>
                <RESULT eventid="1076" points="99" reactiontime="+98" swimtime="00:01:00.75" resultid="3149" heatid="7685" lane="8" entrytime="00:00:56.28" />
                <RESULT eventid="1190" points="102" reactiontime="+104" swimtime="00:01:11.20" resultid="3150" heatid="7763" lane="3" entrytime="00:01:08.01" />
                <RESULT eventid="1222" points="178" reactiontime="+91" swimtime="00:05:23.53" resultid="3151" heatid="7785" lane="1" entrytime="00:05:25.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.19" />
                    <SPLIT distance="100" swimtime="00:02:33.74" />
                    <SPLIT distance="150" swimtime="00:04:00.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="165" reactiontime="+87" swimtime="00:02:24.66" resultid="3152" heatid="7881" lane="3" entrytime="00:02:27.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="83" reactiontime="+114" swimtime="00:02:45.79" resultid="3153" heatid="7932" lane="4" entrytime="00:02:47.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="87" reactiontime="+108" swimtime="00:05:54.60" resultid="3154" heatid="8010" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.09" />
                    <SPLIT distance="100" swimtime="00:02:53.57" />
                    <SPLIT distance="150" swimtime="00:04:26.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="197" reactiontime="+86" swimtime="00:01:00.67" resultid="3155" heatid="8030" lane="3" entrytime="00:00:59.08" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Teodozja" gender="F" lastname="Gdula" nation="POL" athleteid="3156">
              <RESULTS>
                <RESULT eventid="1238" points="125" reactiontime="+85" swimtime="00:02:22.71" resultid="3157" heatid="7797" lane="8" entrytime="00:02:23.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="239" reactiontime="+103" swimtime="00:02:19.20" resultid="3158" heatid="7874" lane="5" entrytime="00:02:14.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="233" reactiontime="+151" swimtime="00:01:02.72" resultid="3159" heatid="8021" lane="6" entrytime="00:01:00.86" />
                <RESULT eventid="1206" points="258" reactiontime="+97" swimtime="00:04:54.37" resultid="5078" heatid="7779" lane="1" entrytime="00:04:44.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.25" />
                    <SPLIT distance="100" swimtime="00:02:23.08" />
                    <SPLIT distance="150" swimtime="00:03:40.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-10" firstname="Barbara" gender="F" lastname="Lipowska" nation="POL" athleteid="3160">
              <RESULTS>
                <RESULT eventid="1206" points="198" reactiontime="+101" swimtime="00:05:04.38" resultid="3161" heatid="7778" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.17" />
                    <SPLIT distance="100" swimtime="00:02:20.75" />
                    <SPLIT distance="150" swimtime="00:03:43.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="118" reactiontime="+94" swimtime="00:02:06.09" resultid="3162" heatid="7796" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" region="DOL" clubid="3298" name="KS Masters Polkowice" shortname="Masters Polkowice">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="ul.Kolejowa 6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1947-04-23" firstname="Bogdan" gender="M" lastname="Jawor" nation="POL" athleteid="3299">
              <RESULTS>
                <RESULT eventid="1076" points="288" reactiontime="+92" swimtime="00:00:42.61" resultid="3300" heatid="7685" lane="5" entrytime="00:00:43.00" entrycourse="SCM" />
                <RESULT eventid="1108" points="252" reactiontime="+93" swimtime="00:04:15.76" resultid="3301" heatid="7720" lane="5" entrytime="00:04:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.70" />
                    <SPLIT distance="100" swimtime="00:02:03.96" />
                    <SPLIT distance="150" swimtime="00:03:15.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="312" reactiontime="+93" swimtime="00:04:28.38" resultid="3302" heatid="7785" lane="4" entrytime="00:04:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.54" />
                    <SPLIT distance="100" swimtime="00:02:09.66" />
                    <SPLIT distance="150" swimtime="00:03:20.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="250" reactiontime="+84" swimtime="00:01:57.19" resultid="3303" heatid="7839" lane="3" entrytime="00:01:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="268" reactiontime="+96" swimtime="00:02:03.08" resultid="3304" heatid="7882" lane="3" entrytime="00:01:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="260" reactiontime="+108" swimtime="00:09:36.67" resultid="3305" heatid="8812" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.69" />
                    <SPLIT distance="100" swimtime="00:02:21.49" />
                    <SPLIT distance="150" swimtime="00:03:37.11" />
                    <SPLIT distance="200" swimtime="00:04:52.25" />
                    <SPLIT distance="250" swimtime="00:06:10.81" />
                    <SPLIT distance="300" swimtime="00:07:28.95" />
                    <SPLIT distance="350" swimtime="00:08:33.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="190" reactiontime="+80" swimtime="00:04:34.18" resultid="3306" heatid="8011" lane="8" entrytime="00:04:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.71" />
                    <SPLIT distance="100" swimtime="00:02:15.48" />
                    <SPLIT distance="150" swimtime="00:03:27.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="290" reactiontime="+91" swimtime="00:00:53.35" resultid="3307" heatid="8031" lane="2" entrytime="00:00:53.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00914" nation="POL" region="14" clubid="2659" name="KS Polonia Warszawa" shortname="Polonia Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1930-01-01" firstname="Lucjan" gender="M" lastname="Prządo" nation="POL" athleteid="2658">
              <RESULTS>
                <RESULT eventid="1076" points="526" reactiontime="+115" swimtime="00:00:41.15" resultid="2660" heatid="7684" lane="2" />
                <RESULT eventid="1190" points="575" reactiontime="+82" swimtime="00:00:52.55" resultid="2661" heatid="7762" lane="5" />
                <RESULT eventid="1222" points="637" reactiontime="+110" swimtime="00:04:16.46" resultid="2662" heatid="7786" lane="8" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.90" />
                    <SPLIT distance="100" swimtime="00:02:00.90" />
                    <SPLIT distance="150" swimtime="00:03:07.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="537" reactiontime="+114" swimtime="00:01:53.49" resultid="2663" heatid="7840" lane="7" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="627" reactiontime="+113" swimtime="00:01:53.22" resultid="2664" heatid="7882" lane="5" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="419" reactiontime="+88" swimtime="00:02:08.44" resultid="2665" heatid="7932" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="754" reactiontime="+107" swimtime="00:00:49.40" resultid="2666" heatid="8031" lane="7" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="3208" name="KS Warta Poznań" shortname="Warta Poznań">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Thiem Jacek" phone="502 499 565" state="WIE" street="Os. Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" athleteid="3209">
              <RESULTS>
                <RESULT eventid="1156" points="378" swimtime="00:24:36.85" resultid="3210" heatid="8722" lane="4" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:01:26.24" />
                    <SPLIT distance="200" swimtime="00:03:01.85" />
                    <SPLIT distance="300" swimtime="00:04:39.98" />
                    <SPLIT distance="400" swimtime="00:06:18.39" />
                    <SPLIT distance="500" swimtime="00:07:57.71" />
                    <SPLIT distance="600" swimtime="00:09:37.22" />
                    <SPLIT distance="700" swimtime="00:11:16.28" />
                    <SPLIT distance="800" swimtime="00:12:56.16" />
                    <SPLIT distance="900" swimtime="00:14:37.49" />
                    <SPLIT distance="1000" swimtime="00:16:18.48" />
                    <SPLIT distance="1100" swimtime="00:18:00.63" />
                    <SPLIT distance="1200" swimtime="00:19:41.33" />
                    <SPLIT distance="1300" swimtime="00:21:22.33" />
                    <SPLIT distance="1400" swimtime="00:23:02.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="433" reactiontime="+104" swimtime="00:03:09.33" resultid="3211" heatid="7862" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                    <SPLIT distance="100" swimtime="00:01:27.68" />
                    <SPLIT distance="150" swimtime="00:02:16.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="380" reactiontime="+109" swimtime="00:02:53.49" resultid="3212" heatid="7958" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="100" swimtime="00:01:25.08" />
                    <SPLIT distance="150" swimtime="00:02:09.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="435" reactiontime="+102" swimtime="00:01:22.43" resultid="3213" heatid="7997" lane="7" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="352" reactiontime="+90" swimtime="00:03:25.30" resultid="3214" heatid="8013" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.98" />
                    <SPLIT distance="100" swimtime="00:01:44.85" />
                    <SPLIT distance="150" swimtime="00:02:36.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" athleteid="3215">
              <RESULTS>
                <RESULT eventid="1140" points="426" swimtime="00:12:44.71" resultid="3216" heatid="8713" lane="6" entrytime="00:12:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:25.73" />
                    <SPLIT distance="200" swimtime="00:02:58.69" />
                    <SPLIT distance="300" swimtime="00:04:33.84" />
                    <SPLIT distance="400" swimtime="00:06:10.79" />
                    <SPLIT distance="500" swimtime="00:07:51.17" />
                    <SPLIT distance="600" swimtime="00:09:29.50" />
                    <SPLIT distance="700" swimtime="00:11:08.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="370" reactiontime="+88" swimtime="00:00:45.37" resultid="3217" heatid="7756" lane="8" entrytime="00:00:46.00" />
                <RESULT eventid="1238" points="404" swimtime="00:01:21.68" resultid="3218" heatid="7801" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="451" reactiontime="+72" swimtime="00:01:32.47" resultid="3219" heatid="7928" lane="1" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="476" swimtime="00:02:51.20" resultid="3220" heatid="7948" lane="6" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="150" swimtime="00:02:06.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="481" reactiontime="+94" swimtime="00:03:16.17" resultid="3221" heatid="8006" lane="5" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:35.09" />
                    <SPLIT distance="150" swimtime="00:02:26.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="426" swimtime="00:06:16.95" resultid="3222" heatid="9050" lane="6" entrytime="00:06:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:25.66" />
                    <SPLIT distance="150" swimtime="00:02:11.86" />
                    <SPLIT distance="200" swimtime="00:03:00.86" />
                    <SPLIT distance="250" swimtime="00:03:50.50" />
                    <SPLIT distance="300" swimtime="00:04:40.18" />
                    <SPLIT distance="350" swimtime="00:05:29.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" athleteid="3223">
              <RESULTS>
                <RESULT eventid="1108" points="542" reactiontime="+86" swimtime="00:02:55.22" resultid="3224" heatid="7725" lane="5" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:14.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="573" reactiontime="+87" swimtime="00:03:06.20" resultid="3225" heatid="7792" lane="4" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:27.27" />
                    <SPLIT distance="150" swimtime="00:02:16.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="540" reactiontime="+90" swimtime="00:01:20.42" resultid="3226" heatid="7845" lane="1" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="552" reactiontime="+104" swimtime="00:01:24.74" resultid="3227" heatid="7890" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="460" reactiontime="+73" swimtime="00:01:23.97" resultid="3228" heatid="7936" lane="4" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="603" reactiontime="+89" swimtime="00:00:37.13" resultid="3229" heatid="8038" lane="2" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" athleteid="3230">
              <RESULTS>
                <RESULT eventid="1156" points="449" swimtime="00:21:30.98" resultid="3231" heatid="8719" lane="1" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="200" swimtime="00:02:34.43" />
                    <SPLIT distance="300" swimtime="00:03:57.13" />
                    <SPLIT distance="400" swimtime="00:05:21.14" />
                    <SPLIT distance="500" swimtime="00:06:47.07" />
                    <SPLIT distance="600" swimtime="00:08:13.17" />
                    <SPLIT distance="700" swimtime="00:09:40.77" />
                    <SPLIT distance="800" swimtime="00:11:11.09" />
                    <SPLIT distance="900" swimtime="00:12:39.46" />
                    <SPLIT distance="1000" swimtime="00:14:08.38" />
                    <SPLIT distance="1100" swimtime="00:15:39.16" />
                    <SPLIT distance="1200" swimtime="00:17:08.78" />
                    <SPLIT distance="1300" swimtime="00:18:38.73" />
                    <SPLIT distance="1400" swimtime="00:20:07.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="646" reactiontime="+80" swimtime="00:00:33.14" resultid="3232" heatid="7772" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1254" points="560" reactiontime="+87" swimtime="00:01:04.17" resultid="3233" heatid="7818" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="603" reactiontime="+82" swimtime="00:01:13.57" resultid="3234" heatid="7940" lane="8" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="577" reactiontime="+80" swimtime="00:02:43.70" resultid="3235" heatid="8016" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                    <SPLIT distance="100" swimtime="00:01:18.56" />
                    <SPLIT distance="150" swimtime="00:02:01.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="Tomaszewski" nation="POL" athleteid="3236">
              <RESULTS>
                <RESULT eventid="1076" points="548" reactiontime="+84" swimtime="00:00:27.04" resultid="3237" heatid="7704" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1190" points="681" reactiontime="+73" swimtime="00:00:30.11" resultid="3238" heatid="7775" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1447" points="620" reactiontime="+77" swimtime="00:01:07.48" resultid="3239" heatid="7940" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-05-14" firstname="Przemysław" gender="M" lastname="Isalski" nation="POL" athleteid="3240">
              <RESULTS>
                <RESULT eventid="1156" points="761" reactiontime="+80" swimtime="00:18:23.98" resultid="3241" heatid="8717" lane="3" entrytime="00:18:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:08.30" />
                    <SPLIT distance="150" swimtime="00:01:45.11" />
                    <SPLIT distance="200" swimtime="00:02:21.58" />
                    <SPLIT distance="250" swimtime="00:02:58.25" />
                    <SPLIT distance="300" swimtime="00:03:35.03" />
                    <SPLIT distance="350" swimtime="00:04:11.90" />
                    <SPLIT distance="400" swimtime="00:04:48.75" />
                    <SPLIT distance="450" swimtime="00:05:25.87" />
                    <SPLIT distance="500" swimtime="00:06:02.80" />
                    <SPLIT distance="550" swimtime="00:06:39.79" />
                    <SPLIT distance="600" swimtime="00:07:17.06" />
                    <SPLIT distance="650" swimtime="00:07:54.64" />
                    <SPLIT distance="700" swimtime="00:08:32.46" />
                    <SPLIT distance="750" swimtime="00:09:10.17" />
                    <SPLIT distance="800" swimtime="00:09:47.67" />
                    <SPLIT distance="850" swimtime="00:10:25.36" />
                    <SPLIT distance="900" swimtime="00:11:02.64" />
                    <SPLIT distance="950" swimtime="00:11:40.01" />
                    <SPLIT distance="1000" swimtime="00:12:17.68" />
                    <SPLIT distance="1050" swimtime="00:12:55.19" />
                    <SPLIT distance="1100" swimtime="00:13:32.24" />
                    <SPLIT distance="1150" swimtime="00:14:09.30" />
                    <SPLIT distance="1200" swimtime="00:14:46.38" />
                    <SPLIT distance="1250" swimtime="00:15:23.12" />
                    <SPLIT distance="1300" swimtime="00:15:59.37" />
                    <SPLIT distance="1350" swimtime="00:16:35.79" />
                    <SPLIT distance="1400" swimtime="00:17:12.58" />
                    <SPLIT distance="1450" swimtime="00:17:48.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="556" reactiontime="+80" swimtime="00:02:09.50" resultid="3242" heatid="7967" lane="7" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="100" swimtime="00:01:02.36" />
                    <SPLIT distance="150" swimtime="00:01:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="645" reactiontime="+82" swimtime="00:04:38.05" resultid="3243" heatid="9059" lane="2" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                    <SPLIT distance="100" swimtime="00:01:05.57" />
                    <SPLIT distance="150" swimtime="00:01:40.64" />
                    <SPLIT distance="200" swimtime="00:02:16.12" />
                    <SPLIT distance="250" swimtime="00:02:51.49" />
                    <SPLIT distance="300" swimtime="00:03:26.96" />
                    <SPLIT distance="350" swimtime="00:04:02.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-19" firstname="Jakub" gender="M" lastname="Stanoch" nation="POL" athleteid="3244">
              <RESULTS>
                <RESULT eventid="1076" points="559" reactiontime="+66" swimtime="00:00:26.85" resultid="3245" heatid="7710" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1318" points="541" reactiontime="+66" swimtime="00:02:32.17" resultid="3246" heatid="7865" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="512" reactiontime="+65" swimtime="00:00:28.58" resultid="3247" heatid="7924" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1591" points="530" reactiontime="+65" swimtime="00:01:05.00" resultid="3248" heatid="8002" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-20" firstname="Rafał" gender="M" lastname="Liszewski" nation="POL" athleteid="3249">
              <RESULTS>
                <RESULT eventid="1076" points="612" reactiontime="+79" swimtime="00:00:26.90" resultid="3250" heatid="7712" lane="8" entrytime="00:00:25.00" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="3251" heatid="7854" lane="3" entrytime="00:01:07.00" />
                <RESULT eventid="1655" points="633" reactiontime="+73" swimtime="00:00:32.91" resultid="3252" heatid="8045" lane="1" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-02" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" athleteid="3253">
              <RESULTS>
                <RESULT eventid="1076" points="828" reactiontime="+74" swimtime="00:00:27.05" resultid="3254" heatid="7704" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1254" points="878" reactiontime="+73" swimtime="00:00:58.92" resultid="3255" heatid="7821" lane="3" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="870" reactiontime="+78" swimtime="00:02:11.74" resultid="3256" heatid="7965" lane="2" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                    <SPLIT distance="100" swimtime="00:01:04.22" />
                    <SPLIT distance="150" swimtime="00:01:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="809" reactiontime="+75" swimtime="00:04:45.89" resultid="3257" heatid="9060" lane="8" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:45.70" />
                    <SPLIT distance="200" swimtime="00:02:23.29" />
                    <SPLIT distance="250" swimtime="00:03:01.07" />
                    <SPLIT distance="300" swimtime="00:03:38.19" />
                    <SPLIT distance="350" swimtime="00:04:13.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-11-17" firstname="Zbigniew" gender="M" lastname="Liber" nation="POL" athleteid="3258">
              <RESULTS>
                <RESULT eventid="1076" points="195" reactiontime="+119" swimtime="00:00:43.75" resultid="3259" heatid="7685" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1222" points="171" reactiontime="+130" swimtime="00:04:38.50" resultid="3260" heatid="7785" lane="3" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.22" />
                    <SPLIT distance="100" swimtime="00:02:15.58" />
                    <SPLIT distance="150" swimtime="00:03:28.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="168" reactiontime="+109" swimtime="00:02:06.04" resultid="3261" heatid="7881" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="166" reactiontime="+116" swimtime="00:00:57.01" resultid="3262" heatid="8030" lane="7" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-09" firstname="Adrian" gender="M" lastname="Sobkowiak" nation="POL" athleteid="3263">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3264" heatid="7694" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="3265" heatid="7844" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="3266" heatid="7887" lane="8" entrytime="00:01:34.00" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="3267" heatid="7909" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="3268" heatid="8035" lane="2" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-13" firstname="Paweł" gender="M" lastname="Konowalski" nation="POL" athleteid="6260">
              <RESULTS>
                <RESULT eventid="1076" points="529" reactiontime="+68" swimtime="00:00:27.36" resultid="6261" heatid="7705" lane="3" entrytime="00:00:27.60" />
                <RESULT eventid="1254" points="527" reactiontime="+72" swimtime="00:01:00.71" resultid="6262" heatid="7819" lane="6" entrytime="00:01:02.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="6263" heatid="7917" lane="2" entrytime="00:00:31.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Warta Poznań B">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+92" swimtime="00:01:55.59" resultid="3269" heatid="7872" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="150" swimtime="00:01:29.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3236" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="3249" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="3244" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3240" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Warta Poznań C">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+76" swimtime="00:02:10.59" resultid="3271" heatid="7869" lane="2" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:43.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3230" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3223" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="6260" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3253" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" reactiontime="+97" swimtime="00:01:55.60" resultid="3272" heatid="7971" lane="8" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="100" swimtime="00:01:01.24" />
                    <SPLIT distance="150" swimtime="00:01:28.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3223" number="1" />
                    <RELAYPOSITION athleteid="3230" number="2" />
                    <RELAYPOSITION athleteid="6260" number="3" />
                    <RELAYPOSITION athleteid="3253" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Warta Poznań B" number="3">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+74" swimtime="00:01:45.71" resultid="3270" heatid="7974" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.32" />
                    <SPLIT distance="100" swimtime="00:00:52.73" />
                    <SPLIT distance="150" swimtime="00:01:19.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3236" number="1" />
                    <RELAYPOSITION athleteid="3249" number="2" />
                    <RELAYPOSITION athleteid="3244" number="3" />
                    <RELAYPOSITION athleteid="3240" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="5133" name="KU AZS UAM Poznań" shortname="AZS UAM Poznań">
          <CONTACT city="Poznań" email="bartekz009@wp.pl" name="Ziemniarski Bartosz" phone="691679381" state="WLKP" street="Bukowska 96/1" zip="60-396" />
          <ATHLETES>
            <ATHLETE birthdate="1986-09-22" firstname="Bartosz" gender="M" lastname="Ziemniarski" nation="POL" license="S03315200001" athleteid="5134">
              <RESULTS>
                <RESULT eventid="1076" points="838" reactiontime="+70" swimtime="00:00:24.22" resultid="5135" heatid="7712" lane="3" entrytime="00:00:24.39" entrycourse="SCM" />
                <RESULT eventid="1254" points="725" reactiontime="+70" swimtime="00:00:54.06" resultid="5136" heatid="7825" lane="2" entrytime="00:00:54.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="681" reactiontime="+70" swimtime="00:00:26.93" resultid="5137" heatid="7924" lane="2" entrytime="00:00:27.39" entrycourse="SCM" />
                <RESULT eventid="1479" points="839" reactiontime="+71" swimtime="00:01:59.31" resultid="5138" heatid="7966" lane="3" entrytime="00:02:09.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                    <SPLIT distance="100" swimtime="00:00:57.47" />
                    <SPLIT distance="150" swimtime="00:01:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="736" reactiontime="+71" swimtime="00:00:59.71" resultid="5139" heatid="8002" lane="8" entrytime="00:01:03.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="Sterczyński" nation="POL" license="S03315200002" athleteid="5140">
              <RESULTS>
                <RESULT eventid="1108" points="642" reactiontime="+65" swimtime="00:02:19.74" resultid="5141" heatid="7733" lane="2" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:04.94" />
                    <SPLIT distance="150" swimtime="00:01:45.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="686" reactiontime="+65" swimtime="00:01:02.56" resultid="5142" heatid="7856" lane="5" entrytime="00:01:00.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="638" reactiontime="+69" swimtime="00:01:03.91" resultid="5143" heatid="7942" lane="3" entrytime="00:01:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-14" firstname="Jarek" gender="M" lastname="Bystry" nation="POL" athleteid="5144">
              <RESULTS>
                <RESULT eventid="1076" points="567" reactiontime="+71" swimtime="00:00:28.65" resultid="5145" heatid="7701" lane="2" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1479" points="452" reactiontime="+78" swimtime="00:02:25.21" resultid="5146" heatid="7961" lane="7" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:09.23" />
                    <SPLIT distance="150" swimtime="00:01:47.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="412" reactiontime="+84" swimtime="00:05:25.44" resultid="5147" heatid="9065" lane="3" entrytime="00:05:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:17.12" />
                    <SPLIT distance="150" swimtime="00:01:58.67" />
                    <SPLIT distance="200" swimtime="00:02:40.67" />
                    <SPLIT distance="250" swimtime="00:03:22.74" />
                    <SPLIT distance="300" swimtime="00:04:05.17" />
                    <SPLIT distance="350" swimtime="00:04:47.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="Stadnik" nation="POL" license="S03315100003" athleteid="5148">
              <RESULTS>
                <RESULT eventid="1059" points="811" reactiontime="+80" swimtime="00:00:28.39" resultid="5149" heatid="7683" lane="2" entrytime="00:00:28.50" entrycourse="SCM" />
                <RESULT eventid="1173" points="706" reactiontime="+88" swimtime="00:00:34.02" resultid="5150" heatid="7761" lane="8" entrytime="00:00:34.50" entrycourse="SCM" />
                <RESULT eventid="1238" points="813" reactiontime="+82" swimtime="00:01:01.98" resultid="5151" heatid="7805" lane="3" entrytime="00:01:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="689" reactiontime="+82" swimtime="00:02:19.43" resultid="5152" heatid="7951" lane="6" entrytime="00:02:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:06.14" />
                    <SPLIT distance="150" swimtime="00:01:43.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AUJKR" nation="POL" region="06" clubid="6259" name="KU AZS UJ Kraków">
          <ATHLETES>
            <ATHLETE birthdate="1993-05-16" firstname="Joanna" gender="F" lastname="Jasińska" nation="POL" athleteid="1966">
              <RESULTS>
                <RESULT eventid="1059" points="797" reactiontime="+73" swimtime="00:00:28.55" resultid="1967" heatid="7683" lane="5" entrytime="00:00:28.17" />
                <RESULT eventid="1092" points="699" reactiontime="+81" swimtime="00:02:41.10" resultid="1968" heatid="7717" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                    <SPLIT distance="150" swimtime="00:02:01.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="739" reactiontime="+76" swimtime="00:01:03.99" resultid="1969" heatid="7805" lane="1" entrytime="00:01:03.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="722" reactiontime="+74" swimtime="00:01:12.57" resultid="1970" heatid="7837" lane="2" entrytime="00:01:12.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="781" reactiontime="+77" swimtime="00:00:31.08" resultid="1971" heatid="7905" lane="6" entrytime="00:00:31.52" />
                <RESULT eventid="1463" points="576" reactiontime="+82" swimtime="00:02:28.02" resultid="1972" heatid="7950" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:11.03" />
                    <SPLIT distance="150" swimtime="00:01:49.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="578" reactiontime="+70" swimtime="00:02:52.66" resultid="1973" heatid="8009" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                    <SPLIT distance="100" swimtime="00:01:21.35" />
                    <SPLIT distance="150" swimtime="00:02:07.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="599" reactiontime="+79" swimtime="00:00:38.94" resultid="1974" heatid="8027" lane="6" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZWRO" nation="POL" region="01" clubid="3027" name="KU AZS Uniwersytet Wrocławski" shortname="AZS Uniw. Wrocławski">
          <CONTACT name="Wawrzyńczak" />
          <ATHLETES>
            <ATHLETE birthdate="1990-09-11" firstname="Karolina" gender="F" lastname="Wawrzyńczak" nation="POL" athleteid="3028">
              <RESULTS>
                <RESULT eventid="1173" points="647" reactiontime="+73" swimtime="00:00:35.02" resultid="3029" heatid="7761" lane="7" entrytime="00:00:34.40" />
                <RESULT eventid="1270" points="564" reactiontime="+88" swimtime="00:01:18.77" resultid="3030" heatid="7836" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="598" reactiontime="+87" swimtime="00:00:33.98" resultid="3031" heatid="7903" lane="5" entrytime="00:00:34.30" />
                <RESULT eventid="1431" points="655" reactiontime="+66" swimtime="00:01:15.05" resultid="3032" heatid="7931" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="579" reactiontime="+89" swimtime="00:01:16.18" resultid="3033" heatid="7991" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKMOS" nation="RUS" clubid="2718" name="MKMP Moscow">
          <ATHLETES>
            <ATHLETE birthdate="1924-01-01" firstname="Vladimir" gender="M" lastname="Rabinovich" nation="RUS" athleteid="2719">
              <RESULTS>
                <RESULT eventid="1076" points="259" reactiontime="+132" swimtime="00:01:00.85" resultid="2720" heatid="7684" lane="5" entrytime="00:00:58.50" />
                <RESULT eventid="1190" points="308" reactiontime="+73" swimtime="00:01:09.83" resultid="2721" heatid="7763" lane="2" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-01-01" firstname="Alexander" gender="M" lastname="Morshin" nation="RUS" athleteid="2722">
              <RESULTS>
                <RESULT eventid="1190" points="454" reactiontime="+85" swimtime="00:00:43.33" resultid="2723" heatid="7767" lane="6" entrytime="00:00:44.30" />
                <RESULT eventid="1383" points="602" reactiontime="+101" swimtime="00:01:34.00" resultid="2724" heatid="7886" lane="3" entrytime="00:01:34.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="647" reactiontime="+98" swimtime="00:00:40.84" resultid="2725" heatid="8035" lane="8" entrytime="00:00:42.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00116" nation="POL" region="16" clubid="3102" name="MKP Szczecin">
          <CONTACT city="Szczecin" email="windmuhle@wp.pl" name="Kowalczyk Piotr" phone="509758055" state="ZACH" street="Kaliny 45/9" zip="71-118" />
          <ATHLETES>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="3103">
              <RESULTS>
                <RESULT eventid="1140" points="705" reactiontime="+82" swimtime="00:10:46.78" resultid="3104" heatid="8712" lane="3" entrytime="00:10:24.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:51.14" />
                    <SPLIT distance="200" swimtime="00:02:30.97" />
                    <SPLIT distance="250" swimtime="00:03:11.44" />
                    <SPLIT distance="300" swimtime="00:03:52.44" />
                    <SPLIT distance="350" swimtime="00:04:33.50" />
                    <SPLIT distance="400" swimtime="00:05:14.63" />
                    <SPLIT distance="450" swimtime="00:05:55.95" />
                    <SPLIT distance="500" swimtime="00:06:37.68" />
                    <SPLIT distance="550" swimtime="00:07:19.34" />
                    <SPLIT distance="600" swimtime="00:08:00.86" />
                    <SPLIT distance="650" swimtime="00:08:42.45" />
                    <SPLIT distance="700" swimtime="00:09:24.09" />
                    <SPLIT distance="750" swimtime="00:10:05.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="683" reactiontime="+78" swimtime="00:01:08.58" resultid="3105" heatid="7804" lane="6" entrytime="00:01:06.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="735" reactiontime="+78" swimtime="00:02:28.17" resultid="3106" heatid="7951" lane="7" entrytime="00:02:24.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="150" swimtime="00:01:50.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="680" reactiontime="+86" swimtime="00:02:54.85" resultid="3107" heatid="8009" lane="6" entrytime="00:02:42.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="100" swimtime="00:01:26.72" />
                    <SPLIT distance="150" swimtime="00:02:11.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="698" reactiontime="+79" swimtime="00:05:19.84" resultid="3108" heatid="9047" lane="2" entrytime="00:05:07.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:54.84" />
                    <SPLIT distance="200" swimtime="00:02:35.65" />
                    <SPLIT distance="250" swimtime="00:03:17.03" />
                    <SPLIT distance="300" swimtime="00:03:58.63" />
                    <SPLIT distance="350" swimtime="00:04:40.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="3109">
              <RESULTS>
                <RESULT eventid="1156" points="664" reactiontime="+82" swimtime="00:19:17.71" resultid="3110" heatid="8717" lane="1" entrytime="00:19:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:47.62" />
                    <SPLIT distance="200" swimtime="00:02:25.13" />
                    <SPLIT distance="250" swimtime="00:03:03.07" />
                    <SPLIT distance="300" swimtime="00:03:41.22" />
                    <SPLIT distance="350" swimtime="00:04:19.79" />
                    <SPLIT distance="400" swimtime="00:04:58.99" />
                    <SPLIT distance="450" swimtime="00:05:37.89" />
                    <SPLIT distance="500" swimtime="00:06:16.77" />
                    <SPLIT distance="550" swimtime="00:06:55.86" />
                    <SPLIT distance="600" swimtime="00:07:34.93" />
                    <SPLIT distance="650" swimtime="00:08:14.21" />
                    <SPLIT distance="700" swimtime="00:08:53.06" />
                    <SPLIT distance="750" swimtime="00:09:32.37" />
                    <SPLIT distance="800" swimtime="00:10:11.24" />
                    <SPLIT distance="850" swimtime="00:10:50.32" />
                    <SPLIT distance="900" swimtime="00:11:29.28" />
                    <SPLIT distance="950" swimtime="00:12:08.29" />
                    <SPLIT distance="1000" swimtime="00:12:47.84" />
                    <SPLIT distance="1050" swimtime="00:13:26.96" />
                    <SPLIT distance="1100" swimtime="00:14:06.45" />
                    <SPLIT distance="1150" swimtime="00:14:46.28" />
                    <SPLIT distance="1200" swimtime="00:15:25.44" />
                    <SPLIT distance="1250" swimtime="00:16:04.91" />
                    <SPLIT distance="1300" swimtime="00:16:44.39" />
                    <SPLIT distance="1350" swimtime="00:17:24.19" />
                    <SPLIT distance="1400" swimtime="00:18:02.84" />
                    <SPLIT distance="1450" swimtime="00:18:42.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="618" reactiontime="+72" swimtime="00:01:00.36" resultid="3111" heatid="7820" lane="7" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="585" reactiontime="+77" swimtime="00:02:13.23" resultid="3112" heatid="7965" lane="3" entrytime="00:02:13.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="100" swimtime="00:01:03.79" />
                    <SPLIT distance="150" swimtime="00:01:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="3113" heatid="8018" lane="7" entrytime="00:02:36.00" />
                <RESULT eventid="1703" points="600" reactiontime="+83" swimtime="00:04:47.30" resultid="3114" heatid="9060" lane="3" entrytime="00:04:47.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:45.80" />
                    <SPLIT distance="200" swimtime="00:02:23.22" />
                    <SPLIT distance="250" swimtime="00:02:59.81" />
                    <SPLIT distance="300" swimtime="00:03:36.08" />
                    <SPLIT distance="350" swimtime="00:04:13.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-08-21" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="3115">
              <RESULTS>
                <RESULT eventid="1206" points="640" swimtime="00:04:55.59" resultid="3116" heatid="7779" lane="8" entrytime="00:04:44.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.79" />
                    <SPLIT distance="100" swimtime="00:02:21.51" />
                    <SPLIT distance="150" swimtime="00:03:40.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="553" swimtime="00:02:16.40" resultid="3117" heatid="7874" lane="3" entrytime="00:02:14.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="369" swimtime="00:01:05.72" resultid="3118" heatid="8021" lane="2" entrytime="00:01:04.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-09" firstname="Piotr" gender="M" lastname="Nowicki" nation="POL" athleteid="3119">
              <RESULTS>
                <RESULT eventid="1076" points="252" reactiontime="+98" swimtime="00:00:37.52" resultid="3120" heatid="7687" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1254" points="249" reactiontime="+81" swimtime="00:01:21.71" resultid="3121" heatid="7809" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="227" reactiontime="+95" swimtime="00:03:02.63" resultid="3122" heatid="7956" lane="7" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:26.89" />
                    <SPLIT distance="150" swimtime="00:02:15.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQGUB" nation="POL" region="04" clubid="6166" name="MKS Aquatic Gubin" shortname="Aquatic Gubin">
          <CONTACT city="Gubin" email="mks@gubin.com.pl" name="PatekZiemowit" phone="693323270" state="LUBUS" street="Piastowska 26" zip="66-620" />
          <ATHLETES>
            <ATHLETE birthdate="1953-05-24" firstname="Anna" gender="F" lastname="Krupińska" nation="POL" athleteid="6167">
              <RESULTS>
                <RESULT eventid="1206" points="424" reactiontime="+110" swimtime="00:04:09.32" resultid="6168" heatid="7780" lane="5" entrytime="00:03:54.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.49" />
                    <SPLIT distance="100" swimtime="00:01:58.91" />
                    <SPLIT distance="150" swimtime="00:03:04.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="450" reactiontime="+116" swimtime="00:01:52.72" resultid="6169" heatid="7876" lane="3" entrytime="00:01:47.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" status="DNS" swimtime="00:00:00.00" resultid="6170" heatid="8024" lane="2" entrytime="00:00:48.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="4123" name="MKS Astoria Bydgoszcz" shortname="Astoria Bydgoszcz">
          <CONTACT email="sikoreczka7@o2.pl" name="Sikorska" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Krzysztof" gender="M" lastname="Kawecki" nation="POL" athleteid="4133">
              <RESULTS>
                <RESULT eventid="1108" points="553" reactiontime="+91" swimtime="00:03:00.50" resultid="4134" heatid="7725" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:26.28" />
                    <SPLIT distance="150" swimtime="00:02:17.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="600" reactiontime="+84" swimtime="00:03:12.75" resultid="4135" heatid="7791" lane="1" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                    <SPLIT distance="100" swimtime="00:01:32.35" />
                    <SPLIT distance="150" swimtime="00:02:22.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="4136" heatid="7889" lane="1" entrytime="00:01:28.00" />
                <RESULT eventid="1543" points="549" reactiontime="+90" swimtime="00:06:35.77" resultid="4137" heatid="8809" lane="1" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                    <SPLIT distance="100" swimtime="00:01:36.48" />
                    <SPLIT distance="150" swimtime="00:02:26.69" />
                    <SPLIT distance="200" swimtime="00:03:16.51" />
                    <SPLIT distance="250" swimtime="00:04:12.51" />
                    <SPLIT distance="300" swimtime="00:05:07.44" />
                    <SPLIT distance="350" swimtime="00:05:51.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="4138" heatid="8014" lane="3" entrytime="00:03:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1928-01-01" firstname="Wacława" gender="F" lastname="Wilczyńska" nation="POL" athleteid="4139">
              <RESULTS>
                <RESULT eventid="1173" points="489" reactiontime="+70" swimtime="00:01:29.81" resultid="4140" heatid="7754" lane="8" entrytime="00:01:23.00" />
                <RESULT eventid="1238" points="519" swimtime="00:02:37.89" resultid="4141" heatid="7796" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="241" swimtime="00:04:09.73" resultid="4142" heatid="7873" lane="4" entrytime="00:03:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:57.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="416" swimtime="00:06:05.06" resultid="4143" heatid="7943" lane="4" entrytime="00:05:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.93" />
                    <SPLIT distance="100" swimtime="00:02:54.52" />
                    <SPLIT distance="150" swimtime="00:04:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="478" reactiontime="+82" swimtime="00:07:00.07" resultid="4144" heatid="8004" lane="3" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:38.55" />
                    <SPLIT distance="100" swimtime="00:03:24.43" />
                    <SPLIT distance="150" swimtime="00:05:11.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Małgorzata" gender="F" lastname="Sikorska" nation="POL" athleteid="4145">
              <RESULTS>
                <RESULT eventid="1140" points="499" swimtime="00:12:05.53" resultid="4146" heatid="8716" lane="2" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="200" swimtime="00:02:52.36" />
                    <SPLIT distance="300" swimtime="00:04:22.49" />
                    <SPLIT distance="400" swimtime="00:05:55.23" />
                    <SPLIT distance="500" swimtime="00:07:27.60" />
                    <SPLIT distance="600" swimtime="00:09:00.09" />
                    <SPLIT distance="700" swimtime="00:10:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="4147" heatid="7802" lane="6" entrytime="00:01:15.00" />
                <RESULT eventid="1463" points="567" reactiontime="+93" swimtime="00:02:41.49" resultid="4148" heatid="7948" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                    <SPLIT distance="150" swimtime="00:01:59.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="537" reactiontime="+100" swimtime="00:06:42.90" resultid="4149" heatid="8802" lane="7" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:37.64" />
                    <SPLIT distance="150" swimtime="00:02:27.39" />
                    <SPLIT distance="200" swimtime="00:03:17.48" />
                    <SPLIT distance="250" swimtime="00:04:16.01" />
                    <SPLIT distance="300" swimtime="00:05:14.66" />
                    <SPLIT distance="350" swimtime="00:05:59.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="573" reactiontime="+87" swimtime="00:03:05.02" resultid="4150" heatid="8006" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                    <SPLIT distance="100" swimtime="00:01:30.87" />
                    <SPLIT distance="150" swimtime="00:02:18.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06414" nation="POL" region="14" clubid="3503" name="MKS Piaseczno">
          <CONTACT city="PIASECZNO" name="ANDRZEJ RUBASZKIEWICZ" />
          <ATHLETES>
            <ATHLETE birthdate="1949-04-10" firstname="Andrzej" gender="M" lastname="Rubaszkiewicz" nation="POL" license="106414200002" athleteid="3510">
              <RESULTS>
                <RESULT eventid="1076" points="794" reactiontime="+76" swimtime="00:00:29.15" resultid="3511" heatid="7697" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1190" points="652" reactiontime="+87" swimtime="00:00:38.22" resultid="3512" heatid="7771" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1254" points="752" reactiontime="+78" swimtime="00:01:05.83" resultid="3513" heatid="7815" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="798" reactiontime="+81" swimtime="00:00:32.27" resultid="3514" heatid="7914" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1479" points="665" reactiontime="+83" swimtime="00:02:37.93" resultid="3515" heatid="7960" lane="4" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:57.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOBIA" nation="POL" region="09" clubid="2285" name="MOS Białystok">
          <CONTACT city="Białystok" email="rafalperkowskibr@gmail.com" name="MOS Białystok Rafał Perkowski" phone="792869333" zip="15-795" />
          <ATHLETES>
            <ATHLETE birthdate="1993-06-04" firstname="Rafał" gender="M" lastname="Perkowski" nation="POL" athleteid="2286">
              <RESULTS>
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="2287" heatid="7789" lane="2" entrytime="00:03:30.00" />
                <RESULT eventid="1286" points="503" reactiontime="+70" swimtime="00:01:12.21" resultid="2288" heatid="7850" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="458" reactiontime="+71" swimtime="00:01:20.10" resultid="2289" heatid="7892" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="2290" heatid="7916" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1655" points="506" reactiontime="+60" swimtime="00:00:35.46" resultid="2291" heatid="8044" lane="7" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOCZE" nation="POL" region="11" clubid="2597" name="MOSiR Częstochowa">
          <ATHLETES>
            <ATHLETE birthdate="1969-07-22" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="2596">
              <RESULTS>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="2598" heatid="7956" lane="6" entrytime="00:02:55.00" />
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="2599" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01012" nation="POL" region="12" clubid="2235" name="MOSiR Ostrowiec Św.">
          <CONTACT email="basen@mosir.ostrowiec.pl" name="Różalski" street="Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" license="M01012200001" athleteid="2236">
              <RESULTS>
                <RESULT eventid="1076" points="737" reactiontime="+87" swimtime="00:00:31.18" resultid="2237" heatid="7692" lane="6" entrytime="00:00:32.50" />
                <RESULT eventid="1108" points="575" reactiontime="+96" swimtime="00:03:14.38" resultid="2238" heatid="7722" lane="2" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:01:36.03" />
                    <SPLIT distance="150" swimtime="00:02:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="667" reactiontime="+88" swimtime="00:01:24.58" resultid="2239" heatid="7842" lane="1" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="429" reactiontime="+91" swimtime="00:03:41.91" resultid="2240" heatid="7861" lane="2" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:43.53" />
                    <SPLIT distance="150" swimtime="00:02:44.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="727" reactiontime="+91" swimtime="00:00:33.98" resultid="2241" heatid="7913" lane="4" entrytime="00:00:34.50" />
                <RESULT eventid="1543" points="528" reactiontime="+99" swimtime="00:07:35.37" resultid="2242" heatid="8811" lane="5" entrytime="00:07:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                    <SPLIT distance="100" swimtime="00:01:45.99" />
                    <SPLIT distance="150" swimtime="00:02:48.50" />
                    <SPLIT distance="200" swimtime="00:03:49.52" />
                    <SPLIT distance="250" swimtime="00:04:52.07" />
                    <SPLIT distance="300" swimtime="00:05:56.56" />
                    <SPLIT distance="350" swimtime="00:06:46.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="490" reactiontime="+96" swimtime="00:01:30.82" resultid="2243" heatid="7995" lane="1" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="505" reactiontime="+94" swimtime="00:06:25.43" resultid="2244" heatid="9068" lane="8" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="100" swimtime="00:01:28.07" />
                    <SPLIT distance="150" swimtime="00:02:18.78" />
                    <SPLIT distance="200" swimtime="00:03:10.17" />
                    <SPLIT distance="250" swimtime="00:04:00.66" />
                    <SPLIT distance="300" swimtime="00:04:50.18" />
                    <SPLIT distance="350" swimtime="00:05:40.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MPPR" nation="SVK" region="SSO" clubid="6313" name="MPK Previdza">
          <ATHLETES>
            <ATHLETE birthdate="1949-01-01" firstname="Maria" gender="F" lastname="Hausnerova" nation="POL" athleteid="6312">
              <RESULTS>
                <RESULT eventid="1059" points="662" reactiontime="+77" swimtime="00:00:36.88" resultid="6314" heatid="7676" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1173" points="752" reactiontime="+70" swimtime="00:00:43.64" resultid="6315" heatid="7756" lane="4" entrytime="00:00:43.90" />
                <RESULT eventid="1238" points="628" swimtime="00:01:23.38" resultid="6316" heatid="7800" lane="1" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="689" reactiontime="+73" swimtime="00:01:34.98" resultid="6317" heatid="7927" lane="3" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" status="WDR" swimtime="00:00:00.00" resultid="6318" entrytime="00:07:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Nina" gender="F" lastname="Hlatka" nation="SVK" athleteid="6319">
              <RESULTS>
                <RESULT eventid="1059" points="661" reactiontime="+82" swimtime="00:00:31.87" resultid="6320" heatid="7680" lane="1" entrytime="00:00:33.10" />
                <RESULT eventid="1238" points="631" reactiontime="+85" swimtime="00:01:10.43" resultid="6321" heatid="7803" lane="7" entrytime="00:01:12.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="598" reactiontime="+85" swimtime="00:02:38.67" resultid="6322" heatid="7949" lane="2" entrytime="00:02:41.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:58.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="518" reactiontime="+86" swimtime="00:00:44.10" resultid="6323" heatid="8025" lane="7" entrytime="00:00:45.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-11-02" firstname="Silvia" gender="F" lastname="Huszarova" nation="SVK" license="SVK15947" athleteid="6381">
              <RESULTS>
                <RESULT eventid="1173" points="528" reactiontime="+78" swimtime="00:00:39.13" resultid="6382" heatid="7756" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1238" points="509" reactiontime="+89" swimtime="00:01:14.42" resultid="6383" heatid="7801" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="557" reactiontime="+91" swimtime="00:01:31.99" resultid="6384" heatid="7877" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="484" reactiontime="+76" swimtime="00:01:26.54" resultid="6385" heatid="7927" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01103" nation="POL" region="03" clubid="5494" name="MTP Lublinianka Lublin" shortname="Lublinianka Lublin">
          <ATHLETES>
            <ATHLETE birthdate="1961-12-08" firstname="Piotr" gender="M" lastname="Kasperek" nation="POL" license="000168" athleteid="5495">
              <RESULTS>
                <RESULT eventid="1156" points="679" reactiontime="+95" swimtime="00:20:15.26" resultid="5496" heatid="8717" lane="7" entrytime="00:19:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:14.17" />
                    <SPLIT distance="150" swimtime="00:01:53.65" />
                    <SPLIT distance="200" swimtime="00:02:33.65" />
                    <SPLIT distance="250" swimtime="00:03:14.30" />
                    <SPLIT distance="300" swimtime="00:03:54.51" />
                    <SPLIT distance="350" swimtime="00:04:34.83" />
                    <SPLIT distance="400" swimtime="00:05:15.27" />
                    <SPLIT distance="450" swimtime="00:05:55.87" />
                    <SPLIT distance="500" swimtime="00:06:36.81" />
                    <SPLIT distance="550" swimtime="00:07:17.47" />
                    <SPLIT distance="600" swimtime="00:07:58.37" />
                    <SPLIT distance="650" swimtime="00:08:39.20" />
                    <SPLIT distance="700" swimtime="00:09:20.22" />
                    <SPLIT distance="750" swimtime="00:10:01.24" />
                    <SPLIT distance="800" swimtime="00:10:42.47" />
                    <SPLIT distance="850" swimtime="00:11:23.21" />
                    <SPLIT distance="900" swimtime="00:12:04.39" />
                    <SPLIT distance="950" swimtime="00:12:45.69" />
                    <SPLIT distance="1000" swimtime="00:13:27.30" />
                    <SPLIT distance="1050" swimtime="00:14:08.65" />
                    <SPLIT distance="1100" swimtime="00:14:50.33" />
                    <SPLIT distance="1150" swimtime="00:15:31.71" />
                    <SPLIT distance="1200" swimtime="00:16:13.22" />
                    <SPLIT distance="1250" swimtime="00:16:54.90" />
                    <SPLIT distance="1300" swimtime="00:17:36.28" />
                    <SPLIT distance="1350" swimtime="00:18:17.25" />
                    <SPLIT distance="1400" swimtime="00:18:58.25" />
                    <SPLIT distance="1450" swimtime="00:19:37.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03001" nation="POL" region="01" clubid="1869" name="MUKP Just Swim Jelenia Góra" shortname="Just Swim J. Góra">
          <CONTACT city="Jelenia Góra" email="marcin.binasiewicz@justswim.pl" name="Binasiewicz Marcin" phone="509071929" state="DOL" zip="58-506" />
          <ATHLETES>
            <ATHLETE birthdate="1983-05-01" firstname="Andrzej" gender="M" lastname="Waszkewicz" nation="POL" license="M0300120009" athleteid="1870">
              <RESULTS>
                <RESULT eventid="1076" points="833" reactiontime="+85" swimtime="00:00:23.52" resultid="1871" heatid="7712" lane="4" entrytime="00:00:23.82" />
                <RESULT eventid="1254" points="797" reactiontime="+86" swimtime="00:00:52.88" resultid="1872" heatid="7825" lane="5" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="728" reactiontime="+87" swimtime="00:00:25.42" resultid="1873" heatid="7925" lane="4" entrytime="00:00:25.20" />
                <RESULT eventid="1591" points="745" reactiontime="+89" swimtime="00:00:58.05" resultid="1874" heatid="8003" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00309" nation="POL" region="09" clubid="2270" name="Masters Białystok">
          <CONTACT email="DOMA44@INTERIA.PL" name="MICHALIK DOMINIKA" phone="608642788" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" license="M00309100100" athleteid="2271">
              <RESULTS>
                <RESULT eventid="1140" points="770" reactiontime="+82" swimtime="00:10:30.81" resultid="2272" heatid="8712" lane="2" entrytime="00:10:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:48.83" />
                    <SPLIT distance="200" swimtime="00:02:27.33" />
                    <SPLIT distance="250" swimtime="00:03:06.24" />
                    <SPLIT distance="300" swimtime="00:03:45.53" />
                    <SPLIT distance="350" swimtime="00:04:24.66" />
                    <SPLIT distance="400" swimtime="00:05:04.04" />
                    <SPLIT distance="450" swimtime="00:05:43.86" />
                    <SPLIT distance="500" swimtime="00:06:24.32" />
                    <SPLIT distance="550" swimtime="00:07:04.78" />
                    <SPLIT distance="600" swimtime="00:07:45.62" />
                    <SPLIT distance="650" swimtime="00:08:27.13" />
                    <SPLIT distance="700" swimtime="00:09:08.96" />
                    <SPLIT distance="750" swimtime="00:09:50.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="587" reactiontime="+82" swimtime="00:01:08.61" resultid="2273" heatid="7804" lane="1" entrytime="00:01:07.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="649" reactiontime="+82" swimtime="00:02:25.41" resultid="2274" heatid="7950" lane="4" entrytime="00:02:28.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:10.92" />
                    <SPLIT distance="150" swimtime="00:01:48.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="729" reactiontime="+81" swimtime="00:05:03.84" resultid="2275" heatid="9048" lane="3" entrytime="00:05:15.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                    <SPLIT distance="150" swimtime="00:01:48.39" />
                    <SPLIT distance="200" swimtime="00:02:26.81" />
                    <SPLIT distance="250" swimtime="00:03:05.49" />
                    <SPLIT distance="300" swimtime="00:03:44.95" />
                    <SPLIT distance="350" swimtime="00:04:24.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Bartosz" gender="M" lastname="Bogdanowicz" nation="POL" athleteid="2276">
              <RESULTS>
                <RESULT eventid="1318" points="434" reactiontime="+89" swimtime="00:02:48.03" resultid="2277" heatid="7864" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:02:09.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="2278" heatid="7941" lane="3" entrytime="00:01:08.00" />
                <RESULT eventid="1543" points="548" reactiontime="+86" swimtime="00:05:33.32" resultid="2279" heatid="8806" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:56.93" />
                    <SPLIT distance="200" swimtime="00:02:38.53" />
                    <SPLIT distance="250" swimtime="00:03:26.90" />
                    <SPLIT distance="300" swimtime="00:04:17.44" />
                    <SPLIT distance="350" swimtime="00:04:56.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="429" reactiontime="+85" swimtime="00:02:34.04" resultid="2280" heatid="8019" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MACHE" nation="POL" region="03" clubid="2742" name="Masters Chełm">
          <ATHLETES>
            <ATHLETE birthdate="1941-10-11" firstname="Janusz" gender="M" lastname="Golik" nation="POL" athleteid="2743">
              <RESULTS>
                <RESULT eventid="1222" points="478" reactiontime="+118" swimtime="00:03:56.83" resultid="2744" heatid="7786" lane="4" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.59" />
                    <SPLIT distance="100" swimtime="00:01:56.05" />
                    <SPLIT distance="150" swimtime="00:02:58.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="353" reactiontime="+120" swimtime="00:04:35.92" resultid="2745" heatid="7859" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.76" />
                    <SPLIT distance="100" swimtime="00:02:16.55" />
                    <SPLIT distance="150" swimtime="00:03:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="492" reactiontime="+112" swimtime="00:01:45.98" resultid="2746" heatid="7891" lane="8" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="198" reactiontime="+121" swimtime="00:02:08.71" resultid="2747" heatid="7933" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="388" reactiontime="+105" swimtime="00:01:51.08" resultid="2748" heatid="7993" lane="7" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="547" reactiontime="+102" swimtime="00:00:45.76" resultid="2749" heatid="8034" lane="1" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-26" firstname="Wiesław" gender="M" lastname="Wepa" nation="POL" athleteid="2750">
              <RESULTS>
                <RESULT eventid="1222" points="321" reactiontime="+88" swimtime="00:03:57.45" resultid="2751" heatid="7786" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.99" />
                    <SPLIT distance="100" swimtime="00:01:55.30" />
                    <SPLIT distance="150" swimtime="00:02:59.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="199" reactiontime="+116" swimtime="00:04:12.78" resultid="2752" heatid="7860" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                    <SPLIT distance="100" swimtime="00:01:56.19" />
                    <SPLIT distance="150" swimtime="00:03:03.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="265" reactiontime="+102" swimtime="00:01:46.05" resultid="2753" heatid="7883" lane="4" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="230" reactiontime="+109" swimtime="00:03:37.37" resultid="2754" heatid="7953" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.99" />
                    <SPLIT distance="100" swimtime="00:01:42.00" />
                    <SPLIT distance="150" swimtime="00:02:40.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="183" reactiontime="+93" swimtime="00:01:53.95" resultid="2755" heatid="7992" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="2756" heatid="9069" lane="8" entrytime="00:07:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-15" firstname="Dariusz" gender="M" lastname="Biskup" nation="POL" athleteid="2757">
              <RESULTS>
                <RESULT eventid="1383" points="133" reactiontime="+136" swimtime="00:01:59.92" resultid="2758" heatid="7881" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="145" reactiontime="+133" swimtime="00:00:52.86" resultid="2759" heatid="8029" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-20" firstname="Hanna" gender="F" lastname="Wepa" nation="POL" athleteid="2760">
              <RESULTS>
                <RESULT eventid="1206" points="189" reactiontime="+109" swimtime="00:05:08.80" resultid="2761" heatid="7778" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.48" />
                    <SPLIT distance="100" swimtime="00:02:30.11" />
                    <SPLIT distance="150" swimtime="00:03:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="69" reactiontime="+118" swimtime="00:02:31.04" resultid="2762" heatid="7796" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="165" reactiontime="+117" swimtime="00:02:26.16" resultid="2763" heatid="7873" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="83" reactiontime="+115" swimtime="00:05:09.15" resultid="2764" heatid="7943" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.61" />
                    <SPLIT distance="100" swimtime="00:02:28.58" />
                    <SPLIT distance="150" swimtime="00:03:48.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="160" reactiontime="+114" swimtime="00:01:07.39" resultid="2765" heatid="8020" lane="6" />
                <RESULT eventid="1687" points="86" reactiontime="+116" swimtime="00:10:47.14" resultid="2766" heatid="9053" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.95" />
                    <SPLIT distance="100" swimtime="00:02:31.82" />
                    <SPLIT distance="150" swimtime="00:03:55.10" />
                    <SPLIT distance="200" swimtime="00:05:18.81" />
                    <SPLIT distance="250" swimtime="00:06:40.79" />
                    <SPLIT distance="300" swimtime="00:08:01.80" />
                    <SPLIT distance="350" swimtime="00:09:25.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAGOR" nation="POL" region="04" clubid="5186" name="Masters Gorzów Wlkp.">
          <CONTACT city="Gorzów Wlkp." email="mastersgorzow@onet.eu" name="Wojciechowicz Marek" phone="602891603" state="LUB" street="Ogińskiego 97/7" zip="66-400" />
          <ATHLETES>
            <ATHLETE birthdate="1970-12-12" firstname="Marek" gender="M" lastname="Wojciechowicz" nation="POL" license="MWOJ" athleteid="5187">
              <RESULTS>
                <RESULT eventid="1076" points="649" reactiontime="+82" swimtime="00:00:27.43" resultid="5188" heatid="7706" lane="8" entrytime="00:00:27.50" entrycourse="SCM" />
                <RESULT eventid="1156" points="549" swimtime="00:20:17.32" resultid="5189" heatid="8719" lane="5" entrytime="00:21:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="200" swimtime="00:02:30.75" />
                    <SPLIT distance="300" swimtime="00:03:49.77" />
                    <SPLIT distance="400" swimtime="00:05:09.38" />
                    <SPLIT distance="500" swimtime="00:06:29.92" />
                    <SPLIT distance="600" swimtime="00:07:51.56" />
                    <SPLIT distance="700" swimtime="00:09:14.12" />
                    <SPLIT distance="800" swimtime="00:10:37.54" />
                    <SPLIT distance="900" swimtime="00:12:01.07" />
                    <SPLIT distance="1000" swimtime="00:13:26.39" />
                    <SPLIT distance="1100" swimtime="00:14:50.89" />
                    <SPLIT distance="1200" swimtime="00:16:14.14" />
                    <SPLIT distance="1300" swimtime="00:17:39.27" />
                    <SPLIT distance="1400" swimtime="00:19:00.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="630" reactiontime="+84" swimtime="00:01:00.74" resultid="5190" heatid="7821" lane="1" entrytime="00:01:01.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="523" reactiontime="+90" swimtime="00:00:31.18" resultid="5191" heatid="7918" lane="6" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1479" points="562" reactiontime="+82" swimtime="00:02:16.90" resultid="5192" heatid="7964" lane="1" entrytime="00:02:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:04.89" />
                    <SPLIT distance="150" swimtime="00:01:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="540" reactiontime="+89" swimtime="00:04:55.39" resultid="5193" heatid="9062" lane="7" entrytime="00:05:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                    <SPLIT distance="150" swimtime="00:01:46.94" />
                    <SPLIT distance="200" swimtime="00:02:24.77" />
                    <SPLIT distance="250" swimtime="00:03:03.38" />
                    <SPLIT distance="300" swimtime="00:03:41.34" />
                    <SPLIT distance="350" swimtime="00:04:19.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" license="MLAS" athleteid="5194">
              <RESULTS>
                <RESULT eventid="1076" points="348" reactiontime="+112" swimtime="00:00:37.05" resultid="5195" heatid="7688" lane="1" entrytime="00:00:36.10" entrycourse="SCM" />
                <RESULT eventid="1156" points="364" swimtime="00:27:01.93" resultid="5196" heatid="8723" lane="1" entrytime="00:28:15.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                    <SPLIT distance="100" swimtime="00:01:30.51" />
                    <SPLIT distance="200" swimtime="00:03:15.99" />
                    <SPLIT distance="300" swimtime="00:05:04.73" />
                    <SPLIT distance="400" swimtime="00:06:54.96" />
                    <SPLIT distance="500" swimtime="00:08:43.78" />
                    <SPLIT distance="600" swimtime="00:10:33.57" />
                    <SPLIT distance="700" swimtime="00:12:23.68" />
                    <SPLIT distance="800" swimtime="00:14:13.50" />
                    <SPLIT distance="900" swimtime="00:16:04.47" />
                    <SPLIT distance="1000" swimtime="00:17:53.54" />
                    <SPLIT distance="1100" swimtime="00:19:43.32" />
                    <SPLIT distance="1200" swimtime="00:21:33.51" />
                    <SPLIT distance="1300" swimtime="00:23:24.38" />
                    <SPLIT distance="1400" swimtime="00:25:15.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="339" reactiontime="+116" swimtime="00:01:23.22" resultid="5197" heatid="7808" lane="3" entrytime="00:01:23.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="325" reactiontime="+115" swimtime="00:03:13.92" resultid="5198" heatid="7954" lane="1" entrytime="00:03:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                    <SPLIT distance="100" swimtime="00:01:29.71" />
                    <SPLIT distance="150" swimtime="00:02:22.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="350" reactiontime="+108" swimtime="00:06:49.74" resultid="5199" heatid="9069" lane="3" entrytime="00:06:52.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                    <SPLIT distance="100" swimtime="00:01:30.99" />
                    <SPLIT distance="150" swimtime="00:02:22.88" />
                    <SPLIT distance="200" swimtime="00:03:16.64" />
                    <SPLIT distance="250" swimtime="00:04:10.87" />
                    <SPLIT distance="300" swimtime="00:05:04.82" />
                    <SPLIT distance="350" swimtime="00:05:59.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-20" firstname="Artur" gender="M" lastname="Rutkowski" nation="POL" license="ARUT" athleteid="5200">
              <RESULTS>
                <RESULT eventid="1108" points="469" reactiontime="+83" swimtime="00:02:43.77" resultid="5201" heatid="7729" lane="3" entrytime="00:02:44.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:16.59" />
                    <SPLIT distance="150" swimtime="00:02:05.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="388" reactiontime="+84" swimtime="00:02:53.61" resultid="5202" heatid="7864" lane="8" entrytime="00:02:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:21.10" />
                    <SPLIT distance="150" swimtime="00:02:07.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="557" reactiontime="+77" swimtime="00:00:31.18" resultid="5203" heatid="7918" lane="5" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1543" points="445" reactiontime="+87" swimtime="00:05:57.36" resultid="5204" heatid="8808" lane="5" entrytime="00:06:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="200" swimtime="00:02:52.70" />
                    <SPLIT distance="250" swimtime="00:03:43.88" />
                    <SPLIT distance="300" swimtime="00:04:36.54" />
                    <SPLIT distance="350" swimtime="00:05:17.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="521" reactiontime="+81" swimtime="00:01:10.64" resultid="5205" heatid="7999" lane="3" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-08" firstname="Dawid" gender="M" lastname="Borus" nation="POL" license="DABOR" athleteid="5206">
              <RESULTS>
                <RESULT eventid="1076" points="579" reactiontime="+77" swimtime="00:00:28.50" resultid="5207" heatid="7703" lane="8" entrytime="00:00:28.30" entrycourse="SCM" />
                <RESULT eventid="1108" points="478" reactiontime="+75" swimtime="00:02:43.53" resultid="5208" heatid="7728" lane="5" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:15.25" />
                    <SPLIT distance="150" swimtime="00:02:03.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="572" reactiontime="+68" swimtime="00:00:32.69" resultid="5209" heatid="7774" lane="1" entrytime="00:00:33.30" entrycourse="SCM" />
                <RESULT eventid="1286" points="617" reactiontime="+79" swimtime="00:01:10.25" resultid="5210" heatid="7851" lane="6" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="5211" heatid="7892" lane="4" entrytime="00:01:20.00" entrycourse="SCM" />
                <RESULT eventid="1447" points="596" reactiontime="+66" swimtime="00:01:10.16" resultid="5212" heatid="7940" lane="2" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="582" reactiontime="+66" swimtime="00:02:37.42" resultid="5213" heatid="8016" lane="2" entrytime="00:02:48.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:16.71" />
                    <SPLIT distance="150" swimtime="00:01:57.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="556" reactiontime="+82" swimtime="00:00:35.85" resultid="5214" heatid="8042" lane="5" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-06-11" firstname="Artur" gender="M" lastname="Łopaciński" nation="POL" license="AŁOP" athleteid="5215">
              <RESULTS>
                <RESULT eventid="1108" points="429" reactiontime="+70" swimtime="00:02:49.53" resultid="5216" heatid="7728" lane="3" entrytime="00:02:46.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:18.07" />
                    <SPLIT distance="150" swimtime="00:02:09.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="540" reactiontime="+67" swimtime="00:01:03.94" resultid="5217" heatid="7818" lane="7" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="495" reactiontime="+69" swimtime="00:01:15.61" resultid="5218" heatid="7850" lane="8" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="491" reactiontime="+67" swimtime="00:00:31.85" resultid="5219" heatid="7917" lane="7" entrytime="00:00:31.30" entrycourse="SCM" />
                <RESULT eventid="1543" points="390" reactiontime="+78" swimtime="00:06:10.76" resultid="5220" heatid="8808" lane="3" entrytime="00:06:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:21.98" />
                    <SPLIT distance="150" swimtime="00:02:10.24" />
                    <SPLIT distance="200" swimtime="00:02:58.08" />
                    <SPLIT distance="250" swimtime="00:03:52.99" />
                    <SPLIT distance="300" swimtime="00:04:47.00" />
                    <SPLIT distance="350" swimtime="00:05:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="5221" heatid="7999" lane="7" entrytime="00:01:12.00" entrycourse="SCM" />
                <RESULT eventid="1703" points="402" reactiontime="+78" swimtime="00:05:25.88" resultid="5222" heatid="9064" lane="4" entrytime="00:05:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="150" swimtime="00:01:57.54" />
                    <SPLIT distance="200" swimtime="00:02:39.89" />
                    <SPLIT distance="250" swimtime="00:03:22.08" />
                    <SPLIT distance="300" swimtime="00:04:04.48" />
                    <SPLIT distance="350" swimtime="00:04:46.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Masters Gorzów C" number="1">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+81" swimtime="00:01:54.04" resultid="5223" heatid="7972" lane="5" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                    <SPLIT distance="100" swimtime="00:00:58.19" />
                    <SPLIT distance="150" swimtime="00:01:26.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5206" number="1" />
                    <RELAYPOSITION athleteid="5215" number="2" />
                    <RELAYPOSITION athleteid="5200" number="3" />
                    <RELAYPOSITION athleteid="5187" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1357" reactiontime="+67" swimtime="00:02:10.11" resultid="5224" heatid="7870" lane="4" entrytime="00:02:11.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:09.10" />
                    <SPLIT distance="150" swimtime="00:01:41.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5206" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="5215" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5200" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="5187" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00306" nation="POL" region="06" clubid="3710" name="Masters Korona Kraków">
          <CONTACT city="Kraków" email="masterskorona@wp.pl" internet="www.masterskorona.pl" name="Mariola Kuliś" phone="500677133" state="MAŁ" street="Kalwaryjska" />
          <ATHLETES>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="3711">
              <RESULTS>
                <RESULT eventid="1059" points="718" reactiontime="+74" swimtime="00:00:31.00" resultid="3712" heatid="7681" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1238" points="610" reactiontime="+79" swimtime="00:01:11.21" resultid="3713" heatid="7803" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="700" reactiontime="+76" swimtime="00:00:39.90" resultid="3714" heatid="8023" lane="3" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-27" firstname="Wacław" gender="M" lastname="Brożek" nation="POL" athleteid="3718">
              <RESULTS>
                <RESULT eventid="1108" points="252" reactiontime="+94" swimtime="00:03:36.23" resultid="3719" heatid="7722" lane="3" entrytime="00:03:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.20" />
                    <SPLIT distance="100" swimtime="00:01:43.69" />
                    <SPLIT distance="150" swimtime="00:02:49.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="285" swimtime="00:25:02.08" resultid="3720" heatid="8723" lane="2" entrytime="00:27:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:01:26.98" />
                    <SPLIT distance="200" swimtime="00:03:02.84" />
                    <SPLIT distance="300" swimtime="00:04:43.01" />
                    <SPLIT distance="400" swimtime="00:06:24.65" />
                    <SPLIT distance="500" swimtime="00:08:06.35" />
                    <SPLIT distance="600" swimtime="00:09:48.32" />
                    <SPLIT distance="700" swimtime="00:11:29.48" />
                    <SPLIT distance="800" swimtime="00:13:12.12" />
                    <SPLIT distance="900" swimtime="00:14:54.04" />
                    <SPLIT distance="1000" swimtime="00:16:36.60" />
                    <SPLIT distance="1100" swimtime="00:18:16.85" />
                    <SPLIT distance="1200" swimtime="00:19:58.70" />
                    <SPLIT distance="1300" swimtime="00:21:40.90" />
                    <SPLIT distance="1400" swimtime="00:23:22.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="144" reactiontime="+52" swimtime="00:00:54.66" resultid="3721" heatid="7764" lane="5" entrytime="00:00:54.00" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="3722" heatid="7841" lane="1" entrytime="00:01:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-04-24" firstname="Krzysztof" gender="M" lastname="Chołda" nation="POL" athleteid="3723">
              <RESULTS>
                <RESULT eventid="1156" points="386" swimtime="00:22:36.75" resultid="3724" heatid="8721" lane="6" entrytime="00:23:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                    <SPLIT distance="100" swimtime="00:01:21.92" />
                    <SPLIT distance="200" swimtime="00:02:49.45" />
                    <SPLIT distance="300" swimtime="00:04:18.08" />
                    <SPLIT distance="400" swimtime="00:05:48.47" />
                    <SPLIT distance="500" swimtime="00:07:19.78" />
                    <SPLIT distance="600" swimtime="00:08:51.91" />
                    <SPLIT distance="700" swimtime="00:10:23.72" />
                    <SPLIT distance="800" swimtime="00:11:56.00" />
                    <SPLIT distance="900" swimtime="00:13:28.53" />
                    <SPLIT distance="1000" swimtime="00:15:00.56" />
                    <SPLIT distance="1100" swimtime="00:16:32.55" />
                    <SPLIT distance="1200" swimtime="00:18:04.57" />
                    <SPLIT distance="1300" swimtime="00:19:36.36" />
                    <SPLIT distance="1400" swimtime="00:21:09.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="373" reactiontime="+100" swimtime="00:01:24.02" resultid="3725" heatid="7844" lane="5" entrytime="00:01:24.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="411" reactiontime="+97" swimtime="00:01:30.39" resultid="3726" heatid="7887" lane="7" entrytime="00:01:33.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="394" reactiontime="+95" swimtime="00:05:35.21" resultid="3727" heatid="9065" lane="8" entrytime="00:05:44.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-08-18" firstname="Jadwiga" gender="F" lastname="Gorecka" nation="POL" athleteid="3728">
              <RESULTS>
                <RESULT eventid="1059" points="654" reactiontime="+75" swimtime="00:00:34.85" resultid="3729" heatid="7676" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1238" points="613" reactiontime="+76" swimtime="00:01:20.63" resultid="3730" heatid="7800" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="507" reactiontime="+89" swimtime="00:01:37.15" resultid="3731" heatid="7829" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="566" reactiontime="+79" swimtime="00:00:41.25" resultid="3732" heatid="7899" lane="7" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-09-19" firstname="Maciej" gender="M" lastname="Grudzień" nation="POL" athleteid="3733">
              <RESULTS>
                <RESULT eventid="1076" points="397" reactiontime="+90" swimtime="00:00:31.06" resultid="3734" heatid="7698" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1108" points="278" reactiontime="+90" swimtime="00:03:04.67" resultid="3735" heatid="7726" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:31.01" />
                    <SPLIT distance="150" swimtime="00:02:23.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="286" reactiontime="+93" swimtime="00:00:42.86" resultid="3736" heatid="8035" lane="4" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-13" firstname="Michał" gender="M" lastname="Gugała" nation="POL" athleteid="3737">
              <RESULTS>
                <RESULT eventid="1076" points="407" reactiontime="+104" swimtime="00:00:29.84" resultid="3738" heatid="7696" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="1156" points="395" swimtime="00:22:53.83" resultid="3739" heatid="8720" lane="7" entrytime="00:22:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="200" swimtime="00:02:53.86" />
                    <SPLIT distance="300" swimtime="00:04:26.05" />
                    <SPLIT distance="400" swimtime="00:05:38.15" />
                    <SPLIT distance="500" swimtime="00:07:30.35" />
                    <SPLIT distance="600" swimtime="00:09:03.18" />
                    <SPLIT distance="700" swimtime="00:10:36.43" />
                    <SPLIT distance="800" swimtime="00:12:10.12" />
                    <SPLIT distance="900" swimtime="00:13:43.49" />
                    <SPLIT distance="1000" swimtime="00:15:17.58" />
                    <SPLIT distance="1100" swimtime="00:16:49.23" />
                    <SPLIT distance="1200" swimtime="00:18:21.40" />
                    <SPLIT distance="1300" swimtime="00:19:54.16" />
                    <SPLIT distance="1400" swimtime="00:21:26.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="3740" heatid="7769" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="3741" heatid="7814" lane="3" entrytime="00:01:09.00" />
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="3742" heatid="7936" lane="7" entrytime="00:01:30.00" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="3743" heatid="7955" lane="1" entrytime="00:02:45.00" />
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="3744" heatid="9066" lane="8" entrytime="00:05:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="3745">
              <RESULTS>
                <RESULT eventid="1059" points="494" reactiontime="+91" swimtime="00:00:34.38" resultid="3746" heatid="7679" lane="3" entrytime="00:00:33.90" />
                <RESULT eventid="1173" points="506" reactiontime="+86" swimtime="00:00:39.67" resultid="3747" heatid="7758" lane="2" entrytime="00:00:39.95" />
                <RESULT eventid="1270" points="402" reactiontime="+96" swimtime="00:01:32.31" resultid="3748" heatid="7831" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="520" reactiontime="+90" swimtime="00:00:37.14" resultid="3749" heatid="7901" lane="4" entrytime="00:00:37.70" />
                <RESULT eventid="1431" status="DNS" swimtime="00:00:00.00" resultid="3750" heatid="7928" lane="5" entrytime="00:01:30.00" />
                <RESULT eventid="1607" points="459" reactiontime="+105" swimtime="00:03:13.62" resultid="3751" heatid="8006" lane="6" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                    <SPLIT distance="100" swimtime="00:01:34.48" />
                    <SPLIT distance="150" swimtime="00:02:26.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-26" firstname="Anna" gender="F" lastname="Kasprzykowska" nation="POL" athleteid="3752">
              <RESULTS>
                <RESULT eventid="1059" points="195" reactiontime="+105" swimtime="00:00:45.06" resultid="3753" heatid="7673" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1399" points="150" reactiontime="+101" swimtime="00:00:54.61" resultid="3754" heatid="7898" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1687" points="161" reactiontime="+104" swimtime="00:08:22.05" resultid="3755" heatid="9052" lane="7" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.76" />
                    <SPLIT distance="100" swimtime="00:01:59.02" />
                    <SPLIT distance="150" swimtime="00:03:03.99" />
                    <SPLIT distance="200" swimtime="00:04:09.05" />
                    <SPLIT distance="250" swimtime="00:05:13.39" />
                    <SPLIT distance="300" swimtime="00:06:18.04" />
                    <SPLIT distance="350" swimtime="00:07:23.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-12" firstname="Wojciech" gender="M" lastname="Hoffman" nation="POL" athleteid="3756">
              <RESULTS>
                <RESULT eventid="1156" points="560" swimtime="00:20:25.28" resultid="3757" heatid="8719" lane="3" entrytime="00:21:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:12.95" />
                    <SPLIT distance="200" swimtime="00:02:30.36" />
                    <SPLIT distance="300" swimtime="00:03:49.75" />
                    <SPLIT distance="400" swimtime="00:05:10.45" />
                    <SPLIT distance="500" swimtime="00:06:31.89" />
                    <SPLIT distance="600" swimtime="00:07:54.65" />
                    <SPLIT distance="700" swimtime="00:09:17.47" />
                    <SPLIT distance="800" swimtime="00:10:40.23" />
                    <SPLIT distance="900" swimtime="00:12:01.52" />
                    <SPLIT distance="1000" swimtime="00:13:28.04" />
                    <SPLIT distance="1100" swimtime="00:14:51.69" />
                    <SPLIT distance="1200" swimtime="00:16:41.68" />
                    <SPLIT distance="1300" swimtime="00:17:39.75" />
                    <SPLIT distance="1400" swimtime="00:19:03.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="513" reactiontime="+66" swimtime="00:00:33.89" resultid="3758" heatid="7771" lane="6" entrytime="00:00:35.50" />
                <RESULT eventid="1254" points="503" reactiontime="+76" swimtime="00:01:04.66" resultid="3759" heatid="7818" lane="5" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="486" reactiontime="+64" swimtime="00:01:15.16" resultid="3760" heatid="7935" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="476" reactiontime="+78" swimtime="00:02:22.68" resultid="3761" heatid="7963" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:47.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="499" reactiontime="+83" swimtime="00:05:05.39" resultid="3762" heatid="9070" lane="8" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                    <SPLIT distance="150" swimtime="00:01:51.73" />
                    <SPLIT distance="200" swimtime="00:02:30.06" />
                    <SPLIT distance="250" swimtime="00:03:08.76" />
                    <SPLIT distance="300" swimtime="00:03:47.70" />
                    <SPLIT distance="350" swimtime="00:04:27.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-02" firstname="Wojciech" gender="M" lastname="Kaczmarczyk" nation="POL" athleteid="3763">
              <RESULTS>
                <RESULT eventid="1076" points="103" reactiontime="+145" swimtime="00:00:51.55" resultid="3764" heatid="7686" lane="7" entrytime="00:00:54.00" />
                <RESULT eventid="1383" points="208" reactiontime="+100" swimtime="00:01:53.40" resultid="3765" heatid="7882" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="249" reactiontime="+111" swimtime="00:00:48.75" resultid="3766" heatid="8031" lane="8" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-04" firstname="Andrzej" gender="M" lastname="Data" nation="POL" athleteid="3767">
              <RESULTS>
                <RESULT eventid="1108" points="359" reactiontime="+102" swimtime="00:03:21.03" resultid="3768" heatid="7723" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:01:34.66" />
                    <SPLIT distance="150" swimtime="00:02:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="380" swimtime="00:24:33.84" resultid="3769" heatid="8721" lane="7" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                    <SPLIT distance="100" swimtime="00:01:23.99" />
                    <SPLIT distance="200" swimtime="00:03:00.71" />
                    <SPLIT distance="300" swimtime="00:04:40.51" />
                    <SPLIT distance="400" swimtime="00:06:20.84" />
                    <SPLIT distance="500" swimtime="00:08:01.45" />
                    <SPLIT distance="600" swimtime="00:09:40.96" />
                    <SPLIT distance="700" swimtime="00:11:20.11" />
                    <SPLIT distance="800" swimtime="00:12:59.77" />
                    <SPLIT distance="900" swimtime="00:14:38.98" />
                    <SPLIT distance="1000" swimtime="00:16:19.10" />
                    <SPLIT distance="1100" swimtime="00:17:58.98" />
                    <SPLIT distance="1200" swimtime="00:19:38.55" />
                    <SPLIT distance="1300" swimtime="00:21:18.69" />
                    <SPLIT distance="1400" swimtime="00:22:58.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="374" reactiontime="+113" swimtime="00:03:34.66" resultid="3770" heatid="7790" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                    <SPLIT distance="100" swimtime="00:01:40.21" />
                    <SPLIT distance="150" swimtime="00:02:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="352" reactiontime="+114" swimtime="00:01:32.72" resultid="3771" heatid="7841" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="360" reactiontime="+99" swimtime="00:00:44.09" resultid="3772" heatid="8034" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1703" points="376" reactiontime="+119" swimtime="00:06:08.88" resultid="3773" heatid="9067" lane="7" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                    <SPLIT distance="150" swimtime="00:02:10.09" />
                    <SPLIT distance="200" swimtime="00:02:57.94" />
                    <SPLIT distance="250" swimtime="00:03:46.87" />
                    <SPLIT distance="300" swimtime="00:04:35.27" />
                    <SPLIT distance="350" swimtime="00:05:24.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-08" firstname="Tomasz" gender="M" lastname="Czerniecki" nation="POL" athleteid="3774">
              <RESULTS>
                <RESULT eventid="1076" points="595" reactiontime="+69" swimtime="00:00:26.30" resultid="3775" heatid="7710" lane="7" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-20" firstname="Joanna" gender="F" lastname="Kieszek" nation="POL" athleteid="3776">
              <RESULTS>
                <RESULT eventid="1059" points="718" reactiontime="+66" swimtime="00:00:29.57" resultid="3777" heatid="7682" lane="5" entrytime="00:00:29.60" />
                <RESULT eventid="1238" points="694" reactiontime="+68" swimtime="00:01:05.36" resultid="3778" heatid="7805" lane="8" entrytime="00:01:04.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="585" reactiontime="+66" swimtime="00:01:17.84" resultid="3779" heatid="7835" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="697" reactiontime="+68" swimtime="00:00:32.28" resultid="3780" heatid="7905" lane="8" entrytime="00:00:32.50" />
                <RESULT eventid="1463" points="585" reactiontime="+71" swimtime="00:02:27.25" resultid="3781" heatid="7949" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="150" swimtime="00:01:49.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="464" reactiontime="+67" swimtime="00:00:42.39" resultid="3782" heatid="8027" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1687" points="468" reactiontime="+72" swimtime="00:05:33.06" resultid="3783" heatid="9048" lane="7" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:15.64" />
                    <SPLIT distance="150" swimtime="00:01:56.64" />
                    <SPLIT distance="200" swimtime="00:02:38.54" />
                    <SPLIT distance="250" swimtime="00:03:21.88" />
                    <SPLIT distance="300" swimtime="00:04:05.31" />
                    <SPLIT distance="350" swimtime="00:04:49.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-07-26" firstname="Anna" gender="F" lastname="Koźmin" nation="POL" athleteid="3784">
              <RESULTS>
                <RESULT eventid="1092" points="343" reactiontime="+111" swimtime="00:04:12.13" resultid="3785" heatid="7714" lane="6" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.80" />
                    <SPLIT distance="100" swimtime="00:02:01.45" />
                    <SPLIT distance="150" swimtime="00:03:08.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="358" reactiontime="+109" swimtime="00:04:23.79" resultid="3786" heatid="7779" lane="2" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.50" />
                    <SPLIT distance="100" swimtime="00:02:02.31" />
                    <SPLIT distance="150" swimtime="00:03:14.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="331" reactiontime="+111" swimtime="00:01:54.29" resultid="3787" heatid="7828" lane="1" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="387" reactiontime="+106" swimtime="00:01:58.59" resultid="3788" heatid="7875" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="455" reactiontime="+105" swimtime="00:00:50.16" resultid="3789" heatid="8022" lane="2" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-16" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="3790">
              <RESULTS>
                <RESULT eventid="1076" points="254" reactiontime="+113" swimtime="00:00:45.79" resultid="3791" heatid="7685" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="3792" heatid="7720" lane="1" entrytime="00:05:10.00" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="3793" heatid="7763" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1286" points="142" reactiontime="+111" swimtime="00:02:30.08" resultid="3794" heatid="7839" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="3795" heatid="7933" lane="1" entrytime="00:02:15.00" />
                <RESULT eventid="1479" points="240" reactiontime="+138" swimtime="00:04:02.11" resultid="3796" heatid="7953" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.82" />
                    <SPLIT distance="100" swimtime="00:01:53.04" />
                    <SPLIT distance="150" swimtime="00:02:59.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="195" reactiontime="+115" swimtime="00:09:36.42" resultid="3797" heatid="9070" lane="5" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.92" />
                    <SPLIT distance="100" swimtime="00:01:55.52" />
                    <SPLIT distance="150" swimtime="00:03:17.28" />
                    <SPLIT distance="200" swimtime="00:05:52.77" />
                    <SPLIT distance="250" swimtime="00:07:11.75" />
                    <SPLIT distance="300" swimtime="00:08:31.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-06-03" firstname="Antoni" gender="M" lastname="Kubis" nation="POL" athleteid="3798">
              <RESULTS>
                <RESULT eventid="1076" points="383" reactiontime="+111" swimtime="00:00:38.76" resultid="3799" heatid="7685" lane="7" entrytime="00:00:47.00" />
                <RESULT eventid="1190" points="261" reactiontime="+88" swimtime="00:00:52.13" resultid="3800" heatid="7765" lane="1" entrytime="00:00:52.00" />
                <RESULT eventid="1286" points="346" reactiontime="+119" swimtime="00:01:45.23" resultid="3801" heatid="7840" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="3802" heatid="7907" lane="7" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-12" firstname="Joanna" gender="F" lastname="Kwatera" nation="POL" athleteid="3803">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="3804" heatid="7715" lane="4" entrytime="00:03:12.00" />
                <RESULT eventid="1206" points="485" reactiontime="+76" swimtime="00:03:15.49" resultid="3805" heatid="7783" lane="8" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:32.30" />
                    <SPLIT distance="150" swimtime="00:02:23.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="398" reactiontime="+75" swimtime="00:01:28.91" resultid="3806" heatid="7831" lane="5" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="475" reactiontime="+72" swimtime="00:01:30.50" resultid="3807" heatid="7879" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="397" reactiontime="+77" swimtime="00:06:54.37" resultid="3808" heatid="8804" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                    <SPLIT distance="100" swimtime="00:01:48.38" />
                    <SPLIT distance="150" swimtime="00:02:43.10" />
                    <SPLIT distance="200" swimtime="00:03:36.68" />
                    <SPLIT distance="250" swimtime="00:04:28.13" />
                    <SPLIT distance="300" swimtime="00:05:20.10" />
                    <SPLIT distance="350" swimtime="00:06:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="412" reactiontime="+77" swimtime="00:00:42.43" resultid="3809" heatid="8026" lane="5" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="3810">
              <RESULTS>
                <RESULT eventid="1076" points="619" reactiontime="+128" swimtime="00:00:33.04" resultid="3811" heatid="7693" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1156" points="550" swimtime="00:26:51.57" resultid="3812" heatid="8722" lane="6" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                    <SPLIT distance="100" swimtime="00:01:41.02" />
                    <SPLIT distance="200" swimtime="00:03:32.74" />
                    <SPLIT distance="300" swimtime="00:05:19.98" />
                    <SPLIT distance="400" swimtime="00:07:09.60" />
                    <SPLIT distance="500" swimtime="00:08:58.31" />
                    <SPLIT distance="600" swimtime="00:10:46.25" />
                    <SPLIT distance="700" swimtime="00:12:33.80" />
                    <SPLIT distance="800" swimtime="00:14:27.51" />
                    <SPLIT distance="900" swimtime="00:16:11.42" />
                    <SPLIT distance="1000" swimtime="00:17:59.23" />
                    <SPLIT distance="1100" swimtime="00:00:19.49" />
                    <SPLIT distance="1200" swimtime="00:21:38.00" />
                    <SPLIT distance="1300" swimtime="00:23:25.05" />
                    <SPLIT distance="1400" swimtime="00:25:10.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="650" reactiontime="+132" swimtime="00:01:13.17" resultid="3813" heatid="7812" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="286" reactiontime="+135" swimtime="00:04:13.88" resultid="3814" heatid="7860" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.06" />
                    <SPLIT distance="100" swimtime="00:02:06.34" />
                    <SPLIT distance="150" swimtime="00:03:16.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="580" reactiontime="+122" swimtime="00:02:54.96" resultid="3815" heatid="7957" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="100" swimtime="00:01:21.97" />
                    <SPLIT distance="150" swimtime="00:02:08.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="408" reactiontime="+135" swimtime="00:08:16.34" resultid="3816" heatid="8811" lane="3" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.16" />
                    <SPLIT distance="100" swimtime="00:02:02.17" />
                    <SPLIT distance="150" swimtime="00:04:17.74" />
                    <SPLIT distance="200" swimtime="00:05:25.08" />
                    <SPLIT distance="250" swimtime="00:06:32.33" />
                    <SPLIT distance="350" swimtime="00:07:28.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="287" reactiontime="+122" swimtime="00:01:48.51" resultid="3817" heatid="7994" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="444" reactiontime="+135" swimtime="00:06:42.48" resultid="3818" heatid="9067" lane="8" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:30.31" />
                    <SPLIT distance="150" swimtime="00:02:21.09" />
                    <SPLIT distance="200" swimtime="00:03:12.64" />
                    <SPLIT distance="250" swimtime="00:04:05.85" />
                    <SPLIT distance="300" swimtime="00:04:58.97" />
                    <SPLIT distance="350" swimtime="00:05:52.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="3819">
              <RESULTS>
                <RESULT eventid="1059" points="160" reactiontime="+114" swimtime="00:00:59.29" resultid="3820" heatid="7672" lane="8" entrytime="00:00:56.00" />
                <RESULT eventid="1092" points="158" reactiontime="+107" swimtime="00:05:37.55" resultid="3821" heatid="7713" lane="4" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.54" />
                    <SPLIT distance="100" swimtime="00:02:55.29" />
                    <SPLIT distance="150" swimtime="00:04:25.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="173" reactiontime="+115" swimtime="00:02:07.13" resultid="3822" heatid="7797" lane="7" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="161" reactiontime="+109" swimtime="00:02:30.27" resultid="3823" heatid="7827" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="122" reactiontime="+119" swimtime="00:01:14.35" resultid="3824" heatid="7897" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1463" points="212" reactiontime="+117" swimtime="00:04:34.82" resultid="3825" heatid="7944" lane="7" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.83" />
                    <SPLIT distance="100" swimtime="00:02:10.55" />
                    <SPLIT distance="150" swimtime="00:03:21.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="274" reactiontime="+118" swimtime="00:01:03.43" resultid="3826" heatid="8021" lane="5" entrytime="00:00:59.00" />
                <RESULT eventid="1687" points="210" reactiontime="+111" swimtime="00:09:52.59" resultid="3827" heatid="9053" lane="4" entrytime="00:10:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.54" />
                    <SPLIT distance="100" swimtime="00:02:09.26" />
                    <SPLIT distance="150" swimtime="00:03:23.19" />
                    <SPLIT distance="200" swimtime="00:04:38.48" />
                    <SPLIT distance="250" swimtime="00:05:51.87" />
                    <SPLIT distance="300" swimtime="00:07:07.04" />
                    <SPLIT distance="350" swimtime="00:08:29.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="3828">
              <RESULTS>
                <RESULT eventid="1076" points="658" reactiontime="+89" swimtime="00:00:29.21" resultid="3829" heatid="7700" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="1190" points="560" reactiontime="+87" swimtime="00:00:35.63" resultid="3830" heatid="7772" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1286" points="658" reactiontime="+94" swimtime="00:01:15.28" resultid="3831" heatid="7847" lane="2" entrytime="00:01:16.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="712" reactiontime="+93" swimtime="00:00:30.85" resultid="3832" heatid="7915" lane="5" entrytime="00:00:32.80" />
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="3833" heatid="7938" lane="4" entrytime="00:01:17.30" />
                <RESULT eventid="1591" points="631" reactiontime="+105" swimtime="00:01:12.81" resultid="3834" heatid="7998" lane="2" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="586" reactiontime="+93" swimtime="00:00:37.49" resultid="3835" heatid="8042" lane="1" entrytime="00:00:36.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-16" firstname="Kamil" gender="M" lastname="Latuszek" nation="POL" athleteid="3836">
              <RESULTS>
                <RESULT eventid="1076" points="714" reactiontime="+74" swimtime="00:00:25.55" resultid="3837" heatid="7709" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="1254" points="622" reactiontime="+73" swimtime="00:00:56.89" resultid="3838" heatid="7823" lane="7" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="612" reactiontime="+78" swimtime="00:02:12.50" resultid="3839" heatid="7964" lane="5" entrytime="00:02:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="100" swimtime="00:01:03.75" />
                    <SPLIT distance="150" swimtime="00:01:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="593" reactiontime="+76" swimtime="00:04:50.96" resultid="3840" heatid="9061" lane="1" entrytime="00:05:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:07.41" />
                    <SPLIT distance="150" swimtime="00:01:44.27" />
                    <SPLIT distance="200" swimtime="00:02:21.33" />
                    <SPLIT distance="250" swimtime="00:02:58.55" />
                    <SPLIT distance="300" swimtime="00:03:36.02" />
                    <SPLIT distance="350" swimtime="00:04:14.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="Palmowska" nation="POL" athleteid="3841">
              <RESULTS>
                <RESULT eventid="1092" points="641" reactiontime="+69" swimtime="00:02:45.97" resultid="3842" heatid="7717" lane="2" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:14.28" />
                    <SPLIT distance="150" swimtime="00:02:04.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="728" reactiontime="+65" swimtime="00:00:34.31" resultid="3843" heatid="7760" lane="4" entrytime="00:00:34.50" />
                <RESULT eventid="1270" points="658" reactiontime="+66" swimtime="00:01:15.21" resultid="3844" heatid="7836" lane="2" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="630" reactiontime="+65" swimtime="00:01:14.35" resultid="3845" heatid="7931" lane="8" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="539" reactiontime="+68" swimtime="00:06:14.03" resultid="3846" heatid="8804" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:22.60" />
                    <SPLIT distance="150" swimtime="00:02:12.55" />
                    <SPLIT distance="200" swimtime="00:03:01.15" />
                    <SPLIT distance="250" swimtime="00:03:52.80" />
                    <SPLIT distance="300" swimtime="00:04:45.33" />
                    <SPLIT distance="350" swimtime="00:05:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="602" reactiontime="+61" swimtime="00:02:41.53" resultid="3847" heatid="8009" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:17.58" />
                    <SPLIT distance="150" swimtime="00:02:00.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="534" reactiontime="+67" swimtime="00:05:30.00" resultid="3848" heatid="9049" lane="6" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="150" swimtime="00:02:01.00" />
                    <SPLIT distance="200" swimtime="00:02:44.29" />
                    <SPLIT distance="250" swimtime="00:03:26.95" />
                    <SPLIT distance="300" swimtime="00:04:09.71" />
                    <SPLIT distance="350" swimtime="00:04:51.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-18" firstname="Bartosz" gender="M" lastname="Próchniewicz" nation="POL" athleteid="3849">
              <RESULTS>
                <RESULT eventid="1076" points="178" reactiontime="+81" swimtime="00:00:42.15" resultid="3850" heatid="7685" lane="6" entrytime="00:00:46.00" />
                <RESULT eventid="1190" points="175" reactiontime="+71" swimtime="00:00:48.52" resultid="3851" heatid="7764" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1447" points="157" reactiontime="+67" swimtime="00:01:49.48" resultid="3852" heatid="7934" lane="1" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-12-18" firstname="Szymon" gender="M" lastname="Pyrć" nation="POL" athleteid="3853">
              <RESULTS>
                <RESULT eventid="1156" points="626" swimtime="00:19:25.10" resultid="3854" heatid="8718" lane="5" entrytime="00:20:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="200" swimtime="00:02:30.89" />
                    <SPLIT distance="300" swimtime="00:03:48.70" />
                    <SPLIT distance="400" swimtime="00:05:06.17" />
                    <SPLIT distance="500" swimtime="00:06:23.97" />
                    <SPLIT distance="600" swimtime="00:07:42.00" />
                    <SPLIT distance="700" swimtime="00:09:00.19" />
                    <SPLIT distance="800" swimtime="00:10:18.32" />
                    <SPLIT distance="900" swimtime="00:11:36.27" />
                    <SPLIT distance="1000" swimtime="00:12:53.71" />
                    <SPLIT distance="1100" swimtime="00:14:11.74" />
                    <SPLIT distance="1200" swimtime="00:15:30.83" />
                    <SPLIT distance="1300" swimtime="00:16:49.19" />
                    <SPLIT distance="1400" swimtime="00:18:08.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="615" reactiontime="+79" swimtime="00:02:28.22" resultid="3855" heatid="7865" lane="1" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                    <SPLIT distance="150" swimtime="00:01:50.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="555" reactiontime="+84" swimtime="00:05:29.84" resultid="3856" heatid="8807" lane="5" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                    <SPLIT distance="150" swimtime="00:01:57.04" />
                    <SPLIT distance="200" swimtime="00:02:40.64" />
                    <SPLIT distance="250" swimtime="00:03:29.12" />
                    <SPLIT distance="300" swimtime="00:04:16.86" />
                    <SPLIT distance="350" swimtime="00:04:54.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="582" reactiontime="+79" swimtime="00:01:07.80" resultid="3857" heatid="8001" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-22" firstname="Alicja" gender="F" lastname="Romańska" nation="POL" athleteid="3858">
              <RESULTS>
                <RESULT eventid="1140" points="280" swimtime="00:14:24.68" resultid="3859" heatid="8715" lane="5" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.04" />
                    <SPLIT distance="100" swimtime="00:01:52.93" />
                    <SPLIT distance="200" swimtime="00:03:41.06" />
                    <SPLIT distance="300" swimtime="00:05:28.01" />
                    <SPLIT distance="400" swimtime="00:07:17.76" />
                    <SPLIT distance="500" swimtime="00:09:06.86" />
                    <SPLIT distance="600" swimtime="00:10:54.00" />
                    <SPLIT distance="700" swimtime="00:12:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="215" reactiontime="+106" swimtime="00:01:36.46" resultid="3860" heatid="7797" lane="4" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="249" reactiontime="+125" swimtime="00:03:23.52" resultid="3861" heatid="7946" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:40.82" />
                    <SPLIT distance="150" swimtime="00:02:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-08-09" firstname="Michał" gender="M" lastname="Binkowski" nation="POL" athleteid="3862">
              <RESULTS>
                <RESULT eventid="1076" points="586" reactiontime="+83" swimtime="00:00:26.44" resultid="3863" heatid="7710" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1254" points="544" reactiontime="+78" swimtime="00:01:00.06" resultid="3864" heatid="7821" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-12-07" firstname="Robert" gender="M" lastname="Kominiak" nation="POL" athleteid="3865">
              <RESULTS>
                <RESULT eventid="1076" points="594" reactiontime="+78" swimtime="00:00:28.75" resultid="3866" heatid="7706" lane="5" entrytime="00:00:27.20" />
                <RESULT eventid="1286" points="561" reactiontime="+80" swimtime="00:01:13.31" resultid="3867" heatid="7848" lane="8" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="633" reactiontime="+84" swimtime="00:01:18.25" resultid="3868" heatid="7893" lane="5" entrytime="00:01:16.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="589" reactiontime="+72" swimtime="00:00:31.53" resultid="3869" heatid="7921" lane="6" entrytime="00:00:29.10" />
                <RESULT eventid="1655" points="727" reactiontime="+75" swimtime="00:00:34.11" resultid="3870" heatid="8044" lane="2" entrytime="00:00:34.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="3871">
              <RESULTS>
                <RESULT eventid="1173" points="199" reactiontime="+72" swimtime="00:00:54.10" resultid="3872" heatid="7754" lane="3" entrytime="00:00:56.00" />
                <RESULT eventid="1206" points="231" reactiontime="+127" swimtime="00:04:30.55" resultid="3873" heatid="7779" lane="7" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.54" />
                    <SPLIT distance="100" swimtime="00:02:09.99" />
                    <SPLIT distance="150" swimtime="00:03:21.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="211" reactiontime="+124" swimtime="00:02:06.94" resultid="3874" heatid="7874" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" status="DNS" swimtime="00:00:00.00" resultid="3875" heatid="7926" lane="5" entrytime="00:02:10.00" />
                <RESULT eventid="1607" points="177" reactiontime="+76" swimtime="00:04:25.63" resultid="3876" heatid="8005" lane="1" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.85" />
                    <SPLIT distance="100" swimtime="00:02:06.86" />
                    <SPLIT distance="150" swimtime="00:03:19.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="180" reactiontime="+123" swimtime="00:01:00.72" resultid="3877" heatid="8021" lane="3" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="3878">
              <RESULTS>
                <RESULT eventid="1092" points="607" reactiontime="+86" swimtime="00:03:00.65" resultid="3879" heatid="7716" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:24.14" />
                    <SPLIT distance="150" swimtime="00:02:18.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="628" reactiontime="+83" swimtime="00:01:22.37" resultid="3880" heatid="7834" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="592" reactiontime="+91" swimtime="00:00:35.74" resultid="3881" heatid="7904" lane="8" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="Wysocka" nation="POL" athleteid="3882">
              <RESULTS>
                <RESULT eventid="1059" points="534" reactiontime="+88" swimtime="00:00:35.12" resultid="3883" heatid="7677" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1206" points="737" reactiontime="+95" swimtime="00:03:16.49" resultid="3884" heatid="7782" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.55" />
                    <SPLIT distance="100" swimtime="00:01:32.78" />
                    <SPLIT distance="150" swimtime="00:02:24.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="681" reactiontime="+94" swimtime="00:01:31.16" resultid="3885" heatid="7879" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="637" reactiontime="+93" swimtime="00:00:42.59" resultid="3886" heatid="8026" lane="3" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="Frączek" nation="POL" athleteid="3887">
              <RESULTS>
                <RESULT eventid="1059" points="726" reactiontime="+81" swimtime="00:00:30.24" resultid="3888" heatid="7682" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1173" points="623" reactiontime="+64" swimtime="00:00:37.03" resultid="3889" heatid="7759" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1270" points="603" reactiontime="+77" swimtime="00:01:20.62" resultid="3890" heatid="7834" lane="4" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="654" reactiontime="+76" swimtime="00:00:34.40" resultid="3891" heatid="7903" lane="2" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="3892">
              <RESULTS>
                <RESULT eventid="1156" points="395" swimtime="00:31:27.23" resultid="3893" heatid="8724" lane="8" entrytime="00:38:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.51" />
                    <SPLIT distance="100" swimtime="00:01:51.94" />
                    <SPLIT distance="200" swimtime="00:03:59.18" />
                    <SPLIT distance="300" swimtime="00:06:08.85" />
                    <SPLIT distance="400" swimtime="00:08:17.45" />
                    <SPLIT distance="500" swimtime="00:10:25.20" />
                    <SPLIT distance="600" swimtime="00:12:32.55" />
                    <SPLIT distance="700" swimtime="00:14:40.45" />
                    <SPLIT distance="800" swimtime="00:16:47.09" />
                    <SPLIT distance="900" swimtime="00:18:54.37" />
                    <SPLIT distance="1000" swimtime="00:21:01.30" />
                    <SPLIT distance="1100" swimtime="00:23:07.11" />
                    <SPLIT distance="1200" swimtime="00:25:13.14" />
                    <SPLIT distance="1300" swimtime="00:27:19.18" />
                    <SPLIT distance="1400" swimtime="00:29:24.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-04-07" firstname="Jacek" gender="M" lastname="Żurek" nation="POL" athleteid="3894">
              <RESULTS>
                <RESULT eventid="1076" points="573" reactiontime="+87" swimtime="00:00:27.49" resultid="3895" heatid="7709" lane="7" entrytime="00:00:26.50" />
                <RESULT eventid="1156" points="528" swimtime="00:19:58.00" resultid="3896" heatid="8718" lane="4" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:09.84" />
                    <SPLIT distance="200" swimtime="00:02:25.29" />
                    <SPLIT distance="300" swimtime="00:03:44.31" />
                    <SPLIT distance="400" swimtime="00:05:04.44" />
                    <SPLIT distance="500" swimtime="00:06:24.65" />
                    <SPLIT distance="600" swimtime="00:07:46.08" />
                    <SPLIT distance="700" swimtime="00:09:07.97" />
                    <SPLIT distance="800" swimtime="00:10:29.60" />
                    <SPLIT distance="900" swimtime="00:11:50.53" />
                    <SPLIT distance="1000" swimtime="00:13:12.09" />
                    <SPLIT distance="1100" swimtime="00:14:33.18" />
                    <SPLIT distance="1200" swimtime="00:15:54.64" />
                    <SPLIT distance="1300" swimtime="00:17:15.88" />
                    <SPLIT distance="1400" swimtime="00:18:37.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="492" reactiontime="+72" swimtime="00:01:01.50" resultid="3897" heatid="7823" lane="1" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="427" reactiontime="+78" swimtime="00:00:31.47" resultid="3898" heatid="7918" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1479" points="551" reactiontime="+78" swimtime="00:02:17.28" resultid="3899" heatid="7964" lane="7" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:04.70" />
                    <SPLIT distance="150" swimtime="00:01:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="566" reactiontime="+76" swimtime="00:04:55.39" resultid="3900" heatid="9060" lane="2" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:07.05" />
                    <SPLIT distance="150" swimtime="00:01:43.83" />
                    <SPLIT distance="200" swimtime="00:02:21.49" />
                    <SPLIT distance="250" swimtime="00:03:00.22" />
                    <SPLIT distance="300" swimtime="00:03:38.87" />
                    <SPLIT distance="350" swimtime="00:04:18.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-17" firstname="Kinga" gender="F" lastname="Sowa" nation="POL" athleteid="3901">
              <RESULTS>
                <RESULT eventid="1059" points="718" reactiontime="+83" swimtime="00:00:29.56" resultid="3902" heatid="7682" lane="6" entrytime="00:00:29.96" />
                <RESULT eventid="1173" points="703" reactiontime="+69" swimtime="00:00:34.07" resultid="3903" heatid="7760" lane="3" entrytime="00:00:34.77" />
                <RESULT eventid="1238" points="586" reactiontime="+96" swimtime="00:01:09.14" resultid="3904" heatid="7804" lane="8" entrytime="00:01:08.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="721" reactiontime="+73" swimtime="00:01:12.68" resultid="3905" heatid="7931" lane="1" entrytime="00:01:15.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-01" firstname="Karolina" gender="F" lastname="Zadrożna" nation="POL" athleteid="3906">
              <RESULTS>
                <RESULT eventid="1140" points="682" reactiontime="+86" swimtime="00:10:22.38" resultid="3907" heatid="8712" lane="6" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:12.97" />
                    <SPLIT distance="150" swimtime="00:01:51.43" />
                    <SPLIT distance="200" swimtime="00:02:30.35" />
                    <SPLIT distance="250" swimtime="00:03:09.27" />
                    <SPLIT distance="300" swimtime="00:03:48.60" />
                    <SPLIT distance="350" swimtime="00:04:27.98" />
                    <SPLIT distance="400" swimtime="00:05:07.47" />
                    <SPLIT distance="450" swimtime="00:05:46.58" />
                    <SPLIT distance="500" swimtime="00:06:26.35" />
                    <SPLIT distance="550" swimtime="00:07:06.25" />
                    <SPLIT distance="600" swimtime="00:07:45.87" />
                    <SPLIT distance="650" swimtime="00:08:25.65" />
                    <SPLIT distance="700" swimtime="00:09:05.22" />
                    <SPLIT distance="750" swimtime="00:09:44.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="669" reactiontime="+81" swimtime="00:01:06.15" resultid="3908" heatid="7804" lane="3" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="265" reactiontime="+85" swimtime="00:03:30.70" resultid="3909" heatid="7858" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:33.60" />
                    <SPLIT distance="150" swimtime="00:02:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="662" reactiontime="+81" swimtime="00:02:21.29" resultid="3910" heatid="7951" lane="3" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:08.33" />
                    <SPLIT distance="150" swimtime="00:01:44.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="440" reactiontime="+83" swimtime="00:06:36.66" resultid="3911" heatid="8802" lane="6" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:01:37.47" />
                    <SPLIT distance="150" swimtime="00:02:31.88" />
                    <SPLIT distance="200" swimtime="00:03:25.43" />
                    <SPLIT distance="250" swimtime="00:04:21.01" />
                    <SPLIT distance="300" swimtime="00:05:18.64" />
                    <SPLIT distance="350" swimtime="00:05:58.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="390" reactiontime="+79" swimtime="00:01:26.92" resultid="3912" heatid="7990" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="634" reactiontime="+79" swimtime="00:05:00.91" resultid="3913" heatid="9047" lane="5" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:49.93" />
                    <SPLIT distance="200" swimtime="00:02:28.56" />
                    <SPLIT distance="250" swimtime="00:03:07.04" />
                    <SPLIT distance="300" swimtime="00:03:45.74" />
                    <SPLIT distance="350" swimtime="00:04:24.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-12-07" firstname="Jarosław" gender="M" lastname="Zadrożny" nation="POL" athleteid="3914">
              <RESULTS>
                <RESULT eventid="1076" points="388" reactiontime="+84" swimtime="00:00:33.14" resultid="3915" heatid="7691" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1156" points="321" swimtime="00:24:02.85" resultid="3916" heatid="8721" lane="1" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:23.60" />
                    <SPLIT distance="200" swimtime="00:02:54.92" />
                    <SPLIT distance="300" swimtime="00:04:30.27" />
                    <SPLIT distance="400" swimtime="00:06:06.96" />
                    <SPLIT distance="500" swimtime="00:07:43.88" />
                    <SPLIT distance="600" swimtime="00:09:21.06" />
                    <SPLIT distance="700" swimtime="00:10:58.21" />
                    <SPLIT distance="800" swimtime="00:12:37.31" />
                    <SPLIT distance="900" swimtime="00:14:16.08" />
                    <SPLIT distance="1000" swimtime="00:15:55.07" />
                    <SPLIT distance="1100" swimtime="00:17:33.50" />
                    <SPLIT distance="1200" swimtime="00:19:11.42" />
                    <SPLIT distance="1300" swimtime="00:20:49.65" />
                    <SPLIT distance="1400" swimtime="00:22:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="229" reactiontime="+98" swimtime="00:04:03.70" resultid="3917" heatid="7784" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.27" />
                    <SPLIT distance="100" swimtime="00:01:59.24" />
                    <SPLIT distance="150" swimtime="00:03:02.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="344" reactiontime="+95" swimtime="00:01:15.46" resultid="3918" heatid="7812" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="3919" heatid="7881" lane="2" />
                <RESULT eventid="1479" points="337" reactiontime="+95" swimtime="00:02:44.84" resultid="3920" heatid="7958" lane="2" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                    <SPLIT distance="100" swimtime="00:01:17.44" />
                    <SPLIT distance="150" swimtime="00:02:02.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="3921" heatid="8029" lane="3" />
                <RESULT eventid="1703" points="341" reactiontime="+98" swimtime="00:05:51.80" resultid="3922" heatid="9066" lane="7" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                    <SPLIT distance="100" swimtime="00:01:19.84" />
                    <SPLIT distance="150" swimtime="00:02:03.99" />
                    <SPLIT distance="200" swimtime="00:02:49.76" />
                    <SPLIT distance="250" swimtime="00:03:36.37" />
                    <SPLIT distance="300" swimtime="00:04:21.33" />
                    <SPLIT distance="350" swimtime="00:05:08.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="3923">
              <RESULTS>
                <RESULT eventid="1059" points="559" reactiontime="+103" swimtime="00:00:36.72" resultid="3924" heatid="7678" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1140" points="460" swimtime="00:14:29.45" resultid="3925" heatid="8714" lane="7" entrytime="00:13:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                    <SPLIT distance="100" swimtime="00:01:38.21" />
                    <SPLIT distance="200" swimtime="00:03:26.63" />
                    <SPLIT distance="300" swimtime="00:05:17.26" />
                    <SPLIT distance="400" swimtime="00:07:06.82" />
                    <SPLIT distance="500" swimtime="00:08:56.96" />
                    <SPLIT distance="600" swimtime="00:10:48.29" />
                    <SPLIT distance="700" swimtime="00:12:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="575" reactiontime="+81" swimtime="00:00:43.74" resultid="3926" heatid="7757" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1302" points="433" reactiontime="+101" swimtime="00:03:57.19" resultid="3927" heatid="7858" lane="6" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.50" />
                    <SPLIT distance="100" swimtime="00:01:52.23" />
                    <SPLIT distance="150" swimtime="00:02:55.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="539" reactiontime="+109" swimtime="00:00:41.93" resultid="3928" heatid="7899" lane="3" entrytime="00:00:41.13" />
                <RESULT eventid="1527" points="496" reactiontime="+110" swimtime="00:07:47.03" resultid="3929" heatid="8803" lane="6" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.57" />
                    <SPLIT distance="100" swimtime="00:01:55.38" />
                    <SPLIT distance="150" swimtime="00:02:53.44" />
                    <SPLIT distance="200" swimtime="00:03:52.74" />
                    <SPLIT distance="250" swimtime="00:04:58.23" />
                    <SPLIT distance="300" swimtime="00:06:02.36" />
                    <SPLIT distance="350" swimtime="00:06:55.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="424" reactiontime="+115" swimtime="00:01:44.65" resultid="3930" heatid="7988" lane="3" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="456" reactiontime="+114" swimtime="00:06:57.63" resultid="3931" heatid="9051" lane="8" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.14" />
                    <SPLIT distance="100" swimtime="00:01:35.64" />
                    <SPLIT distance="150" swimtime="00:02:29.65" />
                    <SPLIT distance="200" swimtime="00:03:23.67" />
                    <SPLIT distance="250" swimtime="00:04:17.83" />
                    <SPLIT distance="300" swimtime="00:05:12.25" />
                    <SPLIT distance="350" swimtime="00:06:06.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="3932">
              <RESULTS>
                <RESULT eventid="1092" points="508" reactiontime="+99" swimtime="00:03:14.59" resultid="3933" heatid="7713" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                    <SPLIT distance="100" swimtime="00:01:30.85" />
                    <SPLIT distance="150" swimtime="00:02:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="378" swimtime="00:13:28.57" resultid="3934" heatid="8716" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                    <SPLIT distance="100" swimtime="00:01:28.70" />
                    <SPLIT distance="200" swimtime="00:03:08.64" />
                    <SPLIT distance="300" swimtime="00:04:52.43" />
                    <SPLIT distance="400" swimtime="00:06:36.56" />
                    <SPLIT distance="500" swimtime="00:08:20.43" />
                    <SPLIT distance="600" swimtime="00:10:05.94" />
                    <SPLIT distance="700" swimtime="00:11:50.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="435" reactiontime="+93" swimtime="00:01:21.74" resultid="3935" heatid="7796" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="529" reactiontime="+93" swimtime="00:03:30.42" resultid="3936" heatid="7857" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="100" swimtime="00:01:34.53" />
                    <SPLIT distance="150" swimtime="00:02:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="470" reactiontime="+98" swimtime="00:00:40.05" resultid="3937" heatid="7897" lane="3" />
                <RESULT eventid="1463" points="406" reactiontime="+102" swimtime="00:03:02.01" resultid="3938" heatid="7943" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:25.71" />
                    <SPLIT distance="150" swimtime="00:02:15.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="494" reactiontime="+99" swimtime="00:01:29.52" resultid="3939" heatid="7987" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="450" reactiontime="+96" swimtime="00:06:13.50" resultid="3940" heatid="9053" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:24.34" />
                    <SPLIT distance="150" swimtime="00:02:12.42" />
                    <SPLIT distance="200" swimtime="00:03:01.20" />
                    <SPLIT distance="250" swimtime="00:03:50.00" />
                    <SPLIT distance="300" swimtime="00:04:39.62" />
                    <SPLIT distance="350" swimtime="00:05:28.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-15" firstname="Mariusz" gender="M" lastname="Kaliszyk" nation="POL" athleteid="3941">
              <RESULTS>
                <RESULT eventid="1076" points="721" reactiontime="+85" swimtime="00:00:26.49" resultid="3942" heatid="7704" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1190" points="682" reactiontime="+65" swimtime="00:00:30.83" resultid="3943" heatid="7774" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1415" points="659" reactiontime="+85" swimtime="00:00:28.87" resultid="3944" heatid="7918" lane="2" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-05-14" firstname="Piotr" gender="M" lastname="Kowalski" nation="POL" athleteid="3945">
              <RESULTS>
                <RESULT eventid="1076" points="387" reactiontime="+78" swimtime="00:00:32.54" resultid="3946" heatid="7688" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1190" points="234" reactiontime="+89" swimtime="00:00:44.03" resultid="3947" heatid="7766" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1254" points="307" reactiontime="+89" swimtime="00:01:16.19" resultid="3948" heatid="7809" lane="8" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="3949" heatid="7955" lane="2" entrytime="00:03:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-15" firstname="Monika" gender="F" lastname="Jaworska" nation="POL" athleteid="3950">
              <RESULTS>
                <RESULT eventid="1270" points="425" reactiontime="+81" swimtime="00:01:26.58" resultid="3951" heatid="7835" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="512" reactiontime="+80" swimtime="00:00:35.77" resultid="3952" heatid="7904" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1574" points="396" reactiontime="+77" swimtime="00:01:26.46" resultid="3953" heatid="7990" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-11-05" firstname="Aleksandra" gender="F" lastname="Jamrozik" nation="POL" athleteid="3954">
              <RESULTS>
                <RESULT eventid="1092" points="701" reactiontime="+80" swimtime="00:02:40.97" resultid="3955" heatid="7718" lane="3" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:01:15.96" />
                    <SPLIT distance="150" swimtime="00:02:03.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="572" reactiontime="+85" swimtime="00:10:59.77" resultid="3956" heatid="8712" lane="1" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:16.20" />
                    <SPLIT distance="150" swimtime="00:01:57.26" />
                    <SPLIT distance="200" swimtime="00:02:38.88" />
                    <SPLIT distance="250" swimtime="00:03:20.54" />
                    <SPLIT distance="300" swimtime="00:04:02.14" />
                    <SPLIT distance="350" swimtime="00:04:44.23" />
                    <SPLIT distance="400" swimtime="00:05:26.25" />
                    <SPLIT distance="450" swimtime="00:06:07.88" />
                    <SPLIT distance="500" swimtime="00:06:49.96" />
                    <SPLIT distance="550" swimtime="00:07:31.85" />
                    <SPLIT distance="600" swimtime="00:08:13.96" />
                    <SPLIT distance="650" swimtime="00:08:56.56" />
                    <SPLIT distance="700" swimtime="00:09:38.72" />
                    <SPLIT distance="750" swimtime="00:10:20.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="724" reactiontime="+68" swimtime="00:02:40.20" resultid="3957" heatid="8009" lane="7" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                    <SPLIT distance="150" swimtime="00:01:59.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="559" reactiontime="+78" swimtime="00:05:13.89" resultid="3958" heatid="9048" lane="6" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:14.84" />
                    <SPLIT distance="150" swimtime="00:01:54.58" />
                    <SPLIT distance="200" swimtime="00:02:34.33" />
                    <SPLIT distance="250" swimtime="00:03:14.82" />
                    <SPLIT distance="300" swimtime="00:03:55.45" />
                    <SPLIT distance="350" swimtime="00:04:35.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-03-21" firstname="Justyna" gender="F" lastname="Jamrozik" nation="POL" athleteid="3959">
              <RESULTS>
                <RESULT eventid="1206" points="540" reactiontime="+89" swimtime="00:03:08.64" resultid="3960" heatid="7783" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:01:30.85" />
                    <SPLIT distance="150" swimtime="00:02:19.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="511" reactiontime="+93" swimtime="00:01:21.81" resultid="3961" heatid="7835" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="520" reactiontime="+87" swimtime="00:01:27.82" resultid="3962" heatid="7879" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="509" reactiontime="+95" swimtime="00:00:36.39" resultid="3963" heatid="7903" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="3964" heatid="7990" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1639" points="490" reactiontime="+88" swimtime="00:00:40.05" resultid="3965" heatid="8027" lane="7" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-10-18" firstname="Dorota" gender="F" lastname="Widz- Szwarc" nation="POL" athleteid="3966">
              <RESULTS>
                <RESULT eventid="1059" points="438" reactiontime="+88" swimtime="00:00:36.54" resultid="3967" heatid="7675" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-03-21" firstname="Janusz" gender="M" lastname="Gołębiewski" nation="POL" athleteid="3968">
              <RESULTS>
                <RESULT eventid="1076" points="102" swimtime="00:01:00.22" resultid="3969" heatid="7684" lane="8" />
                <RESULT eventid="1222" status="DNF" swimtime="00:00:00.00" resultid="3970" heatid="7784" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="183" swimtime="00:01:02.21" resultid="3971" heatid="8029" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Masters Korona Kraków B" number="1">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+73" swimtime="00:01:48.52" resultid="3981" heatid="7974" lane="2" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.18" />
                    <SPLIT distance="100" swimtime="00:00:52.44" />
                    <SPLIT distance="150" swimtime="00:01:21.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3836" number="1" />
                    <RELAYPOSITION athleteid="3862" number="2" />
                    <RELAYPOSITION athleteid="3756" number="3" />
                    <RELAYPOSITION athleteid="3894" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1357" reactiontime="+66" swimtime="00:02:05.75" resultid="3982" heatid="7872" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3756" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3836" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="3853" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="3862" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Masters Korona Kraków C" number="1">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+84" swimtime="00:01:49.74" resultid="3983" heatid="7974" lane="3" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                    <SPLIT distance="100" swimtime="00:00:55.31" />
                    <SPLIT distance="150" swimtime="00:01:23.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3941" number="1" />
                    <RELAYPOSITION athleteid="3853" number="2" />
                    <RELAYPOSITION athleteid="3865" number="3" />
                    <RELAYPOSITION athleteid="3774" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Masters Korona Kraków D" number="1">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+98" swimtime="00:02:07.00" resultid="3984" heatid="7972" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:04.98" />
                    <SPLIT distance="150" swimtime="00:01:37.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3723" number="1" />
                    <RELAYPOSITION athleteid="3914" number="2" />
                    <RELAYPOSITION athleteid="3810" number="3" />
                    <RELAYPOSITION athleteid="3828" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1357" reactiontime="+62" swimtime="00:02:08.66" resultid="3985" heatid="7871" lane="8" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:35.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3941" number="1" />
                    <RELAYPOSITION athleteid="3865" number="2" />
                    <RELAYPOSITION athleteid="3828" number="3" />
                    <RELAYPOSITION athleteid="3810" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Masters Korona Kraków B" number="1">
              <RESULTS>
                <RESULT eventid="1495" reactiontime="+89" swimtime="00:02:17.87" resultid="3972" heatid="7969" lane="7" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:09.70" />
                    <SPLIT distance="150" swimtime="00:01:43.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3959" number="1" />
                    <RELAYPOSITION athleteid="3803" number="2" />
                    <RELAYPOSITION athleteid="3745" number="3" />
                    <RELAYPOSITION athleteid="3878" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" reactiontime="+65" swimtime="00:02:24.94" resultid="3973" heatid="7867" lane="5" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:01:51.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3841" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="3959" number="2" reactiontime="+74" />
                    <RELAYPOSITION athleteid="3887" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="3745" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Masters Korona Kraków D" number="1">
              <RESULTS>
                <RESULT eventid="1495" reactiontime="+75" swimtime="00:02:12.26" resultid="3986" heatid="7969" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:07.79" />
                    <SPLIT distance="150" swimtime="00:01:42.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3711" number="1" />
                    <RELAYPOSITION athleteid="3923" number="2" />
                    <RELAYPOSITION athleteid="3882" number="3" />
                    <RELAYPOSITION athleteid="3887" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" reactiontime="+61" swimtime="00:02:28.44" resultid="3987" heatid="7867" lane="2" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:18.73" />
                    <SPLIT distance="150" swimtime="00:01:54.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3711" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3882" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3878" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3932" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Masters Korona Kraków B" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+66" swimtime="00:01:56.63" resultid="3976" heatid="7737" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:00:56.97" />
                    <SPLIT distance="150" swimtime="00:01:30.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3841" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3862" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="3745" number="3" reactiontime="+83" />
                    <RELAYPOSITION athleteid="3836" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" reactiontime="+91" swimtime="00:02:17.15" resultid="3977" heatid="8052" lane="7" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3745" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="3959" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3853" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="3836" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Masters Korona Kraków C" number="1">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+66" swimtime="00:02:06.83" resultid="3974" heatid="8052" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:07.91" />
                    <SPLIT distance="150" swimtime="00:01:36.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3841" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3865" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="3941" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3887" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1124" reactiontime="+73" swimtime="00:01:53.49" resultid="3975" heatid="7737" lane="6" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:00:57.35" />
                    <SPLIT distance="150" swimtime="00:01:27.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3711" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3941" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3887" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3774" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Masters Korona Kraków D" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+92" swimtime="00:02:07.59" resultid="3978" heatid="7737" lane="8" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                    <SPLIT distance="100" swimtime="00:01:04.30" />
                    <SPLIT distance="150" swimtime="00:01:38.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3828" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="3932" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3882" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3865" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" reactiontime="+69" swimtime="00:02:19.24" resultid="3979" heatid="8051" lane="7" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:17.46" />
                    <SPLIT distance="150" swimtime="00:01:47.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3711" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3882" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="3828" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3723" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Masters Korona Kraków E" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+107" swimtime="00:02:23.75" resultid="3980" heatid="7734" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="150" swimtime="00:01:50.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3923" number="1" reactiontime="+107" />
                    <RELAYPOSITION athleteid="3728" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3798" number="3" reactiontime="+90" />
                    <RELAYPOSITION athleteid="3810" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAKRA" nation="POL" region="03" clubid="3163" name="Masters Kraśnik">
          <CONTACT city="Kraśnik" email="jurek@krasnik.info" internet="www.masterskrasnik.za.pl" name="Michalczyk Jerzy" phone="601698977" street="Żwirki i Wigury 2" zip="23-210" />
          <ATHLETES>
            <ATHLETE birthdate="1975-02-09" firstname="Marcin" gender="M" lastname="Mazurek" nation="POL" athleteid="3164">
              <RESULTS>
                <RESULT eventid="1254" points="317" reactiontime="+93" swimtime="00:01:15.39" resultid="3166" heatid="7811" lane="7" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="272" reactiontime="+87" swimtime="00:02:51.97" resultid="3167" heatid="7959" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                    <SPLIT distance="150" swimtime="00:02:05.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="301" reactiontime="+108" swimtime="00:00:35.39" resultid="6226" heatid="7699" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-04" firstname="Zdzisław" gender="M" lastname="Bąk" nation="POL" athleteid="3168">
              <RESULTS>
                <RESULT eventid="1076" points="473" reactiontime="+96" swimtime="00:00:32.60" resultid="3169" heatid="7690" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1254" points="421" reactiontime="+112" swimtime="00:01:15.25" resultid="3170" heatid="7810" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="347" reactiontime="+105" swimtime="00:02:58.86" resultid="3171" heatid="7953" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:11.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="3172">
              <RESULTS>
                <RESULT comment="G8 - Ukończenie wyścigu nie w położeniu na plecach  (Czas: 17:51)" eventid="1108" reactiontime="+93" status="DSQ" swimtime="00:03:55.62" resultid="3173" heatid="7721" lane="1" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.34" />
                    <SPLIT distance="100" swimtime="00:01:47.14" />
                    <SPLIT distance="150" swimtime="00:03:00.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="380" reactiontime="+71" swimtime="00:00:43.43" resultid="3174" heatid="7766" lane="1" entrytime="00:00:47.20" />
                <RESULT eventid="1415" points="268" reactiontime="+84" swimtime="00:00:44.20" resultid="3175" heatid="7907" lane="5" entrytime="00:00:49.20" />
                <RESULT eventid="1543" points="288" reactiontime="+96" swimtime="00:08:10.67" resultid="3176" heatid="8811" lane="7" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.91" />
                    <SPLIT distance="100" swimtime="00:01:54.02" />
                    <SPLIT distance="150" swimtime="00:02:55.79" />
                    <SPLIT distance="200" swimtime="00:03:54.96" />
                    <SPLIT distance="250" swimtime="00:05:10.29" />
                    <SPLIT distance="300" swimtime="00:06:22.73" />
                    <SPLIT distance="350" swimtime="00:07:18.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="356" reactiontime="+75" swimtime="00:03:38.66" resultid="3177" heatid="8011" lane="4" entrytime="00:03:57.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.89" />
                    <SPLIT distance="100" swimtime="00:01:46.76" />
                    <SPLIT distance="150" swimtime="00:02:43.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-09-07" firstname="Andrzej" gender="M" lastname="Cis" nation="POL" athleteid="3178">
              <RESULTS>
                <RESULT eventid="1076" points="568" reactiontime="+76" swimtime="00:00:30.68" resultid="3179" heatid="7695" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1108" points="398" reactiontime="+69" swimtime="00:03:14.27" resultid="3180" heatid="7724" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="100" swimtime="00:01:32.59" />
                    <SPLIT distance="150" swimtime="00:02:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="460" reactiontime="+64" swimtime="00:00:38.06" resultid="3181" heatid="7770" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1254" points="543" reactiontime="+64" swimtime="00:01:09.14" resultid="3182" heatid="7813" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1415" reactiontime="+41" status="DSQ" swimtime="00:00:34.79" resultid="3183" heatid="7911" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1543" points="304" reactiontime="+78" swimtime="00:07:38.62" resultid="3184" heatid="8810" lane="3" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                    <SPLIT distance="100" swimtime="00:01:46.56" />
                    <SPLIT distance="150" swimtime="00:02:47.17" />
                    <SPLIT distance="200" swimtime="00:03:47.67" />
                    <SPLIT distance="250" swimtime="00:04:52.79" />
                    <SPLIT distance="300" swimtime="00:05:57.67" />
                    <SPLIT distance="350" swimtime="00:06:50.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="419" reactiontime="+72" swimtime="00:03:13.67" resultid="3185" heatid="8013" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:36.24" />
                    <SPLIT distance="100" swimtime="00:02:27.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-27" firstname="Janusz" gender="M" lastname="Wasiuk" nation="POL" athleteid="3186">
              <RESULTS>
                <RESULT eventid="1222" points="495" reactiontime="+110" swimtime="00:03:41.11" resultid="3188" heatid="7787" lane="2" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.05" />
                    <SPLIT distance="100" swimtime="00:01:44.68" />
                    <SPLIT distance="150" swimtime="00:02:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="348" reactiontime="+141" swimtime="00:03:47.08" resultid="3189" heatid="7859" lane="3" entrytime="00:04:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.87" />
                    <SPLIT distance="100" swimtime="00:01:47.62" />
                    <SPLIT distance="150" swimtime="00:02:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="485" reactiontime="+109" swimtime="00:01:39.43" resultid="3190" heatid="7884" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="330" reactiontime="+126" swimtime="00:08:24.63" resultid="3191" heatid="8812" lane="4" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.80" />
                    <SPLIT distance="100" swimtime="00:01:48.17" />
                    <SPLIT distance="150" swimtime="00:03:05.61" />
                    <SPLIT distance="200" swimtime="00:04:20.79" />
                    <SPLIT distance="250" swimtime="00:05:24.26" />
                    <SPLIT distance="300" swimtime="00:06:26.86" />
                    <SPLIT distance="350" swimtime="00:07:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="268" reactiontime="+134" swimtime="00:01:45.93" resultid="3192" heatid="7993" lane="1" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="474" reactiontime="+104" swimtime="00:00:43.34" resultid="3193" heatid="8032" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="3194">
              <RESULTS>
                <RESULT eventid="1076" points="260" reactiontime="+95" swimtime="00:00:40.84" resultid="3195" heatid="7687" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1222" points="320" reactiontime="+90" swimtime="00:03:57.74" resultid="3196" heatid="7786" lane="7" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.75" />
                    <SPLIT distance="100" swimtime="00:01:53.21" />
                    <SPLIT distance="150" swimtime="00:02:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="274" reactiontime="+90" swimtime="00:01:44.88" resultid="3197" heatid="7883" lane="7" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="222" reactiontime="+85" swimtime="00:00:47.07" resultid="3198" heatid="7907" lane="4" entrytime="00:00:48.00" />
                <RESULT eventid="1591" points="173" reactiontime="+86" swimtime="00:01:56.18" resultid="3199" heatid="7993" lane="3" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-12-19" firstname="Waldemar" gender="M" lastname="Rusowicz" nation="POL" athleteid="3200">
              <RESULTS>
                <RESULT eventid="1108" points="242" reactiontime="+88" swimtime="00:03:57.80" resultid="3201" heatid="7720" lane="6" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.88" />
                    <SPLIT distance="100" swimtime="00:02:02.37" />
                    <SPLIT distance="150" swimtime="00:03:02.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="218" reactiontime="+83" swimtime="00:00:52.24" resultid="3202" heatid="7767" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1222" points="413" reactiontime="+88" swimtime="00:03:38.25" resultid="3203" heatid="7788" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                    <SPLIT distance="100" swimtime="00:01:44.98" />
                    <SPLIT distance="150" swimtime="00:02:42.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="309" reactiontime="+94" swimtime="00:01:40.68" resultid="3204" heatid="7885" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="220" reactiontime="+81" swimtime="00:01:53.69" resultid="3205" heatid="7934" lane="3" entrytime="00:01:45.00" />
                <RESULT eventid="1623" points="340" reactiontime="+75" swimtime="00:03:42.06" resultid="3206" heatid="8011" lane="2" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.69" />
                    <SPLIT distance="100" swimtime="00:01:49.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="300" reactiontime="+90" swimtime="00:00:45.52" resultid="3207" heatid="8033" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EULVI" nation="UKR" clubid="3308" name="Masters Swimming Club Euro Lviv" shortname="Masters SC Euro Lviv">
          <CONTACT city="Lviv" email="riff@mail.lviv.ua" fax="+380322430304" name="Ruslan Friauf" phone="+380676734796" street="Karpincya, 18A/3" zip="79012" />
          <ATHLETES>
            <ATHLETE birthdate="1932-06-01" firstname="Serhiy" gender="M" lastname="Simankov" nation="UKR" athleteid="3309">
              <RESULTS>
                <RESULT eventid="1076" points="511" reactiontime="+120" swimtime="00:00:41.56" resultid="3310" heatid="7686" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1415" points="714" reactiontime="+123" swimtime="00:00:49.68" resultid="3311" heatid="7907" lane="8" entrytime="00:00:52.00" />
                <RESULT comment="M8 - Przenoszenie ramion do przodu pod powierzchnią wody podczas ostatniego cyklu pracy ramion przed nawrotem lub na zakończenie wyścigu  (Czas: 9:17)" eventid="1591" reactiontime="+124" status="DSQ" swimtime="00:02:06.10" resultid="3312" heatid="7992" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-11-07" firstname="Bohdan" gender="M" lastname="Yatsura" nation="UKR" athleteid="3313">
              <RESULTS>
                <RESULT eventid="1076" points="415" reactiontime="+89" swimtime="00:00:34.96" resultid="3314" heatid="7690" lane="1" entrytime="00:00:34.01" />
                <RESULT eventid="1415" points="352" reactiontime="+76" swimtime="00:00:40.38" resultid="3315" heatid="7909" lane="4" entrytime="00:00:39.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-04-06" firstname="Sergiy" gender="M" lastname="Mashkin" nation="UKR" athleteid="3316">
              <RESULTS>
                <RESULT eventid="1190" points="728" reactiontime="+77" swimtime="00:00:34.98" resultid="3317" heatid="7772" lane="8" entrytime="00:00:35.05" />
                <RESULT eventid="1286" points="748" reactiontime="+81" swimtime="00:01:16.18" resultid="3318" heatid="7850" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="739" reactiontime="+87" swimtime="00:01:15.91" resultid="3319" heatid="7939" lane="6" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="810" reactiontime="+79" swimtime="00:02:46.30" resultid="3320" heatid="8017" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:20.78" />
                    <SPLIT distance="150" swimtime="00:02:03.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-11" firstname="Nataliya" gender="F" lastname="Hertsyk" nation="UKR" athleteid="3321">
              <RESULTS>
                <RESULT eventid="1059" points="405" reactiontime="+117" swimtime="00:00:38.49" resultid="3322" heatid="7676" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1399" points="402" reactiontime="+101" swimtime="00:00:42.20" resultid="3323" heatid="7901" lane="8" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-08-08" firstname="Andrii" gender="M" lastname="Hertsyk" nation="UKR" athleteid="3324">
              <RESULTS>
                <RESULT eventid="1383" points="465" reactiontime="+89" swimtime="00:01:29.76" resultid="3325" heatid="7887" lane="4" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="454" reactiontime="+98" swimtime="00:00:40.80" resultid="3326" heatid="8037" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-13" firstname="Oleksandr" gender="M" lastname="Syrbu" nation="UKR" athleteid="3327">
              <RESULTS>
                <RESULT eventid="1076" points="793" reactiontime="+73" swimtime="00:00:25.67" resultid="3328" heatid="7711" lane="7" entrytime="00:00:25.80" />
                <RESULT eventid="1254" points="765" reactiontime="+76" swimtime="00:00:56.91" resultid="3329" heatid="7824" lane="7" entrytime="00:00:57.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="795" reactiontime="+76" swimtime="00:00:27.12" resultid="3330" heatid="7924" lane="7" entrytime="00:00:27.40" />
                <RESULT eventid="1479" points="572" reactiontime="+80" swimtime="00:02:16.10" resultid="3331" heatid="7966" lane="4" entrytime="00:02:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:06.85" />
                    <SPLIT distance="150" swimtime="00:01:41.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="656" reactiontime="+77" swimtime="00:01:05.14" resultid="3332" heatid="8002" lane="7" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-06-05" firstname="Mykhailo" gender="M" lastname="Shelest" nation="UKR" athleteid="3333">
              <RESULTS>
                <RESULT eventid="1383" points="495" reactiontime="+96" swimtime="00:01:26.09" resultid="3334" heatid="7889" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="531" reactiontime="+92" swimtime="00:00:37.65" resultid="3335" heatid="8040" lane="6" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-18" firstname="Dmytro" gender="M" lastname="Melnyk" nation="UKR" athleteid="3336">
              <RESULTS>
                <RESULT eventid="1076" points="751" reactiontime="+69" swimtime="00:00:26.09" resultid="3337" heatid="7709" lane="2" entrytime="00:00:26.45" />
                <RESULT eventid="1383" points="633" reactiontime="+69" swimtime="00:01:14.56" resultid="3338" heatid="7894" lane="1" entrytime="00:01:15.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="645" reactiontime="+64" swimtime="00:00:33.40" resultid="3339" heatid="8046" lane="1" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-06-23" firstname="Nadiya" gender="F" lastname="Sannikova" nation="UKR" athleteid="3340">
              <RESULTS>
                <RESULT eventid="1639" points="465" reactiontime="+104" swimtime="00:00:48.45" resultid="3341" heatid="8024" lane="1" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-02" firstname="Serhiy" gender="M" lastname="Zhykh" nation="UKR" athleteid="3342">
              <RESULTS>
                <RESULT eventid="1076" points="657" reactiontime="+81" swimtime="00:00:29.22" resultid="3343" heatid="7702" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="1190" points="645" reactiontime="+80" swimtime="00:00:33.99" resultid="3344" heatid="7774" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="3345" heatid="7850" lane="4" entrytime="00:01:12.50" />
                <RESULT eventid="1415" points="651" reactiontime="+82" swimtime="00:00:31.78" resultid="3346" heatid="7919" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1447" points="663" reactiontime="+67" swimtime="00:01:14.34" resultid="3347" heatid="7940" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-23" firstname="Oleksandr" gender="M" lastname="Shavrov" nation="UKR" athleteid="3348">
              <RESULTS>
                <RESULT eventid="1222" points="572" reactiontime="+77" swimtime="00:02:51.60" resultid="3349" heatid="7794" lane="7" entrytime="00:02:54.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                    <SPLIT distance="150" swimtime="00:02:05.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="604" reactiontime="+77" swimtime="00:01:15.71" resultid="3350" heatid="7893" lane="7" entrytime="00:01:19.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="609" reactiontime="+75" swimtime="00:00:34.06" resultid="3351" heatid="8044" lane="3" entrytime="00:00:34.65" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-13" firstname="Bogdan" gender="M" lastname="Osidach" nation="UKR" athleteid="3352">
              <RESULTS>
                <RESULT eventid="1076" points="404" reactiontime="+88" swimtime="00:00:32.08" resultid="3353" heatid="7697" lane="3" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-05-09" firstname="Lidiya" gender="F" lastname="Tymoshenko" nation="UKR" athleteid="3354">
              <RESULTS>
                <RESULT eventid="1059" points="318" reactiontime="+111" swimtime="00:00:47.10" resultid="3355" heatid="7674" lane="8" entrytime="00:00:44.60" />
                <RESULT eventid="1173" points="251" reactiontime="+91" swimtime="00:01:02.91" resultid="3356" heatid="7754" lane="6" entrytime="00:01:01.12" />
                <RESULT eventid="1639" points="385" reactiontime="+108" swimtime="00:00:53.02" resultid="3357" heatid="8022" lane="6" entrytime="00:00:52.59" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-07-08" firstname="Ihor" gender="M" lastname="Rudnyk" nation="UKR" athleteid="3358">
              <RESULTS>
                <RESULT eventid="1076" points="475" reactiontime="+95" swimtime="00:00:32.55" resultid="3359" heatid="7694" lane="7" entrytime="00:00:31.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="Friauf" nation="UKR" athleteid="3360">
              <RESULTS>
                <RESULT comment="G8 - Ukończenie wyścigu nie w położeniu na plecach  (Czas: 18:11)" eventid="1108" reactiontime="+75" status="DSQ" swimtime="00:03:01.38" resultid="3361" heatid="7727" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:24.24" />
                    <SPLIT distance="150" swimtime="00:02:15.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="414" reactiontime="+74" swimtime="00:00:36.42" resultid="3362" heatid="7771" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1286" points="467" reactiontime="+77" swimtime="00:01:17.08" resultid="3363" heatid="7843" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="3364" heatid="7937" lane="3" entrytime="00:01:23.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="3365" heatid="8041" lane="8" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-11-30" firstname="Tetiana" gender="F" lastname="Kozakova" nation="UKR" athleteid="3377">
              <RESULTS>
                <RESULT eventid="1173" points="441" reactiontime="+108" swimtime="00:00:52.13" resultid="3378" heatid="7755" lane="6" entrytime="00:00:51.00" />
                <RESULT eventid="1270" points="317" reactiontime="+108" swimtime="00:01:55.99" resultid="3379" heatid="7828" lane="8" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-10" firstname="Serhiy" gender="M" lastname="Fedorov" nation="UKR" athleteid="3380">
              <RESULTS>
                <RESULT eventid="1076" points="749" status="EXH" swimtime="00:00:28.71" resultid="3381" heatid="7699" lane="8" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-03" firstname="Romana" gender="F" lastname="Sirenko" nation="UKR" athleteid="3382">
              <RESULTS>
                <RESULT eventid="1092" points="511" reactiontime="+116" swimtime="00:03:01.61" resultid="3383" heatid="7716" lane="6" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:24.36" />
                    <SPLIT distance="150" swimtime="00:02:17.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="562" reactiontime="+108" swimtime="00:01:22.26" resultid="3384" heatid="7834" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="582" reactiontime="+107" swimtime="00:00:35.35" resultid="3385" heatid="7902" lane="3" entrytime="00:00:35.50" />
                <RESULT eventid="1527" points="480" reactiontime="+99" swimtime="00:06:42.93" resultid="3386" heatid="8803" lane="3" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                    <SPLIT distance="100" swimtime="00:01:39.28" />
                    <SPLIT distance="150" swimtime="00:02:28.76" />
                    <SPLIT distance="200" swimtime="00:03:18.13" />
                    <SPLIT distance="250" swimtime="00:04:13.67" />
                    <SPLIT distance="300" swimtime="00:05:09.50" />
                    <SPLIT distance="350" swimtime="00:05:56.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="411" reactiontime="+106" swimtime="00:01:27.85" resultid="3387" heatid="7989" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-11-13" firstname="Ihor" gender="M" lastname="Yaskevych" nation="UKR" athleteid="3388">
              <RESULTS>
                <RESULT eventid="1383" points="481" reactiontime="+82" swimtime="00:01:25.79" resultid="3389" heatid="7888" lane="4" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="492" reactiontime="+81" swimtime="00:00:38.85" resultid="3390" heatid="8039" lane="6" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-10-14" firstname="Stepan" gender="M" lastname="Delyatynskyy" nation="UKR" athleteid="3391">
              <RESULTS>
                <RESULT eventid="1076" points="566" reactiontime="+81" swimtime="00:00:29.22" resultid="3392" heatid="7703" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1254" points="518" reactiontime="+82" swimtime="00:01:05.88" resultid="3393" heatid="7818" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="466" reactiontime="+78" swimtime="00:00:39.55" resultid="3394" heatid="8040" lane="2" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-05" firstname="Lyudmyla" gender="F" lastname="Khiresh" nation="UKR" athleteid="3395">
              <RESULTS>
                <RESULT eventid="1059" points="632" reactiontime="+91" swimtime="00:00:35.24" resultid="3396" heatid="7677" lane="3" entrytime="00:00:35.50" />
                <RESULT eventid="1173" points="793" reactiontime="+93" swimtime="00:00:39.30" resultid="3397" heatid="7758" lane="6" entrytime="00:00:39.50" />
                <RESULT eventid="1270" points="739" reactiontime="+92" swimtime="00:01:25.67" resultid="3398" heatid="7831" lane="4" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="814" reactiontime="+87" swimtime="00:01:25.41" resultid="3399" heatid="7929" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-03-29" firstname="Tetyana" gender="F" lastname="Zelikova" nation="UKR" athleteid="3400">
              <RESULTS>
                <RESULT eventid="1639" points="446" reactiontime="+99" swimtime="00:00:49.14" resultid="3401" heatid="8024" lane="4" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-27" firstname="Iurii" gender="M" lastname="Martyniuk" nation="UKR" athleteid="3402">
              <RESULTS>
                <RESULT eventid="1076" points="467" reactiontime="+92" swimtime="00:00:30.61" resultid="3403" heatid="7700" lane="3" entrytime="00:00:29.27" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="3404" heatid="7815" lane="8" entrytime="00:01:08.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-06" firstname="Yuriy" gender="M" lastname="Chyrkov" nation="UKR" athleteid="3405">
              <RESULTS>
                <RESULT eventid="1076" points="583" reactiontime="+103" swimtime="00:00:32.31" resultid="3406" heatid="7693" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1108" points="554" reactiontime="+109" swimtime="00:03:19.87" resultid="3407" heatid="7724" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.01" />
                    <SPLIT distance="100" swimtime="00:01:33.81" />
                    <SPLIT distance="150" swimtime="00:02:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="523" reactiontime="+70" swimtime="00:00:41.14" resultid="3408" heatid="7769" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1254" points="528" reactiontime="+93" swimtime="00:01:14.05" resultid="3409" heatid="7811" lane="3" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="500" reactiontime="+75" swimtime="00:01:31.57" resultid="3410" heatid="7936" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G3 - Nieutrzymanie pozycji na plecach (z wyjątkiem wykonania cyklu nawrotu)  (Czas: 10:30)" eventid="1623" reactiontime="+72" status="DSQ" swimtime="00:03:24.53" resultid="3411" heatid="8012" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                    <SPLIT distance="100" swimtime="00:01:41.67" />
                    <SPLIT distance="150" swimtime="00:02:35.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-05-31" firstname="Zenoviy" gender="M" lastname="Kushnir" nation="UKR" athleteid="3412">
              <RESULTS>
                <RESULT eventid="1190" points="208" reactiontime="+97" swimtime="00:00:56.22" resultid="3413" heatid="7764" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="1447" points="196" reactiontime="+88" swimtime="00:02:04.41" resultid="3414" heatid="7933" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="205" reactiontime="+90" swimtime="00:04:27.01" resultid="3415" heatid="8011" lane="7" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.85" />
                    <SPLIT distance="100" swimtime="00:02:13.93" />
                    <SPLIT distance="150" swimtime="00:03:23.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-06" firstname="Mariia" gender="F" lastname="Vasylko" nation="UKR" athleteid="3416">
              <RESULTS>
                <RESULT eventid="1173" points="320" reactiontime="+91" swimtime="00:00:48.52" resultid="3417" heatid="7754" lane="5" entrytime="00:00:56.00" />
                <RESULT eventid="1270" status="DNS" swimtime="00:00:00.00" resultid="3418" heatid="7830" lane="8" entrytime="00:01:36.00" />
                <RESULT eventid="1639" status="DNS" swimtime="00:00:00.00" resultid="3419" heatid="8025" lane="1" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-10-27" firstname="Yuriy" gender="M" lastname="Denisov" nation="UKR" athleteid="3420">
              <RESULTS>
                <RESULT eventid="1076" points="489" reactiontime="+110" swimtime="00:00:33.09" resultid="3421" heatid="7694" lane="2" entrytime="00:00:31.58" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-02-10" firstname="Taras" gender="M" lastname="Babyak" nation="UKR" athleteid="3422">
              <RESULTS>
                <RESULT eventid="1076" points="539" reactiontime="+93" swimtime="00:00:28.05" resultid="3423" heatid="7702" lane="4" entrytime="00:00:28.50" />
                <RESULT eventid="1254" points="454" reactiontime="+101" swimtime="00:01:03.20" resultid="3424" heatid="7813" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-03-11" firstname="Taras" gender="M" lastname="Kunets" nation="UKR" athleteid="3425">
              <RESULTS>
                <RESULT eventid="1076" points="549" reactiontime="+89" swimtime="00:00:27.89" resultid="3426" heatid="7702" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="1190" points="349" reactiontime="+91" swimtime="00:00:35.56" resultid="3427" heatid="7773" lane="6" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-11-09" firstname="Ostap" gender="M" lastname="Kunets" nation="UKR" athleteid="3428">
              <RESULTS>
                <RESULT eventid="1076" points="445" reactiontime="+97" swimtime="00:00:29.91" resultid="3429" heatid="7702" lane="6" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-28" firstname="Nina" gender="F" lastname="Golub" nation="UKR" athleteid="3430">
              <RESULTS>
                <RESULT eventid="1059" points="180" reactiontime="+111" swimtime="00:00:58.99" resultid="3431" heatid="7672" lane="6" entrytime="00:00:54.49" />
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="3432" heatid="8716" lane="5" entrytime="00:20:45.31" />
                <RESULT eventid="1238" points="196" reactiontime="+117" swimtime="00:02:08.51" resultid="3433" heatid="7797" lane="2" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="177" reactiontime="+126" swimtime="00:04:58.47" resultid="3434" heatid="7944" lane="2" entrytime="00:04:44.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.70" />
                    <SPLIT distance="100" swimtime="00:02:23.04" />
                    <SPLIT distance="150" swimtime="00:03:41.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" status="WDR" swimtime="00:00:00.00" resultid="3435" entrytime="00:09:59.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-09-04" firstname="Oleksandra" gender="F" lastname="Galkina" nation="UKR" athleteid="3436">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="3437" heatid="7673" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-05" firstname="Mykhailo" gender="M" lastname="Galkin" nation="UKR" athleteid="3438">
              <RESULTS>
                <RESULT eventid="1190" points="465" reactiontime="+79" swimtime="00:00:42.99" resultid="3439" heatid="7767" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1447" points="443" reactiontime="+83" swimtime="00:01:34.86" resultid="3440" heatid="7935" lane="7" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="523" reactiontime="+121" swimtime="00:03:01.14" resultid="3441" heatid="7956" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                    <SPLIT distance="100" swimtime="00:01:30.19" />
                    <SPLIT distance="150" swimtime="00:02:16.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="431" reactiontime="+87" swimtime="00:03:28.56" resultid="3442" heatid="8012" lane="3" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.15" />
                    <SPLIT distance="100" swimtime="00:01:43.44" />
                    <SPLIT distance="150" swimtime="00:02:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="3443" heatid="9067" lane="2" entrytime="00:06:06.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="MSC Euro Lviv A">
              <RESULTS>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="8772" heatid="7970" lane="8">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3422" number="1" />
                    <RELAYPOSITION athleteid="3428" number="2" />
                    <RELAYPOSITION athleteid="3425" number="3" />
                    <RELAYPOSITION athleteid="3336" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="MSC Euro Lviv C">
              <RESULTS>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="8769" heatid="7869" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3342" number="1" />
                    <RELAYPOSITION athleteid="3348" number="2" />
                    <RELAYPOSITION athleteid="3360" number="3" />
                    <RELAYPOSITION athleteid="3391" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="MSC Euro Lviv D">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+78" status="EXH" swimtime="00:02:06.17" resultid="8768" heatid="7872" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:07.62" />
                    <SPLIT distance="150" swimtime="00:01:34.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3316" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3336" number="2" reactiontime="+5" />
                    <RELAYPOSITION athleteid="3327" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3405" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" reactiontime="+78" status="EXH" swimtime="00:01:52.36" resultid="8771" heatid="7973" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                    <SPLIT distance="100" swimtime="00:00:57.60" />
                    <SPLIT distance="150" swimtime="00:01:26.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3391" number="1" />
                    <RELAYPOSITION athleteid="3380" number="2" />
                    <RELAYPOSITION athleteid="3316" number="3" />
                    <RELAYPOSITION athleteid="3327" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="MSC Euro Lviv D">
              <RESULTS>
                <RESULT eventid="1334" reactiontime="+82" status="EXH" swimtime="00:02:38.97" resultid="8762" heatid="7866" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:27.37" />
                    <SPLIT distance="150" swimtime="00:02:02.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3395" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3400" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="3382" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3321" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" name="MSC Euro Lviv E">
              <RESULTS>
                <RESULT eventid="1495" reactiontime="+93" status="EXH" swimtime="00:02:54.94" resultid="8770" heatid="7968" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:32.29" />
                    <SPLIT distance="150" swimtime="00:02:16.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3395" number="1" />
                    <RELAYPOSITION athleteid="3430" number="2" />
                    <RELAYPOSITION athleteid="3354" number="3" />
                    <RELAYPOSITION athleteid="3321" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="MSC Euro Lviv D">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+87" status="EXH" swimtime="00:02:07.24" resultid="8642" heatid="7736" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                    <SPLIT distance="100" swimtime="00:01:04.71" />
                    <SPLIT distance="150" swimtime="00:01:38.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3316" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3395" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3382" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="3342" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="X" name="MSC Euro Lviv F">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+108" status="EXH" swimtime="00:03:01.71" resultid="8641" heatid="7734" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:33.77" />
                    <SPLIT distance="150" swimtime="00:02:19.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3438" number="1" reactiontime="+108" />
                    <RELAYPOSITION athleteid="3430" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3354" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="3309" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00908" nation="POL" region="08" clubid="2771" name="Motyl Senior MOSiR St. Wola">
          <CONTACT city="Stalowa Wola" internet="lorkowska@wp.pl" name="Chmielewski Andrzej" phone="15-8422562 wew.45" state="PODK" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1970-06-07" firstname="Wiesław" gender="M" lastname="Bar" nation="POL" athleteid="2772">
              <RESULTS>
                <RESULT eventid="1076" points="645" reactiontime="+91" swimtime="00:00:27.50" resultid="2773" heatid="7706" lane="7" entrytime="00:00:27.44" />
                <RESULT eventid="1156" points="547" swimtime="00:20:18.68" resultid="2774" heatid="8718" lane="8" entrytime="00:21:19.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="200" swimtime="00:02:31.66" />
                    <SPLIT distance="300" swimtime="00:03:51.24" />
                    <SPLIT distance="400" swimtime="00:05:11.36" />
                    <SPLIT distance="500" swimtime="00:06:32.74" />
                    <SPLIT distance="600" swimtime="00:07:54.11" />
                    <SPLIT distance="700" swimtime="00:09:16.04" />
                    <SPLIT distance="800" swimtime="00:10:38.26" />
                    <SPLIT distance="1000" swimtime="00:13:23.97" />
                    <SPLIT distance="1100" swimtime="00:14:47.55" />
                    <SPLIT distance="1200" swimtime="00:16:10.64" />
                    <SPLIT distance="1300" swimtime="00:17:35.34" />
                    <SPLIT distance="1400" swimtime="00:18:59.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="605" reactiontime="+86" swimtime="00:01:01.54" resultid="2775" heatid="7821" lane="8" entrytime="00:01:01.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="601" reactiontime="+89" swimtime="00:01:10.86" resultid="2776" heatid="7851" lane="8" entrytime="00:01:12.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="540" reactiontime="+70" swimtime="00:01:12.51" resultid="2777" heatid="7939" lane="8" entrytime="00:01:16.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="560" reactiontime="+98" swimtime="00:02:17.10" resultid="2778" heatid="7963" lane="5" entrytime="00:02:18.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:07.65" />
                    <SPLIT distance="150" swimtime="00:01:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="462" reactiontime="+91" swimtime="00:01:13.24" resultid="2779" heatid="7999" lane="8" entrytime="00:01:12.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="553" reactiontime="+90" swimtime="00:04:53.21" resultid="2780" heatid="9062" lane="6" entrytime="00:05:03.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:10.43" />
                    <SPLIT distance="150" swimtime="00:01:48.50" />
                    <SPLIT distance="200" swimtime="00:02:25.96" />
                    <SPLIT distance="250" swimtime="00:03:03.91" />
                    <SPLIT distance="300" swimtime="00:03:41.00" />
                    <SPLIT distance="350" swimtime="00:04:17.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="2781">
              <RESULTS>
                <RESULT eventid="1076" points="753" reactiontime="+86" swimtime="00:00:26.07" resultid="2782" heatid="7708" lane="6" entrytime="00:00:26.69" />
                <RESULT eventid="1108" points="637" reactiontime="+91" swimtime="00:02:27.96" resultid="2783" heatid="7730" lane="4" entrytime="00:02:33.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:08.31" />
                    <SPLIT distance="150" swimtime="00:01:53.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="743" reactiontime="+77" swimtime="00:00:29.96" resultid="2784" heatid="7776" lane="8" entrytime="00:00:30.12" />
                <RESULT eventid="1254" points="703" reactiontime="+84" swimtime="00:00:57.82" resultid="2785" heatid="7822" lane="4" entrytime="00:00:59.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="723" reactiontime="+76" swimtime="00:01:05.86" resultid="2786" heatid="7942" lane="7" entrytime="00:01:05.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="696" reactiontime="+80" swimtime="00:02:26.63" resultid="2787" heatid="8019" lane="7" entrytime="00:02:28.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:10.56" />
                    <SPLIT distance="150" swimtime="00:01:48.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="492" reactiontime="+88" swimtime="00:00:36.57" resultid="2788" heatid="8039" lane="5" entrytime="00:00:38.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="2789">
              <RESULTS>
                <RESULT eventid="1076" points="826" reactiontime="+72" swimtime="00:00:25.32" resultid="2790" heatid="7709" lane="1" entrytime="00:00:26.50" />
                <RESULT eventid="1108" points="847" reactiontime="+72" swimtime="00:02:15.14" resultid="2791" heatid="7732" lane="4" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="100" swimtime="00:01:04.58" />
                    <SPLIT distance="150" swimtime="00:01:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="853" reactiontime="+73" swimtime="00:01:03.06" resultid="2792" heatid="7842" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="739" reactiontime="+77" swimtime="00:02:19.38" resultid="2793" heatid="7865" lane="4" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:07.07" />
                    <SPLIT distance="150" swimtime="00:01:43.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="800" reactiontime="+76" swimtime="00:01:10.68" resultid="2794" heatid="7895" lane="1" entrytime="00:01:11.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="792" reactiontime="+76" swimtime="00:00:27.16" resultid="2795" heatid="7923" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="1591" points="882" reactiontime="+72" swimtime="00:00:59.02" resultid="2796" heatid="8002" lane="5" entrytime="00:01:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="766" reactiontime="+72" swimtime="00:00:32.23" resultid="2797" heatid="8046" lane="8" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzimierz" gender="M" lastname="Jarzyna" nation="POL" athleteid="2807">
              <RESULTS>
                <RESULT eventid="1076" points="568" reactiontime="+94" swimtime="00:00:32.59" resultid="2808" heatid="7690" lane="5" entrytime="00:00:33.69" />
                <RESULT eventid="1108" points="581" reactiontime="+94" swimtime="00:03:16.76" resultid="2809" heatid="7722" lane="6" entrytime="00:03:31.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.12" />
                    <SPLIT distance="100" swimtime="00:01:36.44" />
                    <SPLIT distance="150" swimtime="00:02:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="508" reactiontime="+78" swimtime="00:00:41.54" resultid="2810" heatid="7767" lane="3" entrytime="00:00:44.21" />
                <RESULT eventid="1286" points="527" reactiontime="+93" swimtime="00:01:29.65" resultid="2811" heatid="7842" lane="8" entrytime="00:01:33.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="518" reactiontime="+79" swimtime="00:01:30.50" resultid="2812" heatid="7936" lane="8" entrytime="00:01:33.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="548" reactiontime="+90" swimtime="00:07:06.05" resultid="2813" heatid="8810" lane="1" entrytime="00:07:27.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.57" />
                    <SPLIT distance="100" swimtime="00:01:47.95" />
                    <SPLIT distance="150" swimtime="00:02:44.13" />
                    <SPLIT distance="200" swimtime="00:03:36.42" />
                    <SPLIT distance="250" swimtime="00:04:36.62" />
                    <SPLIT distance="300" swimtime="00:05:36.15" />
                    <SPLIT distance="350" swimtime="00:06:24.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="582" reactiontime="+84" swimtime="00:03:18.15" resultid="2814" heatid="8013" lane="7" entrytime="00:03:26.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                    <SPLIT distance="100" swimtime="00:02:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="529" reactiontime="+96" swimtime="00:06:11.93" resultid="2815" heatid="9068" lane="1" entrytime="00:06:39.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:28.64" />
                    <SPLIT distance="150" swimtime="00:02:17.30" />
                    <SPLIT distance="200" swimtime="00:03:06.60" />
                    <SPLIT distance="250" swimtime="00:03:54.35" />
                    <SPLIT distance="300" swimtime="00:04:42.21" />
                    <SPLIT distance="350" swimtime="00:05:28.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="2825">
              <RESULTS>
                <RESULT eventid="1076" points="604" reactiontime="+94" swimtime="00:00:30.05" resultid="2826" heatid="7696" lane="3" entrytime="00:00:30.61" />
                <RESULT eventid="1108" points="623" reactiontime="+89" swimtime="00:02:47.30" resultid="2827" heatid="7727" lane="7" entrytime="00:02:53.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                    <SPLIT distance="150" swimtime="00:02:09.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="617" reactiontime="+86" swimtime="00:01:06.28" resultid="2828" heatid="7815" lane="6" entrytime="00:01:07.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="490" reactiontime="+93" swimtime="00:03:01.64" resultid="2829" heatid="7862" lane="5" entrytime="00:03:10.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                    <SPLIT distance="100" swimtime="00:01:25.93" />
                    <SPLIT distance="150" swimtime="00:02:14.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="2830" heatid="7960" lane="2" entrytime="00:02:33.21" />
                <RESULT comment="K16 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu  (Czas: 21:40)" eventid="1543" reactiontime="+94" status="DSQ" swimtime="00:06:00.73" resultid="2831" heatid="8808" lane="7" entrytime="00:06:12.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:11.59" />
                    <SPLIT distance="200" swimtime="00:02:56.66" />
                    <SPLIT distance="250" swimtime="00:03:48.73" />
                    <SPLIT distance="300" swimtime="00:04:40.26" />
                    <SPLIT distance="350" swimtime="00:05:21.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="447" reactiontime="+90" swimtime="00:01:21.67" resultid="2832" heatid="7995" lane="3" entrytime="00:01:30.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="618" reactiontime="+89" swimtime="00:02:50.15" resultid="2833" heatid="8016" lane="8" entrytime="00:02:52.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                    <SPLIT distance="100" swimtime="00:01:22.63" />
                    <SPLIT distance="150" swimtime="00:02:06.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="2834">
              <RESULTS>
                <RESULT eventid="1076" points="586" reactiontime="+75" swimtime="00:00:28.34" resultid="2835" heatid="7700" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1108" points="466" reactiontime="+81" swimtime="00:02:44.12" resultid="2836" heatid="7727" lane="3" entrytime="00:02:50.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                    <SPLIT distance="100" swimtime="00:01:18.29" />
                    <SPLIT distance="150" swimtime="00:02:04.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="529" reactiontime="+66" swimtime="00:00:33.54" resultid="2837" heatid="7773" lane="4" entrytime="00:00:33.85" />
                <RESULT eventid="1286" points="537" reactiontime="+86" swimtime="00:01:12.63" resultid="2838" heatid="7849" lane="1" entrytime="00:01:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="485" reactiontime="+81" swimtime="00:01:21.46" resultid="2839" heatid="7891" lane="1" entrytime="00:01:23.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="377" reactiontime="+89" swimtime="00:06:17.78" resultid="2840" heatid="8808" lane="6" entrytime="00:06:09.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="100" swimtime="00:01:28.02" />
                    <SPLIT distance="150" swimtime="00:02:15.75" />
                    <SPLIT distance="200" swimtime="00:03:03.62" />
                    <SPLIT distance="250" swimtime="00:03:55.00" />
                    <SPLIT distance="300" swimtime="00:04:47.74" />
                    <SPLIT distance="350" swimtime="00:05:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="2841" heatid="8016" lane="1" entrytime="00:02:51.50" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="2842" heatid="8042" lane="8" entrytime="00:00:36.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="2843">
              <RESULTS>
                <RESULT eventid="1059" points="526" reactiontime="+92" swimtime="00:00:34.40" resultid="2844" heatid="7678" lane="8" entrytime="00:00:35.01" />
                <RESULT eventid="1092" points="559" reactiontime="+99" swimtime="00:03:05.70" resultid="2845" heatid="7715" lane="3" entrytime="00:03:15.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:29.60" />
                    <SPLIT distance="150" swimtime="00:02:22.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="569" reactiontime="+91" swimtime="00:03:25.57" resultid="2846" heatid="7781" lane="3" entrytime="00:03:30.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                    <SPLIT distance="100" swimtime="00:01:38.74" />
                    <SPLIT distance="150" swimtime="00:02:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="547" reactiontime="+92" swimtime="00:01:26.26" resultid="2847" heatid="7832" lane="1" entrytime="00:01:28.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="544" reactiontime="+92" swimtime="00:01:36.62" resultid="2848" heatid="7878" lane="8" entrytime="00:01:38.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" status="WDR" swimtime="00:00:00.00" resultid="2849" entrytime="00:06:59.90" />
                <RESULT eventid="1574" points="430" reactiontime="+88" swimtime="00:01:30.12" resultid="2850" heatid="7989" lane="2" entrytime="00:01:32.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="532" reactiontime="+89" swimtime="00:00:43.71" resultid="2851" heatid="8025" lane="5" entrytime="00:00:45.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-12" firstname="Adam" gender="M" lastname="Przybylski" nation="POL" athleteid="2852">
              <RESULTS>
                <RESULT eventid="1076" points="681" reactiontime="+81" swimtime="00:00:27.48" resultid="2853" heatid="7703" lane="1" entrytime="00:00:28.12" />
                <RESULT eventid="1190" points="551" reactiontime="+69" swimtime="00:00:34.95" resultid="2854" heatid="7769" lane="7" entrytime="00:00:40.12" />
                <RESULT eventid="1254" points="615" reactiontime="+79" swimtime="00:01:02.22" resultid="2855" heatid="7819" lane="5" entrytime="00:01:02.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="597" reactiontime="+78" swimtime="00:00:31.39" resultid="2856" heatid="7910" lane="3" entrytime="00:00:38.12" />
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="2857" heatid="7939" lane="1" entrytime="00:01:16.12" />
                <RESULT eventid="1591" points="462" reactiontime="+84" swimtime="00:01:16.03" resultid="2858" heatid="7995" lane="7" entrytime="00:01:35.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="518" reactiontime="+72" swimtime="00:02:49.65" resultid="2859" heatid="8016" lane="7" entrytime="00:02:49.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:20.17" />
                    <SPLIT distance="150" swimtime="00:02:05.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-15" firstname="Michał" gender="M" lastname="Skrok" nation="POL" athleteid="2860">
              <RESULTS>
                <RESULT eventid="1108" points="706" reactiontime="+76" swimtime="00:02:22.92" resultid="2861" heatid="7731" lane="2" entrytime="00:02:30.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:10.03" />
                    <SPLIT distance="150" swimtime="00:01:49.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="732" reactiontime="+78" swimtime="00:02:38.09" resultid="2862" heatid="7795" lane="1" entrytime="00:02:40.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:15.67" />
                    <SPLIT distance="150" swimtime="00:01:56.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="735" reactiontime="+72" swimtime="00:01:05.43" resultid="2863" heatid="7852" lane="4" entrytime="00:01:08.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="701" reactiontime="+76" swimtime="00:01:12.04" resultid="2864" heatid="7894" lane="4" entrytime="00:01:12.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="2865" heatid="8808" lane="2" entrytime="00:06:10.40" />
                <RESULT eventid="1623" points="622" reactiontime="+75" swimtime="00:02:32.23" resultid="2866" heatid="8018" lane="2" entrytime="00:02:35.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:15.06" />
                    <SPLIT distance="150" swimtime="00:01:54.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="716" reactiontime="+72" swimtime="00:00:32.27" resultid="2867" heatid="8046" lane="4" entrytime="00:00:32.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Paweł" gender="M" lastname="Cieśliński" nation="POL" athleteid="2868">
              <RESULTS>
                <RESULT eventid="1108" points="377" reactiontime="+100" swimtime="00:02:56.16" resultid="2869" heatid="7726" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:01:26.13" />
                    <SPLIT distance="150" swimtime="00:02:15.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="501" reactiontime="+93" swimtime="00:02:59.39" resultid="2870" heatid="7793" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:26.42" />
                    <SPLIT distance="150" swimtime="00:02:13.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="333" reactiontime="+93" swimtime="00:03:02.54" resultid="2871" heatid="7863" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                    <SPLIT distance="100" swimtime="00:01:28.53" />
                    <SPLIT distance="150" swimtime="00:02:17.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="468" reactiontime="+90" swimtime="00:01:22.42" resultid="2872" heatid="7892" lane="1" entrytime="00:01:21.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="WDR" swimtime="00:00:00.00" resultid="2873" entrytime="00:06:20.00" />
                <RESULT eventid="1591" points="306" reactiontime="+99" swimtime="00:01:24.34" resultid="2874" heatid="7997" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="438" reactiontime="+80" swimtime="00:00:37.99" resultid="2875" heatid="8040" lane="4" entrytime="00:00:37.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-04" firstname="Paweł" gender="M" lastname="Opaliński" nation="POL" athleteid="2876">
              <RESULTS>
                <RESULT eventid="1076" points="690" reactiontime="+79" swimtime="00:00:26.84" resultid="2877" heatid="7700" lane="4" entrytime="00:00:29.01" />
                <RESULT eventid="1222" points="642" reactiontime="+86" swimtime="00:02:45.16" resultid="2878" heatid="7795" lane="8" entrytime="00:02:41.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:02:01.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="624" reactiontime="+80" swimtime="00:01:00.18" resultid="2879" heatid="7822" lane="2" entrytime="00:00:59.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="653" reactiontime="+83" swimtime="00:01:13.77" resultid="2880" heatid="7894" lane="5" entrytime="00:01:13.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="572" reactiontime="+76" swimtime="00:02:14.22" resultid="2881" heatid="7965" lane="5" entrytime="00:02:12.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:04.33" />
                    <SPLIT distance="150" swimtime="00:01:39.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="616" reactiontime="+76" swimtime="00:00:33.93" resultid="2882" heatid="8045" lane="8" entrytime="00:00:34.02" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Motyl Senior MOSiR St. Wola C">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+88" swimtime="00:01:55.53" resultid="2884" heatid="7872" lane="5" entrytime="00:01:58.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:01.93" />
                    <SPLIT distance="150" swimtime="00:01:28.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2781" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="2860" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2789" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="2852" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" reactiontime="+89" swimtime="00:01:46.14" resultid="2887" heatid="7974" lane="6" entrytime="00:01:48.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                    <SPLIT distance="100" swimtime="00:00:53.40" />
                    <SPLIT distance="150" swimtime="00:01:20.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2781" number="1" />
                    <RELAYPOSITION athleteid="2876" number="2" />
                    <RELAYPOSITION athleteid="2852" number="3" />
                    <RELAYPOSITION athleteid="2789" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NARYD" nation="POL" region="11" clubid="6231" name="Naprzód Rydułtowy">
          <ATHLETES>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="6230">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="6232" heatid="7685" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1108" points="328" reactiontime="+99" swimtime="00:04:17.61" resultid="6233" heatid="7720" lane="3" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.08" />
                    <SPLIT distance="100" swimtime="00:02:05.27" />
                    <SPLIT distance="150" swimtime="00:03:17.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="6234" heatid="7764" lane="6" entrytime="00:00:55.00" />
                <RESULT eventid="1318" points="344" reactiontime="+86" swimtime="00:04:38.24" resultid="6235" heatid="7860" lane="2" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.53" />
                    <SPLIT distance="100" swimtime="00:02:11.12" />
                    <SPLIT distance="150" swimtime="00:03:23.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="217" reactiontime="+84" swimtime="00:02:04.85" resultid="6236" heatid="7934" lane="8" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.38" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z1 - Nieprawidłowa kolejność stylów pływania (prawidłowa: motylkowy, grzbietowy, klasyczny, dowolny)  (Czas: 22:17)" eventid="1543" reactiontime="+98" status="DSQ" swimtime="00:08:52.59" resultid="6237" heatid="8812" lane="5" entrytime="00:09:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.69" />
                    <SPLIT distance="100" swimtime="00:02:25.45" />
                    <SPLIT distance="150" swimtime="00:03:42.46" />
                    <SPLIT distance="200" swimtime="00:04:57.72" />
                    <SPLIT distance="250" swimtime="00:06:13.77" />
                    <SPLIT distance="300" swimtime="00:07:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="6238" heatid="7992" lane="3" entrytime="00:02:09.00" />
                <RESULT eventid="1623" points="309" reactiontime="+77" swimtime="00:04:28.85" resultid="6239" heatid="8010" lane="4" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.92" />
                    <SPLIT distance="100" swimtime="00:02:09.80" />
                    <SPLIT distance="150" swimtime="00:03:20.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZSTP" nation="RUS" clubid="2675" name="Nevskie Zvezdy St. Petersburg">
          <ATHLETES>
            <ATHLETE birthdate="1972-06-06" firstname="Marina" gender="F" lastname="Perepelkina" nation="RUS" athleteid="2676">
              <RESULTS>
                <RESULT eventid="1366" points="704" reactiontime="+85" swimtime="00:01:25.08" resultid="2677" heatid="7880" lane="6" entrytime="00:01:24.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="668" reactiontime="+87" swimtime="00:00:39.27" resultid="2679" heatid="8028" lane="2" entrytime="00:00:38.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-11-08" firstname="Igor" gender="M" lastname="Andreev" nation="RUS" athleteid="2678">
              <RESULTS>
                <RESULT eventid="1190" points="469" reactiontime="+80" swimtime="00:00:42.88" resultid="2680" heatid="7768" lane="8" entrytime="00:00:43.00" />
                <RESULT eventid="1415" points="604" reactiontime="+95" swimtime="00:00:36.15" resultid="2681" heatid="7911" lane="7" entrytime="00:00:37.20" />
                <RESULT eventid="1591" points="491" reactiontime="+99" swimtime="00:01:30.76" resultid="2682" heatid="7995" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-04-17" firstname="Alexander" gender="M" lastname="Kharchenko" nation="RUS" athleteid="2683">
              <RESULTS>
                <RESULT eventid="1108" points="606" reactiontime="+80" swimtime="00:03:11.00" resultid="2684" heatid="7723" lane="5" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:30.19" />
                    <SPLIT distance="150" swimtime="00:02:25.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="615" reactiontime="+89" swimtime="00:03:34.18" resultid="2685" heatid="7791" lane="8" entrytime="00:03:19.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                    <SPLIT distance="100" swimtime="00:01:40.76" />
                    <SPLIT distance="150" swimtime="00:02:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="677" reactiontime="+86" swimtime="00:01:30.40" resultid="2686" heatid="7888" lane="5" entrytime="00:01:28.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="721" reactiontime="+82" swimtime="00:00:39.40" resultid="2687" heatid="8039" lane="7" entrytime="00:00:38.79" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-10-19" firstname="Igor" gender="M" lastname="Lukonenko" nation="RUS" athleteid="2688">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="2689" heatid="7732" lane="7" entrytime="00:02:25.00" />
                <RESULT eventid="1190" points="632" reactiontime="+77" swimtime="00:00:34.23" resultid="2690" heatid="7771" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1415" points="693" reactiontime="+92" swimtime="00:00:31.12" resultid="2691" heatid="7916" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="1655" points="597" reactiontime="+97" swimtime="00:00:37.26" resultid="2692" heatid="8040" lane="8" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-10-06" firstname="Sergey" gender="M" lastname="Frolov" nation="RUS" athleteid="2693">
              <RESULTS>
                <RESULT eventid="1156" points="508" swimtime="00:20:38.61" resultid="2694" heatid="8718" lane="7" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                    <SPLIT distance="200" swimtime="00:02:38.84" />
                    <SPLIT distance="400" swimtime="00:05:24.78" />
                    <SPLIT distance="500" swimtime="00:06:48.07" />
                    <SPLIT distance="600" swimtime="00:08:11.77" />
                    <SPLIT distance="700" swimtime="00:09:36.24" />
                    <SPLIT distance="800" swimtime="00:11:01.44" />
                    <SPLIT distance="900" swimtime="00:12:25.51" />
                    <SPLIT distance="1000" swimtime="00:13:48.58" />
                    <SPLIT distance="1100" swimtime="00:15:11.84" />
                    <SPLIT distance="1200" swimtime="00:16:34.53" />
                    <SPLIT distance="1300" swimtime="00:17:56.66" />
                    <SPLIT distance="1400" swimtime="00:19:19.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="503" reactiontime="+89" swimtime="00:02:24.17" resultid="2695" heatid="7964" lane="2" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                    <SPLIT distance="150" swimtime="00:01:45.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="504" reactiontime="+85" swimtime="00:05:08.82" resultid="2696" heatid="9060" lane="1" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:12.84" />
                    <SPLIT distance="150" swimtime="00:01:52.30" />
                    <SPLIT distance="200" swimtime="00:02:32.09" />
                    <SPLIT distance="300" swimtime="00:03:50.98" />
                    <SPLIT distance="350" swimtime="00:04:30.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZWAR" nation="POL" region="14" clubid="6116" name="Niezrzeszeni.pl ">
          <CONTACT city="Warszawa" email="niezrzeszenipl@gmail.com" internet="niezrzeszeni.pl" name="Wawer" phone="505960036" state="MAZOW" street="Tołstoja 1 m 407" zip="01-910" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="6117">
              <RESULTS>
                <RESULT eventid="1156" points="389" swimtime="00:26:27.21" resultid="6118" heatid="8723" lane="4" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:32.45" />
                    <SPLIT distance="200" swimtime="00:03:15.26" />
                    <SPLIT distance="300" swimtime="00:05:00.15" />
                    <SPLIT distance="400" swimtime="00:06:46.88" />
                    <SPLIT distance="500" swimtime="00:08:33.74" />
                    <SPLIT distance="600" swimtime="00:10:21.45" />
                    <SPLIT distance="700" swimtime="00:12:10.27" />
                    <SPLIT distance="800" swimtime="00:13:58.19" />
                    <SPLIT distance="900" swimtime="00:15:45.36" />
                    <SPLIT distance="1000" swimtime="00:17:33.38" />
                    <SPLIT distance="1100" swimtime="00:19:21.24" />
                    <SPLIT distance="1200" swimtime="00:21:09.02" />
                    <SPLIT distance="1300" swimtime="00:22:56.21" />
                    <SPLIT distance="1400" swimtime="00:24:45.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="384" reactiontime="+114" swimtime="00:03:43.56" resultid="6119" heatid="7787" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.79" />
                    <SPLIT distance="100" swimtime="00:01:45.37" />
                    <SPLIT distance="150" swimtime="00:02:44.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="320" reactiontime="+106" swimtime="00:01:24.77" resultid="6120" heatid="7808" lane="2" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="368" reactiontime="+111" swimtime="00:03:06.07" resultid="6121" heatid="7954" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                    <SPLIT distance="100" swimtime="00:01:28.82" />
                    <SPLIT distance="150" swimtime="00:02:17.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="WDR" swimtime="00:00:00.00" resultid="6122" />
                <RESULT eventid="1655" points="291" reactiontime="+110" swimtime="00:00:46.01" resultid="6123" heatid="8032" lane="2" entrytime="00:00:46.00" />
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="6124" heatid="9068" lane="3" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-08-26" firstname="Małgorzata" gender="F" lastname="Piechura" nation="POL" athleteid="6125">
              <RESULTS>
                <RESULT eventid="1059" points="238" reactiontime="+106" swimtime="00:00:43.84" resultid="6126" heatid="7673" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1206" points="358" reactiontime="+120" swimtime="00:03:53.90" resultid="6127" heatid="7778" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.68" />
                    <SPLIT distance="100" swimtime="00:01:54.63" />
                    <SPLIT distance="150" swimtime="00:02:54.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="207" reactiontime="+117" swimtime="00:01:55.04" resultid="6128" heatid="7826" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="133" reactiontime="+113" swimtime="00:00:58.47" resultid="6129" heatid="7897" lane="5" />
                <RESULT eventid="1463" points="190" reactiontime="+117" swimtime="00:03:46.41" resultid="6130" heatid="7945" lane="7" entrytime="00:03:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.17" />
                    <SPLIT distance="100" swimtime="00:01:46.19" />
                    <SPLIT distance="150" swimtime="00:02:45.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="194" reactiontime="+115" swimtime="00:07:57.93" resultid="6131" heatid="9052" lane="2" entrytime="00:07:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.40" />
                    <SPLIT distance="100" swimtime="00:01:47.96" />
                    <SPLIT distance="150" swimtime="00:02:48.68" />
                    <SPLIT distance="200" swimtime="00:03:48.96" />
                    <SPLIT distance="250" swimtime="00:05:56.47" />
                    <SPLIT distance="300" swimtime="00:06:59.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OROPO" nation="POL" region="07" clubid="3639" name="Odrzańskie Ratownictwo Spec. Opole" shortname="ORS Opole">
          <CONTACT email="wkania62@gmail.com" name="Kania Waldemar" />
          <ATHLETES>
            <ATHLETE birthdate="1973-01-01" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="3640">
              <RESULTS>
                <RESULT eventid="1173" points="525" reactiontime="+71" swimtime="00:00:39.20" resultid="3641" heatid="7758" lane="1" entrytime="00:00:40.01" />
                <RESULT eventid="1270" points="535" reactiontime="+101" swimtime="00:01:23.90" resultid="3642" heatid="7833" lane="1" entrytime="00:01:25.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="497" reactiontime="+82" swimtime="00:01:25.78" resultid="3643" heatid="7929" lane="3" entrytime="00:01:26.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="551" reactiontime="+75" swimtime="00:03:02.19" resultid="3644" heatid="8008" lane="8" entrytime="00:03:03.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:27.74" />
                    <SPLIT distance="150" swimtime="00:02:15.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="439" reactiontime="+105" swimtime="00:06:04.12" resultid="3645" heatid="9049" lane="5" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:08.24" />
                    <SPLIT distance="200" swimtime="00:02:55.66" />
                    <SPLIT distance="250" swimtime="00:03:43.21" />
                    <SPLIT distance="300" swimtime="00:04:30.50" />
                    <SPLIT distance="350" swimtime="00:05:18.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Waldemar" gender="M" lastname="Kania" nation="POL" athleteid="3646">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3647" heatid="7695" lane="2" entrytime="00:00:31.01" />
                <RESULT eventid="1156" points="532" swimtime="00:21:57.96" resultid="3648" heatid="8719" lane="7" entrytime="00:21:59.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:21.46" />
                    <SPLIT distance="200" swimtime="00:02:50.65" />
                    <SPLIT distance="300" swimtime="00:04:20.01" />
                    <SPLIT distance="400" swimtime="00:05:48.88" />
                    <SPLIT distance="500" swimtime="00:07:17.33" />
                    <SPLIT distance="600" swimtime="00:08:45.25" />
                    <SPLIT distance="700" swimtime="00:10:12.99" />
                    <SPLIT distance="800" swimtime="00:11:41.49" />
                    <SPLIT distance="900" swimtime="00:13:10.23" />
                    <SPLIT distance="1000" swimtime="00:14:39.69" />
                    <SPLIT distance="1100" swimtime="00:16:09.56" />
                    <SPLIT distance="1200" swimtime="00:17:38.16" />
                    <SPLIT distance="1300" swimtime="00:19:07.12" />
                    <SPLIT distance="1400" swimtime="00:20:34.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="508" reactiontime="+89" swimtime="00:01:10.71" resultid="3649" heatid="7813" lane="2" entrytime="00:01:10.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="525" reactiontime="+88" swimtime="00:02:35.88" resultid="3650" heatid="7960" lane="7" entrytime="00:02:34.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:15.30" />
                    <SPLIT distance="150" swimtime="00:01:56.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="3651" heatid="8013" lane="2" entrytime="00:03:24.01" />
                <RESULT eventid="1703" points="520" reactiontime="+92" swimtime="00:05:31.18" resultid="3652" heatid="9064" lane="7" entrytime="00:05:30.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="100" swimtime="00:01:18.20" />
                    <SPLIT distance="150" swimtime="00:02:00.71" />
                    <SPLIT distance="200" swimtime="00:02:43.49" />
                    <SPLIT distance="250" swimtime="00:03:25.72" />
                    <SPLIT distance="300" swimtime="00:04:08.02" />
                    <SPLIT distance="350" swimtime="00:04:50.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Grzegorz" gender="M" lastname="Stanek" nation="POL" athleteid="3653">
              <RESULTS>
                <RESULT eventid="1108" points="884" reactiontime="+77" swimtime="00:02:22.34" resultid="3654" heatid="7732" lane="6" entrytime="00:02:24.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:05.30" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="832" reactiontime="+76" swimtime="00:01:04.31" resultid="3655" heatid="7854" lane="5" entrytime="00:01:06.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="975" reactiontime="+82" swimtime="00:05:06.71" resultid="3656" heatid="8806" lane="6" entrytime="00:05:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:09.70" />
                    <SPLIT distance="150" swimtime="00:01:49.79" />
                    <SPLIT distance="200" swimtime="00:02:29.14" />
                    <SPLIT distance="250" swimtime="00:03:12.68" />
                    <SPLIT distance="300" swimtime="00:03:56.95" />
                    <SPLIT distance="350" swimtime="00:04:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="679" reactiontime="+80" swimtime="00:04:39.71" resultid="3657" heatid="9060" lane="4" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:08.20" />
                    <SPLIT distance="150" swimtime="00:01:43.94" />
                    <SPLIT distance="200" swimtime="00:02:19.65" />
                    <SPLIT distance="250" swimtime="00:02:55.17" />
                    <SPLIT distance="300" swimtime="00:03:30.26" />
                    <SPLIT distance="350" swimtime="00:04:05.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Wojciech" gender="M" lastname="Stanek" nation="POL" athleteid="3658">
              <RESULTS>
                <RESULT eventid="1108" points="516" reactiontime="+80" swimtime="00:02:38.32" resultid="3659" heatid="7728" lane="6" entrytime="00:02:46.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:17.37" />
                    <SPLIT distance="150" swimtime="00:02:01.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="448" reactiontime="+84" swimtime="00:01:15.04" resultid="3660" heatid="7847" lane="8" entrytime="00:01:17.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="448" reactiontime="+86" swimtime="00:05:50.61" resultid="3661" heatid="8807" lane="2" entrytime="00:05:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:19.35" />
                    <SPLIT distance="150" swimtime="00:02:10.26" />
                    <SPLIT distance="200" swimtime="00:02:56.79" />
                    <SPLIT distance="250" swimtime="00:03:44.40" />
                    <SPLIT distance="300" swimtime="00:04:32.53" />
                    <SPLIT distance="350" swimtime="00:05:12.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="496" reactiontime="+75" swimtime="00:05:10.03" resultid="3662" heatid="9063" lane="5" entrytime="00:05:19.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                    <SPLIT distance="100" swimtime="00:01:14.08" />
                    <SPLIT distance="150" swimtime="00:01:52.67" />
                    <SPLIT distance="200" swimtime="00:02:32.73" />
                    <SPLIT distance="250" swimtime="00:03:12.06" />
                    <SPLIT distance="300" swimtime="00:03:51.38" />
                    <SPLIT distance="350" swimtime="00:04:30.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Marcin" gender="M" lastname="Wilczyński" nation="POL" athleteid="3663">
              <RESULTS>
                <RESULT eventid="1222" points="664" reactiontime="+95" swimtime="00:02:43.72" resultid="3664" heatid="7794" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:18.79" />
                    <SPLIT distance="150" swimtime="00:02:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="683" reactiontime="+93" swimtime="00:01:14.49" resultid="3665" heatid="7894" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="WDR" swimtime="00:00:00.00" resultid="3666" entrytime="00:05:33.00" />
                <RESULT eventid="1655" points="651" reactiontime="+86" swimtime="00:00:34.02" resultid="3667" heatid="8045" lane="7" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OMTPO" nation="POL" region="15" clubid="6171" name="One Man Team Poznań">
          <CONTACT city="Poznań" email="gmo@o2.pl" name="Monczak" phone="608639696" state="WLKP" zip="61-160" />
          <ATHLETES>
            <ATHLETE birthdate="1973-05-25" firstname="Grzegorz" gender="M" lastname="Monczak" nation="POL" athleteid="6172">
              <RESULTS>
                <RESULT eventid="1108" points="597" reactiontime="+76" swimtime="00:02:31.86" resultid="6173" heatid="7730" lane="6" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:13.54" />
                    <SPLIT distance="150" swimtime="00:01:58.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="714" reactiontime="+76" swimtime="00:18:35.11" resultid="6174" heatid="8717" lane="2" entrytime="00:18:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:09.27" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                    <SPLIT distance="200" swimtime="00:02:22.89" />
                    <SPLIT distance="250" swimtime="00:03:00.30" />
                    <SPLIT distance="300" swimtime="00:03:37.38" />
                    <SPLIT distance="350" swimtime="00:04:14.51" />
                    <SPLIT distance="400" swimtime="00:04:51.73" />
                    <SPLIT distance="450" swimtime="00:05:29.50" />
                    <SPLIT distance="500" swimtime="00:06:07.00" />
                    <SPLIT distance="550" swimtime="00:06:44.94" />
                    <SPLIT distance="600" swimtime="00:07:22.82" />
                    <SPLIT distance="650" swimtime="00:07:59.98" />
                    <SPLIT distance="700" swimtime="00:08:37.56" />
                    <SPLIT distance="750" swimtime="00:09:15.02" />
                    <SPLIT distance="800" swimtime="00:09:52.30" />
                    <SPLIT distance="850" swimtime="00:10:29.48" />
                    <SPLIT distance="900" swimtime="00:11:06.83" />
                    <SPLIT distance="950" swimtime="00:11:44.54" />
                    <SPLIT distance="1000" swimtime="00:12:21.72" />
                    <SPLIT distance="1050" swimtime="00:12:59.10" />
                    <SPLIT distance="1100" swimtime="00:13:36.46" />
                    <SPLIT distance="1150" swimtime="00:14:14.01" />
                    <SPLIT distance="1200" swimtime="00:14:51.12" />
                    <SPLIT distance="1250" swimtime="00:15:28.22" />
                    <SPLIT distance="1300" swimtime="00:16:05.44" />
                    <SPLIT distance="1350" swimtime="00:16:42.95" />
                    <SPLIT distance="1400" swimtime="00:17:20.55" />
                    <SPLIT distance="1450" swimtime="00:17:58.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="684" reactiontime="+69" swimtime="00:00:59.09" resultid="6175" heatid="7822" lane="3" entrytime="00:00:59.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="589" reactiontime="+74" swimtime="00:01:11.34" resultid="6176" heatid="7851" lane="1" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="486" reactiontime="+77" swimtime="00:00:31.95" resultid="6177" heatid="7918" lane="7" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1479" points="644" reactiontime="+77" swimtime="00:02:10.84" resultid="6178" heatid="7966" lane="7" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:05.32" />
                    <SPLIT distance="150" swimtime="00:01:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="6179" heatid="7999" lane="1" entrytime="00:01:12.00" entrycourse="SCM" />
                <RESULT eventid="1703" points="653" reactiontime="+79" swimtime="00:04:37.30" resultid="6180" heatid="9059" lane="1" entrytime="00:04:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:42.58" />
                    <SPLIT distance="200" swimtime="00:02:17.86" />
                    <SPLIT distance="250" swimtime="00:02:53.42" />
                    <SPLIT distance="300" swimtime="00:03:28.96" />
                    <SPLIT distance="350" swimtime="00:04:04.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORRAD" nation="POL" region="11" clubid="3444" name="Orka Masters Radlin">
          <CONTACT email="otelom.080966@interia.pl" name="OTLIK Marian" zip="44-314" />
          <ATHLETES>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="3445">
              <RESULTS>
                <RESULT eventid="1108" points="553" reactiontime="+78" swimtime="00:03:20.00" resultid="3446" heatid="7723" lane="6" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:32.28" />
                    <SPLIT distance="150" swimtime="00:02:35.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="650" swimtime="00:24:40.50" resultid="3447" heatid="8722" lane="1" entrytime="00:26:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:27.84" />
                    <SPLIT distance="200" swimtime="00:03:05.02" />
                    <SPLIT distance="300" swimtime="00:04:44.90" />
                    <SPLIT distance="400" swimtime="00:06:25.03" />
                    <SPLIT distance="500" swimtime="00:08:05.35" />
                    <SPLIT distance="600" swimtime="00:09:45.30" />
                    <SPLIT distance="700" swimtime="00:11:24.61" />
                    <SPLIT distance="800" swimtime="00:13:04.41" />
                    <SPLIT distance="900" swimtime="00:14:44.73" />
                    <SPLIT distance="1000" swimtime="00:16:25.31" />
                    <SPLIT distance="1100" swimtime="00:18:05.93" />
                    <SPLIT distance="1200" swimtime="00:19:46.97" />
                    <SPLIT distance="1300" swimtime="00:21:23.67" />
                    <SPLIT distance="1400" swimtime="00:23:04.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="534" reactiontime="+79" swimtime="00:00:40.85" resultid="3448" heatid="7769" lane="8" entrytime="00:00:41.00" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="3449" heatid="7843" lane="8" entrytime="00:01:29.00" />
                <RESULT eventid="1479" points="506" reactiontime="+83" swimtime="00:02:52.91" resultid="3450" heatid="7956" lane="2" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:21.42" />
                    <SPLIT distance="150" swimtime="00:02:07.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="546" reactiontime="+92" swimtime="00:07:06.57" resultid="3451" heatid="8810" lane="2" entrytime="00:07:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.33" />
                    <SPLIT distance="100" swimtime="00:01:41.71" />
                    <SPLIT distance="150" swimtime="00:02:35.27" />
                    <SPLIT distance="200" swimtime="00:03:28.82" />
                    <SPLIT distance="250" swimtime="00:04:32.49" />
                    <SPLIT distance="300" swimtime="00:05:34.88" />
                    <SPLIT distance="350" swimtime="00:06:21.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="588" reactiontime="+79" swimtime="00:03:17.48" resultid="3452" heatid="8013" lane="6" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                    <SPLIT distance="100" swimtime="00:01:34.24" />
                    <SPLIT distance="150" swimtime="00:02:27.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="529" reactiontime="+91" swimtime="00:06:11.95" resultid="3453" heatid="9067" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:24.50" />
                    <SPLIT distance="150" swimtime="00:02:12.59" />
                    <SPLIT distance="200" swimtime="00:03:00.72" />
                    <SPLIT distance="250" swimtime="00:03:48.43" />
                    <SPLIT distance="300" swimtime="00:04:36.95" />
                    <SPLIT distance="350" swimtime="00:05:25.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-08-07" firstname="Leon" gender="M" lastname="Irczyk" nation="POL" athleteid="3454">
              <RESULTS>
                <RESULT eventid="1108" points="292" reactiontime="+115" swimtime="00:04:07.40" resultid="3455" heatid="7722" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.47" />
                    <SPLIT distance="100" swimtime="00:02:06.72" />
                    <SPLIT distance="150" swimtime="00:03:08.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="307" swimtime="00:31:39.94" resultid="3456" heatid="8725" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.40" />
                    <SPLIT distance="100" swimtime="00:01:50.43" />
                    <SPLIT distance="200" swimtime="00:03:57.46" />
                    <SPLIT distance="300" swimtime="00:06:03.95" />
                    <SPLIT distance="400" swimtime="00:08:15.00" />
                    <SPLIT distance="500" swimtime="00:10:22.84" />
                    <SPLIT distance="600" swimtime="00:12:30.97" />
                    <SPLIT distance="700" swimtime="00:14:40.90" />
                    <SPLIT distance="800" swimtime="00:16:49.93" />
                    <SPLIT distance="900" swimtime="00:19:00.61" />
                    <SPLIT distance="1000" swimtime="00:21:08.82" />
                    <SPLIT distance="1100" swimtime="00:23:18.62" />
                    <SPLIT distance="1200" swimtime="00:25:24.10" />
                    <SPLIT distance="1300" swimtime="00:27:30.75" />
                    <SPLIT distance="1400" swimtime="00:29:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="449" reactiontime="+125" swimtime="00:03:48.39" resultid="3457" heatid="7786" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.04" />
                    <SPLIT distance="100" swimtime="00:01:50.42" />
                    <SPLIT distance="150" swimtime="00:02:49.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="168" reactiontime="+109" swimtime="00:04:49.11" resultid="3458" heatid="7859" lane="5" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.76" />
                    <SPLIT distance="100" swimtime="00:02:10.99" />
                    <SPLIT distance="150" swimtime="00:03:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="417" reactiontime="+107" swimtime="00:01:44.59" resultid="3459" heatid="7883" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="284" reactiontime="+127" swimtime="00:08:50.72" resultid="3460" heatid="8812" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.60" />
                    <SPLIT distance="100" swimtime="00:02:07.07" />
                    <SPLIT distance="150" swimtime="00:03:27.02" />
                    <SPLIT distance="200" swimtime="00:04:41.41" />
                    <SPLIT distance="250" swimtime="00:05:44.69" />
                    <SPLIT distance="300" swimtime="00:06:46.53" />
                    <SPLIT distance="350" swimtime="00:07:50.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="343" reactiontime="+114" swimtime="00:00:48.30" resultid="3461" heatid="8031" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1703" points="246" reactiontime="+118" swimtime="00:07:59.88" resultid="3462" heatid="9070" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.91" />
                    <SPLIT distance="100" swimtime="00:01:49.35" />
                    <SPLIT distance="150" swimtime="00:02:49.42" />
                    <SPLIT distance="200" swimtime="00:03:51.22" />
                    <SPLIT distance="250" swimtime="00:04:54.10" />
                    <SPLIT distance="300" swimtime="00:05:57.23" />
                    <SPLIT distance="350" swimtime="00:07:00.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-07-08" firstname="Sławomir" gender="M" lastname="Szurek" nation="POL" athleteid="3463">
              <RESULTS>
                <RESULT eventid="1108" points="350" reactiontime="+85" swimtime="00:03:01.30" resultid="3464" heatid="7725" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="100" swimtime="00:01:24.54" />
                    <SPLIT distance="150" swimtime="00:02:18.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="359" swimtime="00:23:22.53" resultid="3465" heatid="8722" lane="3" entrytime="00:25:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:24.03" />
                    <SPLIT distance="200" swimtime="00:02:56.09" />
                    <SPLIT distance="300" swimtime="00:04:29.81" />
                    <SPLIT distance="400" swimtime="00:06:02.49" />
                    <SPLIT distance="500" swimtime="00:07:35.83" />
                    <SPLIT distance="600" swimtime="00:09:10.26" />
                    <SPLIT distance="700" swimtime="00:10:45.26" />
                    <SPLIT distance="800" swimtime="00:12:20.71" />
                    <SPLIT distance="900" swimtime="00:13:56.13" />
                    <SPLIT distance="1000" swimtime="00:15:31.54" />
                    <SPLIT distance="1100" swimtime="00:17:06.07" />
                    <SPLIT distance="1200" swimtime="00:18:41.15" />
                    <SPLIT distance="1300" swimtime="00:20:16.41" />
                    <SPLIT distance="1400" swimtime="00:21:51.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="388" reactiontime="+82" swimtime="00:01:11.37" resultid="3466" heatid="7811" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="353" reactiontime="+86" swimtime="00:01:24.61" resultid="3467" heatid="7843" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="350" reactiontime="+84" swimtime="00:00:35.64" resultid="3468" heatid="7913" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1479" points="347" reactiontime="+83" swimtime="00:02:40.75" resultid="3469" heatid="7956" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:17.89" />
                    <SPLIT distance="150" swimtime="00:02:00.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-09" firstname="Tomasz" gender="M" lastname="Żurczak" nation="POL" athleteid="3470">
              <RESULTS>
                <RESULT eventid="1156" points="359" swimtime="00:23:22.57" resultid="3471" heatid="8724" lane="6" entrytime="00:30:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                    <SPLIT distance="100" swimtime="00:01:22.66" />
                    <SPLIT distance="200" swimtime="00:02:55.28" />
                    <SPLIT distance="300" swimtime="00:04:28.63" />
                    <SPLIT distance="400" swimtime="00:06:02.15" />
                    <SPLIT distance="500" swimtime="00:07:36.77" />
                    <SPLIT distance="600" swimtime="00:09:11.26" />
                    <SPLIT distance="700" swimtime="00:10:45.45" />
                    <SPLIT distance="800" swimtime="00:12:19.93" />
                    <SPLIT distance="900" swimtime="00:13:54.72" />
                    <SPLIT distance="1000" swimtime="00:15:37.32" />
                    <SPLIT distance="1100" swimtime="00:17:03.86" />
                    <SPLIT distance="1200" swimtime="00:18:39.17" />
                    <SPLIT distance="1300" swimtime="00:20:14.81" />
                    <SPLIT distance="1400" swimtime="00:21:48.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="324" reactiontime="+94" swimtime="00:03:27.85" resultid="3472" heatid="7788" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.99" />
                    <SPLIT distance="100" swimtime="00:01:38.38" />
                    <SPLIT distance="150" swimtime="00:02:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="247" reactiontime="+97" swimtime="00:01:35.25" resultid="3473" heatid="7841" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="359" reactiontime="+100" swimtime="00:01:32.31" resultid="3474" heatid="7884" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="285" reactiontime="+104" swimtime="00:02:51.60" resultid="3475" heatid="7955" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:02:06.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-08" firstname="Marian" gender="M" lastname="Otlik" nation="POL" athleteid="3476">
              <RESULTS>
                <RESULT eventid="1076" status="WDR" swimtime="00:00:00.00" resultid="3477" heatid="7697" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="3478" heatid="7724" lane="3" entrytime="00:03:15.00" />
                <RESULT eventid="1254" status="WDR" swimtime="00:00:00.00" resultid="3479" heatid="7813" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="1286" status="WDR" swimtime="00:00:00.00" resultid="3480" heatid="7844" lane="3" entrytime="00:01:25.00" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="3481" heatid="7884" lane="6" entrytime="00:01:40.00" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="3482" heatid="7956" lane="1" entrytime="00:03:00.00" />
                <RESULT eventid="1655" status="WDR" swimtime="00:00:00.00" resultid="3483" heatid="8037" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="3484" entrytime="00:06:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-08-06" firstname="Renata" gender="F" lastname="Macionczyk" nation="POL" athleteid="3485">
              <RESULTS>
                <RESULT eventid="1059" points="418" reactiontime="+87" swimtime="00:00:36.31" resultid="3486" heatid="7676" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1206" points="339" reactiontime="+88" swimtime="00:03:53.25" resultid="3487" heatid="7780" lane="7" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.93" />
                    <SPLIT distance="100" swimtime="00:01:53.76" />
                    <SPLIT distance="150" swimtime="00:02:54.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="299" reactiontime="+90" swimtime="00:01:26.35" resultid="3488" heatid="7799" lane="7" entrytime="00:01:29.00" />
                <RESULT eventid="1366" points="303" reactiontime="+90" swimtime="00:01:49.91" resultid="3489" heatid="7876" lane="7" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" status="DNS" swimtime="00:00:00.00" resultid="3490" heatid="7946" lane="6" entrytime="00:03:20.00" />
                <RESULT eventid="1639" points="351" reactiontime="+87" swimtime="00:00:48.00" resultid="3491" heatid="8024" lane="7" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-08-30" firstname="Monika" gender="F" lastname="Rek-Dylich" nation="POL" athleteid="3492">
              <RESULTS>
                <RESULT eventid="1059" points="441" reactiontime="+90" swimtime="00:00:34.34" resultid="3493" heatid="7680" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1173" points="340" reactiontime="+76" swimtime="00:00:43.47" resultid="3494" heatid="7756" lane="3" entrytime="00:00:44.00" />
                <RESULT eventid="1238" points="350" reactiontime="+101" swimtime="00:01:21.53" resultid="3495" heatid="7800" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-24" firstname="Piotr" gender="M" lastname="Sobik" nation="POL" athleteid="3496">
              <RESULTS>
                <RESULT eventid="1318" status="WDR" swimtime="00:00:00.00" resultid="3497" heatid="7862" lane="1" entrytime="00:03:30.00" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="3498" heatid="7915" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1591" status="WDR" swimtime="00:00:00.00" resultid="3499" heatid="7996" lane="3" entrytime="00:01:23.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Orka Masters Radlin D">
              <RESULTS>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="3500" heatid="7970" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3463" number="1" />
                    <RELAYPOSITION athleteid="3454" number="2" />
                    <RELAYPOSITION athleteid="3445" number="3" />
                    <RELAYPOSITION athleteid="3470" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1357" reactiontime="+80" swimtime="00:02:38.51" resultid="3501" heatid="7868" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                    <SPLIT distance="100" swimtime="00:01:23.88" />
                    <SPLIT distance="150" swimtime="00:01:59.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3445" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3470" number="2" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3463" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3454" number="4" reactiontime="+80" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Orka Masters Radlin B">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+92" swimtime="00:02:17.79" resultid="3502" heatid="7734" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="150" swimtime="00:01:46.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3470" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="3485" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3492" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3463" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KIPRI" nation="LAT" clubid="2220" name="PK Kipsala Riga">
          <ATHLETES>
            <ATHLETE birthdate="1974-01-01" firstname="Galina" gender="F" lastname="Shikina" nation="LAT" athleteid="2227">
              <RESULTS>
                <RESULT eventid="1059" points="541" reactiontime="+113" swimtime="00:00:33.33" resultid="2228" heatid="7679" lane="6" entrytime="00:00:33.97" />
                <RESULT eventid="1173" points="552" reactiontime="+84" swimtime="00:00:38.87" resultid="2229" heatid="7757" lane="4" entrytime="00:00:40.43" />
                <RESULT eventid="1238" points="487" reactiontime="+82" swimtime="00:01:13.45" resultid="2230" heatid="7802" lane="1" entrytime="00:01:15.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="468" reactiontime="+78" swimtime="00:05:51.62" resultid="2231" heatid="9049" lane="1" entrytime="00:05:53.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:21.01" />
                    <SPLIT distance="150" swimtime="00:02:05.35" />
                    <SPLIT distance="200" swimtime="00:02:50.61" />
                    <SPLIT distance="250" swimtime="00:03:37.62" />
                    <SPLIT distance="300" swimtime="00:04:23.87" />
                    <SPLIT distance="350" swimtime="00:05:09.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Vyacheslav" gender="M" lastname="Shikin" nation="LAT" athleteid="2232">
              <RESULTS>
                <RESULT eventid="1076" points="372" reactiontime="+84" swimtime="00:00:33.03" resultid="2233" heatid="7692" lane="7" entrytime="00:00:32.54" />
                <RESULT eventid="1254" points="287" reactiontime="+83" swimtime="00:01:18.93" resultid="2234" heatid="7810" lane="3" entrytime="00:01:17.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PKOGR" nation="LAT" clubid="2221" name="PK Ogre">
          <ATHLETES>
            <ATHLETE birthdate="1992-01-01" firstname="Leonid" gender="M" lastname="Belushko" nation="LAT" athleteid="2222">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2223" heatid="7705" lane="6" entrytime="00:00:27.68" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="2224" heatid="7820" lane="4" entrytime="00:01:01.32" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="2225" heatid="7920" lane="6" entrytime="00:00:29.78" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="2226" heatid="8000" lane="5" entrytime="00:01:09.21" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STRAL" nation="CZE" clubid="2019" name="PK Straz pod Ralskem" shortname="Straz pod Ralskem">
          <ATHLETES>
            <ATHLETE birthdate="1988-03-30" firstname="Jiri" gender="M" lastname="Janovsky" nation="CZE" athleteid="2020">
              <RESULTS>
                <RESULT eventid="1108" points="668" reactiontime="+77" swimtime="00:02:17.88" resultid="2021" heatid="7733" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="150" swimtime="00:01:45.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="685" reactiontime="+78" swimtime="00:02:36.95" resultid="2022" heatid="7795" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:56.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="668" reactiontime="+75" swimtime="00:01:03.14" resultid="2023" heatid="7855" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="685" reactiontime="+80" swimtime="00:01:10.35" resultid="2024" heatid="7895" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="681" reactiontime="+77" swimtime="00:00:32.12" resultid="2025" heatid="8046" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1703" points="763" reactiontime="+79" swimtime="00:04:27.48" resultid="2026" heatid="9059" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                    <SPLIT distance="100" swimtime="00:01:03.11" />
                    <SPLIT distance="150" swimtime="00:01:37.24" />
                    <SPLIT distance="200" swimtime="00:02:11.35" />
                    <SPLIT distance="250" swimtime="00:02:45.62" />
                    <SPLIT distance="300" swimtime="00:03:20.43" />
                    <SPLIT distance="350" swimtime="00:03:54.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-08-16" firstname="Jakub" gender="M" lastname="Lechner" nation="CZE" athleteid="2027">
              <RESULTS>
                <RESULT eventid="1076" points="572" reactiontime="+82" swimtime="00:00:27.50" resultid="2028" heatid="7705" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="1318" points="318" reactiontime="+95" swimtime="00:03:06.50" resultid="2029" heatid="7863" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:19.73" />
                    <SPLIT distance="150" swimtime="00:02:08.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="442" reactiontime="+84" swimtime="00:05:58.22" resultid="2030" heatid="8807" lane="3" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                    <SPLIT distance="150" swimtime="00:02:03.77" />
                    <SPLIT distance="200" swimtime="00:02:49.78" />
                    <SPLIT distance="250" swimtime="00:03:40.89" />
                    <SPLIT distance="300" swimtime="00:04:33.31" />
                    <SPLIT distance="350" swimtime="00:05:17.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="338" reactiontime="+83" swimtime="00:02:46.81" resultid="2031" heatid="8015" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:23.03" />
                    <SPLIT distance="150" swimtime="00:02:04.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-06" firstname="Jan" gender="M" lastname="Milda" nation="CZE" athleteid="2032">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2033" heatid="7711" lane="8" entrytime="00:00:26.00" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="2034" heatid="7823" lane="5" entrytime="00:00:58.00" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="2035" heatid="7921" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="2036" heatid="8045" lane="6" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-03-15" firstname="Jiri" gender="M" lastname="Janovsky " nameprefix="Jr." nation="CZE" athleteid="2037">
              <RESULTS>
                <RESULT eventid="1156" points="486" swimtime="00:20:56.60" resultid="2038" heatid="8719" lane="2" entrytime="00:21:41.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="200" swimtime="00:02:43.26" />
                    <SPLIT distance="300" swimtime="00:04:06.40" />
                    <SPLIT distance="400" swimtime="00:05:30.20" />
                    <SPLIT distance="500" swimtime="00:06:54.19" />
                    <SPLIT distance="600" swimtime="00:08:18.69" />
                    <SPLIT distance="700" swimtime="00:09:43.14" />
                    <SPLIT distance="800" swimtime="00:11:08.36" />
                    <SPLIT distance="900" swimtime="00:12:33.49" />
                    <SPLIT distance="1000" swimtime="00:13:57.95" />
                    <SPLIT distance="1100" swimtime="00:15:22.39" />
                    <SPLIT distance="1200" swimtime="00:16:46.77" />
                    <SPLIT distance="1300" swimtime="00:18:10.91" />
                    <SPLIT distance="1400" swimtime="00:19:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="487" reactiontime="+79" swimtime="00:00:36.42" resultid="2039" heatid="7771" lane="4" entrytime="00:00:35.10" />
                <RESULT eventid="1254" points="450" reactiontime="+97" swimtime="00:01:09.02" resultid="2040" heatid="7815" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="477" reactiontime="+98" swimtime="00:02:26.74" resultid="2041" heatid="7962" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:11.74" />
                    <SPLIT distance="150" swimtime="00:01:49.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="515" reactiontime="+95" swimtime="00:05:06.77" resultid="2042" heatid="9063" lane="3" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                    <SPLIT distance="150" swimtime="00:01:52.33" />
                    <SPLIT distance="200" swimtime="00:02:30.92" />
                    <SPLIT distance="250" swimtime="00:03:10.21" />
                    <SPLIT distance="300" swimtime="00:03:49.26" />
                    <SPLIT distance="350" swimtime="00:04:28.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Straz pod Ralskem B" number="1">
              <RESULTS>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="2043" heatid="7868" lane="7">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2037" number="1" />
                    <RELAYPOSITION athleteid="2020" number="2" />
                    <RELAYPOSITION athleteid="2027" number="3" />
                    <RELAYPOSITION athleteid="2032" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="UMBBB" nation="SVK" region="SSO" clubid="1919" name="PO KTV UMB Banska Bystrica">
          <ATHLETES>
            <ATHLETE birthdate="1963-04-17" firstname="Branislav" gender="M" lastname="Hakel" nation="SVK" license="15901" athleteid="1920">
              <RESULTS>
                <RESULT eventid="1286" points="846" reactiontime="+65" swimtime="00:01:09.24" resultid="1921" heatid="7855" lane="5" entrytime="00:01:04.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="796" reactiontime="+53" swimtime="00:02:15.70" resultid="1922" heatid="7967" lane="6" entrytime="00:02:04.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:05.14" />
                    <SPLIT distance="150" swimtime="00:01:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="892" reactiontime="+65" swimtime="00:01:04.88" resultid="1923" heatid="8001" lane="4" entrytime="00:01:03.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="877" reactiontime="+58" swimtime="00:00:32.78" resultid="1924" heatid="8047" lane="8" entrytime="00:00:32.25" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PVKBA" nation="SVK" region="BAO" clubid="3594" name="Plavecký Veteránsky Klub Bratislava" shortname="PVK Bratislava">
          <ATHLETES>
            <ATHLETE birthdate="1960-01-01" firstname="Ivica" gender="F" lastname="Forrova" nation="SVK" athleteid="3595">
              <RESULTS>
                <RESULT eventid="1059" points="577" reactiontime="+88" swimtime="00:00:34.22" resultid="3596" heatid="7679" lane="4" entrytime="00:00:33.50" />
                <RESULT eventid="1270" points="503" reactiontime="+85" swimtime="00:01:31.28" resultid="3597" heatid="7832" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="525" reactiontime="+90" swimtime="00:01:39.44" resultid="3598" heatid="7877" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="489" reactiontime="+82" swimtime="00:01:31.65" resultid="3599" heatid="7928" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" status="DNS" swimtime="00:00:00.00" resultid="3600" heatid="8007" lane="1" entrytime="00:03:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Jaroslav" gender="M" lastname="Sykora" nation="SVK" athleteid="3601">
              <RESULTS>
                <RESULT eventid="1076" points="683" reactiontime="+81" swimtime="00:00:26.97" resultid="3602" heatid="7706" lane="6" entrytime="00:00:27.30" />
                <RESULT eventid="1108" points="516" reactiontime="+91" swimtime="00:02:39.38" resultid="3603" heatid="7729" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="100" swimtime="00:01:12.06" />
                    <SPLIT distance="150" swimtime="00:02:01.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="593" reactiontime="+63" swimtime="00:00:32.30" resultid="3604" heatid="7774" lane="3" entrytime="00:00:32.50" />
                <RESULT eventid="1286" points="659" reactiontime="+83" swimtime="00:01:08.71" resultid="3605" heatid="7852" lane="3" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1415" reactiontime="+63" status="DSQ" swimtime="00:00:29.26" resultid="3606" heatid="7920" lane="2" entrytime="00:00:29.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Jozef" gender="M" lastname="Krcik" nation="SVK" athleteid="3607">
              <RESULTS>
                <RESULT eventid="1156" points="723" swimtime="00:21:30.93" resultid="3608" heatid="8720" lane="4" entrytime="00:22:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:20.23" />
                    <SPLIT distance="200" swimtime="00:02:45.08" />
                    <SPLIT distance="300" swimtime="00:04:10.96" />
                    <SPLIT distance="400" swimtime="00:05:37.53" />
                    <SPLIT distance="500" swimtime="00:07:04.53" />
                    <SPLIT distance="600" swimtime="00:08:31.35" />
                    <SPLIT distance="700" swimtime="00:09:58.44" />
                    <SPLIT distance="800" swimtime="00:11:25.67" />
                    <SPLIT distance="900" swimtime="00:12:53.15" />
                    <SPLIT distance="1000" swimtime="00:14:20.83" />
                    <SPLIT distance="1100" swimtime="00:15:47.96" />
                    <SPLIT distance="1200" swimtime="00:17:13.56" />
                    <SPLIT distance="1300" swimtime="00:18:40.00" />
                    <SPLIT distance="1400" swimtime="00:20:06.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="589" reactiontime="+97" swimtime="00:01:22.50" resultid="3609" heatid="7844" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="613" reactiontime="+93" swimtime="00:02:36.92" resultid="3610" heatid="7959" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:02:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="697" reactiontime="+99" swimtime="00:05:25.86" resultid="3611" heatid="9064" lane="2" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:17.38" />
                    <SPLIT distance="150" swimtime="00:01:58.25" />
                    <SPLIT distance="200" swimtime="00:02:39.92" />
                    <SPLIT distance="300" swimtime="00:04:04.26" />
                    <SPLIT distance="350" swimtime="00:04:46.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Laura" gender="F" lastname="Majernikova" nation="SVK" athleteid="3612">
              <RESULTS>
                <RESULT eventid="1140" points="359" swimtime="00:13:30.01" resultid="3613" heatid="8715" lane="3" entrytime="00:15:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                    <SPLIT distance="100" swimtime="00:01:28.07" />
                    <SPLIT distance="200" swimtime="00:03:08.14" />
                    <SPLIT distance="300" swimtime="00:04:51.39" />
                    <SPLIT distance="400" swimtime="00:06:34.84" />
                    <SPLIT distance="500" swimtime="00:08:19.26" />
                    <SPLIT distance="600" swimtime="00:10:05.56" />
                    <SPLIT distance="700" swimtime="00:11:50.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="423" reactiontime="+87" swimtime="00:01:33.95" resultid="3614" heatid="7829" lane="6" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Monika" gender="F" lastname="Novakova" nation="SVK" athleteid="3615">
              <RESULTS>
                <RESULT eventid="1092" points="466" reactiontime="+86" swimtime="00:03:07.23" resultid="3616" heatid="7715" lane="7" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:01:28.04" />
                    <SPLIT distance="150" swimtime="00:02:23.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="453" reactiontime="+81" swimtime="00:03:31.84" resultid="3617" heatid="7781" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.82" />
                    <SPLIT distance="100" swimtime="00:01:41.54" />
                    <SPLIT distance="150" swimtime="00:02:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="405" reactiontime="+94" swimtime="00:03:20.14" resultid="3618" heatid="7858" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="100" swimtime="00:01:33.07" />
                    <SPLIT distance="150" swimtime="00:02:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" status="DNS" swimtime="00:00:00.00" resultid="3619" heatid="8803" lane="7" entrytime="00:07:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Peter" gender="M" lastname="Mansil" nation="SVK" athleteid="3620">
              <RESULTS>
                <RESULT eventid="1076" points="638" reactiontime="+98" swimtime="00:00:30.29" resultid="3621" heatid="7692" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1286" points="582" reactiontime="+105" swimtime="00:01:22.82" resultid="3622" heatid="7844" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="507" reactiontime="+88" swimtime="00:00:38.24" resultid="3623" heatid="8034" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1383" points="474" reactiontime="+99" swimtime="00:01:27.36" resultid="3624" heatid="7886" lane="4" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Peter" gender="M" lastname="Moravec" nation="SVK" athleteid="3625">
              <RESULTS>
                <RESULT eventid="1222" points="457" reactiontime="+89" swimtime="00:03:31.13" resultid="3626" heatid="7788" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:36.60" />
                    <SPLIT distance="150" swimtime="00:02:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="383" reactiontime="+95" swimtime="00:01:33.77" resultid="3627" heatid="7886" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="3628" heatid="8035" lane="5" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Peter" gender="M" lastname="Nahalka" nation="SVK" athleteid="3629">
              <RESULTS>
                <RESULT eventid="1156" status="WDR" swimtime="00:00:00.00" resultid="3630" entrytime="00:29:30.00" />
                <RESULT eventid="1222" status="WDR" swimtime="00:00:00.00" resultid="3631" heatid="7789" lane="3" entrytime="00:03:29.50" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="3632" heatid="7886" lane="5" entrytime="00:01:34.00" />
                <RESULT eventid="1655" status="WDR" swimtime="00:00:00.00" resultid="3633" heatid="8036" lane="3" entrytime="00:00:41.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Petr" gender="M" lastname="Soukup" nation="SVK" athleteid="3634">
              <RESULTS>
                <RESULT eventid="1076" points="670" reactiontime="+92" swimtime="00:00:27.62" resultid="3635" heatid="7705" lane="7" entrytime="00:00:27.80" />
                <RESULT eventid="1254" points="681" reactiontime="+87" swimtime="00:01:00.13" resultid="3636" heatid="7821" lane="5" entrytime="00:01:00.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="606" reactiontime="+92" swimtime="00:02:15.54" resultid="3637" heatid="7964" lane="3" entrytime="00:02:15.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                    <SPLIT distance="150" swimtime="00:01:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="3638" heatid="8043" lane="3" entrytime="00:00:35.60" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="PVK Bratislava D">
              <RESULTS>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="8761" heatid="7868" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3601" number="1" />
                    <RELAYPOSITION athleteid="3620" number="2" />
                    <RELAYPOSITION athleteid="3634" number="3" />
                    <RELAYPOSITION athleteid="3607" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="PVK Bratislava C">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+80" status="EXH" swimtime="00:02:05.40" resultid="8643" heatid="7734" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.62" />
                    <SPLIT distance="100" swimtime="00:01:03.54" />
                    <SPLIT distance="150" swimtime="00:01:37.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3601" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3612" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="3615" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="3634" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="POMOS" nation="RUS" clubid="2703" name="Poseidon Moscow">
          <ATHLETES>
            <ATHLETE birthdate="1946-01-01" firstname="Alexander" gender="M" lastname="Bashmakov" nation="RUS" athleteid="2704">
              <RESULTS>
                <RESULT eventid="1076" points="816" reactiontime="+91" swimtime="00:00:30.14" resultid="2705" heatid="7700" lane="7" entrytime="00:00:29.50" />
                <RESULT eventid="1254" points="782" reactiontime="+90" swimtime="00:01:08.81" resultid="2706" heatid="7814" lane="2" entrytime="00:01:09.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="768" reactiontime="+93" swimtime="00:02:39.34" resultid="2707" heatid="7958" lane="4" entrytime="00:02:40.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:16.76" />
                    <SPLIT distance="150" swimtime="00:01:57.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="502" reactiontime="+86" swimtime="00:03:18.25" resultid="2708" heatid="8014" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                    <SPLIT distance="100" swimtime="00:01:35.02" />
                    <SPLIT distance="150" swimtime="00:02:27.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Vladislav" gender="M" lastname="Zagrabenko" nation="RUS" athleteid="2709">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2710" heatid="7696" lane="7" entrytime="00:00:30.85" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="2711" heatid="7896" lane="1" entrytime="00:01:08.50" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="2712" heatid="8047" lane="5" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Sergey" gender="M" lastname="Petrov" nation="RUS" athleteid="2713">
              <RESULTS>
                <RESULT eventid="1222" points="575" reactiontime="+75" swimtime="00:02:51.76" resultid="2714" heatid="7794" lane="2" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:19.76" />
                    <SPLIT distance="150" swimtime="00:02:04.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="688" reactiontime="+76" swimtime="00:01:14.31" resultid="2715" heatid="7894" lane="8" entrytime="00:01:15.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="615" reactiontime="+74" swimtime="00:00:29.55" resultid="2716" heatid="7922" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="1655" points="745" reactiontime="+72" swimtime="00:00:32.53" resultid="2717" heatid="8045" lane="4" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PRKAL" nation="RUS" clubid="2119" name="Pregel Kaliningrad">
          <ATHLETES>
            <ATHLETE birthdate="1938-02-01" firstname="Luiza" gender="F" lastname="Shcherbich" nation="RUS" athleteid="2120">
              <RESULTS>
                <RESULT eventid="1059" points="245" reactiontime="+153" swimtime="00:01:01.42" resultid="2121" heatid="7671" lane="4" entrytime="00:00:59.50" />
                <RESULT eventid="1206" status="DNS" swimtime="00:00:00.00" resultid="2122" heatid="7778" lane="5" entrytime="00:05:29.00" />
                <RESULT eventid="1270" status="DNS" swimtime="00:00:00.00" resultid="2123" heatid="7827" lane="8" entrytime="00:02:19.00" />
                <RESULT eventid="1366" points="318" reactiontime="+119" swimtime="00:02:43.91" resultid="2124" heatid="7874" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="304" reactiontime="+114" swimtime="00:01:10.10" resultid="2125" heatid="8021" lane="1" entrytime="00:01:09.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-16" firstname="Natalia" gender="F" lastname="Aleskchenko" nation="RUS" athleteid="2126">
              <RESULTS>
                <RESULT eventid="1059" points="659" reactiontime="+89" swimtime="00:00:34.75" resultid="2127" heatid="7678" lane="5" entrytime="00:00:34.80" />
                <RESULT eventid="1092" points="797" reactiontime="+94" swimtime="00:03:04.45" resultid="2128" heatid="7716" lane="1" entrytime="00:03:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:28.17" />
                    <SPLIT distance="150" swimtime="00:02:21.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="700" reactiontime="+92" swimtime="00:01:27.23" resultid="2129" heatid="7832" lane="3" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="748" reactiontime="+88" swimtime="00:00:37.60" resultid="2130" heatid="7901" lane="5" entrytime="00:00:37.80" />
                <RESULT eventid="1463" points="760" reactiontime="+95" swimtime="00:02:47.19" resultid="2131" heatid="7948" lane="5" entrytime="00:02:48.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:21.50" />
                    <SPLIT distance="150" swimtime="00:02:05.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="733" reactiontime="+92" swimtime="00:01:27.22" resultid="2132" heatid="7989" lane="6" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" status="DNS" swimtime="00:00:00.00" resultid="2133" heatid="9049" lane="8" entrytime="00:05:52.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-30" firstname="Marina" gender="F" lastname="Kilina" nation="RUS" athleteid="2134">
              <RESULTS>
                <RESULT eventid="1059" points="630" reactiontime="+103" swimtime="00:00:33.23" resultid="2135" heatid="7679" lane="5" entrytime="00:00:33.80" />
                <RESULT eventid="1092" points="582" reactiontime="+94" swimtime="00:03:06.02" resultid="2136" heatid="7716" lane="7" entrytime="00:03:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:01:27.63" />
                    <SPLIT distance="150" swimtime="00:02:21.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="656" reactiontime="+74" swimtime="00:00:38.21" resultid="2137" heatid="7758" lane="3" entrytime="00:00:39.50" />
                <RESULT eventid="1270" points="692" reactiontime="+94" swimtime="00:01:22.10" resultid="2138" heatid="7833" lane="8" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="618" reactiontime="+86" swimtime="00:01:24.78" resultid="2139" heatid="7929" lane="6" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" status="DNS" swimtime="00:00:00.00" resultid="2140" heatid="8006" lane="3" entrytime="00:03:16.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-07-02" firstname="Svetlana" gender="F" lastname="Smirnova" nation="RUS" athleteid="2141">
              <RESULTS>
                <RESULT eventid="1639" points="190" reactiontime="+111" swimtime="00:00:59.71" resultid="2142" heatid="8023" lane="4" entrytime="00:00:49.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-23" firstname="Akim" gender="M" lastname="Denisenko" nation="RUS" athleteid="2143">
              <RESULTS>
                <RESULT eventid="1076" points="482" reactiontime="+85" swimtime="00:00:34.42" resultid="2144" heatid="7690" lane="6" entrytime="00:00:33.80" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="2145" heatid="7767" lane="2" entrytime="00:00:44.50" />
                <RESULT eventid="1286" points="378" reactiontime="+91" swimtime="00:01:40.19" resultid="2146" heatid="7842" lane="5" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="357" reactiontime="+81" swimtime="00:00:42.17" resultid="2147" heatid="7908" lane="4" entrytime="00:00:41.50" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="2148" heatid="8032" lane="6" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-07-20" firstname="Alexander" gender="M" lastname="Tervinskiy" nation="RUS" athleteid="2149">
              <RESULTS>
                <RESULT eventid="1076" points="543" reactiontime="+83" swimtime="00:00:31.95" resultid="2150" heatid="7690" lane="3" entrytime="00:00:33.80" />
                <RESULT eventid="1190" points="487" reactiontime="+85" swimtime="00:00:39.99" resultid="2151" heatid="7768" lane="7" entrytime="00:00:42.30" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="2152" heatid="7843" lane="2" entrytime="00:01:26.80" />
                <RESULT eventid="1383" points="414" reactiontime="+85" swimtime="00:01:31.35" resultid="2153" heatid="7886" lane="2" entrytime="00:01:34.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="501" reactiontime="+78" swimtime="00:00:38.38" resultid="2154" heatid="8035" lane="1" entrytime="00:00:42.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-08-21" firstname="Grigoriy" gender="M" lastname="Lopin" nation="RUS" athleteid="2155">
              <RESULTS>
                <RESULT eventid="1108" points="322" reactiontime="+120" swimtime="00:03:28.49" resultid="2156" heatid="7723" lane="3" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                    <SPLIT distance="100" swimtime="00:01:33.75" />
                    <SPLIT distance="150" swimtime="00:02:35.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="381" reactiontime="+122" swimtime="00:03:33.30" resultid="2157" heatid="7789" lane="5" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.71" />
                    <SPLIT distance="100" swimtime="00:01:39.06" />
                    <SPLIT distance="150" swimtime="00:02:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="434" reactiontime="+114" swimtime="00:01:31.82" resultid="2158" heatid="7886" lane="6" entrytime="00:01:34.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="470" reactiontime="+100" swimtime="00:00:40.35" resultid="2159" heatid="8036" lane="8" entrytime="00:00:41.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-07-31" firstname="Sergey" gender="M" lastname="Dirindyaev" nation="RUS" athleteid="2160">
              <RESULTS>
                <RESULT eventid="1076" points="585" reactiontime="+102" swimtime="00:00:30.37" resultid="2161" heatid="7696" lane="2" entrytime="00:00:30.80" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="2162" heatid="7768" lane="5" entrytime="00:00:41.80" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="2163" heatid="7814" lane="1" entrytime="00:01:09.50" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="2164" heatid="7912" lane="4" entrytime="00:00:35.50" />
                <RESULT eventid="1655" points="437" reactiontime="+71" swimtime="00:00:41.34" resultid="2165" heatid="8036" lane="1" entrytime="00:00:41.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-04-17" firstname="Vadim" gender="M" lastname="Ezhkov" nation="RUS" athleteid="2166">
              <RESULTS>
                <RESULT eventid="1076" points="515" reactiontime="+75" swimtime="00:00:30.16" resultid="2167" heatid="7696" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1222" points="592" reactiontime="+73" swimtime="00:02:57.69" resultid="2168" heatid="7793" lane="8" entrytime="00:03:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                    <SPLIT distance="100" swimtime="00:01:23.68" />
                    <SPLIT distance="150" swimtime="00:02:10.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="579" reactiontime="+74" swimtime="00:01:20.61" resultid="2169" heatid="7890" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="548" reactiontime="+72" swimtime="00:00:32.30" resultid="2170" heatid="7914" lane="1" entrytime="00:00:34.50" />
                <RESULT eventid="1655" points="633" reactiontime="+70" swimtime="00:00:35.73" resultid="2171" heatid="8041" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-12-05" firstname="Vladimir" gender="M" lastname="Chekutov" nation="RUS" athleteid="2172">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2173" heatid="7702" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="2174" heatid="7774" lane="8" entrytime="00:00:33.50" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="2176" heatid="7850" lane="6" entrytime="00:01:13.50" />
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="2177" heatid="7939" lane="4" entrytime="00:01:14.50" />
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="2178" heatid="8016" lane="3" entrytime="00:02:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-03-26" firstname="Alexander" gender="M" lastname="Smirnov" nation="RUS" athleteid="2179">
              <RESULTS>
                <RESULT eventid="1156" points="573" swimtime="00:19:49.74" resultid="2180" heatid="8718" lane="2" entrytime="00:20:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="200" swimtime="00:02:34.10" />
                    <SPLIT distance="300" swimtime="00:03:53.07" />
                    <SPLIT distance="400" swimtime="00:05:12.45" />
                    <SPLIT distance="500" swimtime="00:06:31.39" />
                    <SPLIT distance="600" swimtime="00:07:50.54" />
                    <SPLIT distance="700" swimtime="00:09:10.01" />
                    <SPLIT distance="800" swimtime="00:10:29.94" />
                    <SPLIT distance="900" swimtime="00:11:50.29" />
                    <SPLIT distance="1000" swimtime="00:13:10.57" />
                    <SPLIT distance="1100" swimtime="00:14:31.14" />
                    <SPLIT distance="1200" swimtime="00:15:52.21" />
                    <SPLIT distance="1300" swimtime="00:17:12.50" />
                    <SPLIT distance="1400" swimtime="00:18:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="605" reactiontime="+83" swimtime="00:02:15.62" resultid="2181" heatid="7963" lane="6" entrytime="00:02:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="604" reactiontime="+85" swimtime="00:04:50.78" resultid="2182" heatid="9062" lane="5" entrytime="00:05:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:09.84" />
                    <SPLIT distance="150" swimtime="00:01:47.60" />
                    <SPLIT distance="200" swimtime="00:02:25.13" />
                    <SPLIT distance="250" swimtime="00:03:02.40" />
                    <SPLIT distance="300" swimtime="00:03:39.95" />
                    <SPLIT distance="350" swimtime="00:04:16.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-09" firstname="Vladimir" gender="M" lastname="Polyakov" nation="RUS" athleteid="2183">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2184" heatid="7696" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="2185" heatid="7812" lane="8" entrytime="00:01:12.50" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="2186" heatid="7913" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="2187" heatid="8036" lane="2" entrytime="00:00:41.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Sergey" gender="M" lastname="Katakchiev" nation="RUS" athleteid="6336">
              <RESULTS>
                <RESULT eventid="1190" points="679" reactiontime="+73" swimtime="00:00:32.60" resultid="6337" heatid="7774" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1286" points="706" reactiontime="+81" swimtime="00:01:07.93" resultid="6338" heatid="7851" lane="3" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="669" reactiontime="+75" swimtime="00:01:11.04" resultid="6339" heatid="7940" lane="6" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="702" reactiontime="+75" swimtime="00:02:33.32" resultid="6340" heatid="8018" lane="8" entrytime="00:02:37.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:13.32" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Tatiana" gender="F" lastname="Logvinova" nation="RUS" athleteid="6777">
              <RESULTS>
                <RESULT eventid="1059" points="439" reactiontime="+86" swimtime="00:00:36.53" resultid="6778" heatid="7677" lane="6" entrytime="00:00:35.50" />
                <RESULT eventid="1173" points="404" reactiontime="+68" swimtime="00:00:44.05" resultid="6779" heatid="7757" lane="1" entrytime="00:00:43.50" />
                <RESULT eventid="1270" points="424" reactiontime="+83" swimtime="00:01:33.86" resultid="6780" heatid="7830" lane="4" entrytime="00:01:31.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" status="DNS" swimtime="00:00:00.00" resultid="6781" heatid="7877" lane="5" entrytime="00:01:39.50" />
                <RESULT eventid="1639" points="480" reactiontime="+92" swimtime="00:00:45.24" resultid="6782" heatid="8026" lane="8" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Pregel Kaliningrad D" number="1">
              <RESULTS>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="2189" heatid="7870" lane="8" entrytime="00:02:18.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6336" number="1" />
                    <RELAYPOSITION athleteid="2179" number="2" />
                    <RELAYPOSITION athleteid="2160" number="3" />
                    <RELAYPOSITION athleteid="2143" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" reactiontime="+97" swimtime="00:02:02.79" resultid="2190" heatid="7971" lane="4" entrytime="00:02:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.27" />
                    <SPLIT distance="100" swimtime="00:00:58.24" />
                    <SPLIT distance="150" swimtime="00:01:29.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6336" number="1" />
                    <RELAYPOSITION athleteid="2179" number="2" />
                    <RELAYPOSITION athleteid="2160" number="3" />
                    <RELAYPOSITION athleteid="2143" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Pregel Kaliningrad D" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+83" swimtime="00:02:05.44" resultid="2188" heatid="7735" lane="3" entrytime="00:02:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                    <SPLIT distance="100" swimtime="00:00:58.43" />
                    <SPLIT distance="150" swimtime="00:01:32.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2172" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2166" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="2126" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="2134" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" status="DNS" swimtime="00:00:00.00" resultid="2191" heatid="8052" lane="6" entrytime="00:02:09.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2172" number="1" />
                    <RELAYPOSITION athleteid="2166" number="2" />
                    <RELAYPOSITION athleteid="2126" number="3" />
                    <RELAYPOSITION athleteid="2134" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02705" nation="POL" region="05" clubid="2296" name="Pływak Tomaszów Maz.">
          <CONTACT email="tsplywak@wp.pl" name="Bucholz" phone="606135860" />
          <ATHLETES>
            <ATHLETE birthdate="1979-03-01" firstname="Gabriela" gender="F" lastname="Kozłowska" nation="POL" athleteid="2297">
              <RESULTS>
                <RESULT eventid="1238" points="361" reactiontime="+86" swimtime="00:01:20.71" resultid="2298" heatid="7799" lane="5" entrytime="00:01:26.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="277" reactiontime="+93" swimtime="00:01:39.83" resultid="2299" heatid="7830" lane="2" entrytime="00:01:35.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-02" firstname="Bernard" gender="M" lastname="Wierzbik" nation="POL" athleteid="2300">
              <RESULTS>
                <RESULT eventid="1286" points="366" reactiontime="+84" swimtime="00:01:22.50" resultid="2301" heatid="7845" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="447" reactiontime="+92" swimtime="00:00:33.55" resultid="2302" heatid="7915" lane="8" entrytime="00:00:33.50" />
                <RESULT eventid="1479" points="293" reactiontime="+94" swimtime="00:02:47.68" resultid="2303" heatid="7960" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:04.46" />
                    <SPLIT distance="100" swimtime="00:02:47.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="351" reactiontime="+95" swimtime="00:01:20.54" resultid="2304" heatid="7997" lane="2" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="REWRO" nation="POL" region="01" clubid="3988" name="Redeco Wrocław">
          <CONTACT city="Wrocław" name="Wolny Dariusz" phone="603630870" state="DOL" street="Rogowska 52a" zip="54-440" />
          <ATHLETES>
            <ATHLETE birthdate="1974-01-25" firstname="Marlena" gender="F" lastname="Jakubów" nation="POL" athleteid="4017">
              <RESULTS>
                <RESULT eventid="1059" points="442" reactiontime="+113" swimtime="00:00:35.64" resultid="4018" heatid="7678" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1092" points="321" reactiontime="+126" swimtime="00:03:32.13" resultid="4019" heatid="7716" lane="8" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.76" />
                    <SPLIT distance="100" swimtime="00:01:42.43" />
                    <SPLIT distance="150" swimtime="00:02:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="365" swimtime="00:00:44.61" resultid="4020" heatid="7756" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1270" points="380" reactiontime="+110" swimtime="00:01:33.70" resultid="4021" heatid="7830" lane="7" entrytime="00:01:35.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="267" swimtime="00:01:42.34" resultid="4022" heatid="7927" lane="2" entrytime="00:01:37.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="300" reactiontime="+121" swimtime="00:03:11.36" resultid="4023" heatid="7947" lane="6" entrytime="00:03:03.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                    <SPLIT distance="100" swimtime="00:01:31.13" />
                    <SPLIT distance="150" swimtime="00:02:23.58" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G4 - Wykonanie więcej niż jednego pociągnięcia ramieniem (lub obydwoma ramionami jednocześnie) po obróceniu się na piersi, w trakcie wykonywania nawrotu  (Czas: 10:04)" eventid="1607" reactiontime="+107" status="DSQ" swimtime="00:03:41.34" resultid="4024" heatid="8007" lane="6" entrytime="00:03:11.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.98" />
                    <SPLIT distance="100" swimtime="00:01:48.70" />
                    <SPLIT distance="150" swimtime="00:02:46.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="268" reactiontime="+105" swimtime="00:07:03.23" resultid="4025" heatid="9051" lane="7" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                    <SPLIT distance="100" swimtime="00:01:34.46" />
                    <SPLIT distance="150" swimtime="00:02:30.41" />
                    <SPLIT distance="200" swimtime="00:03:25.46" />
                    <SPLIT distance="250" swimtime="00:04:22.97" />
                    <SPLIT distance="300" swimtime="00:05:17.88" />
                    <SPLIT distance="350" swimtime="00:06:14.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-27" firstname="Hanna" gender="F" lastname="Sikacz" nation="POL" athleteid="4026">
              <RESULTS>
                <RESULT eventid="1140" points="491" swimtime="00:12:12.71" resultid="4027" heatid="8713" lane="1" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:24.86" />
                    <SPLIT distance="200" swimtime="00:02:55.73" />
                    <SPLIT distance="300" swimtime="00:04:27.77" />
                    <SPLIT distance="400" swimtime="00:05:59.89" />
                    <SPLIT distance="500" swimtime="00:07:35.57" />
                    <SPLIT distance="600" swimtime="00:09:10.33" />
                    <SPLIT distance="700" swimtime="00:10:43.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="459" reactiontime="+76" swimtime="00:01:14.48" resultid="4028" heatid="7801" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="408" reactiontime="+75" swimtime="00:01:27.72" resultid="4029" heatid="7830" lane="5" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="425" reactiontime="+74" swimtime="00:02:47.45" resultid="4030" heatid="7948" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:02:02.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="409" reactiontime="+81" swimtime="00:06:50.05" resultid="4031" heatid="8802" lane="8" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:41.90" />
                    <SPLIT distance="150" swimtime="00:02:34.02" />
                    <SPLIT distance="200" swimtime="00:03:26.85" />
                    <SPLIT distance="250" swimtime="00:04:22.81" />
                    <SPLIT distance="300" swimtime="00:05:20.83" />
                    <SPLIT distance="350" swimtime="00:06:07.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="395" reactiontime="+77" swimtime="00:03:12.97" resultid="4032" heatid="8007" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                    <SPLIT distance="100" swimtime="00:01:33.20" />
                    <SPLIT distance="150" swimtime="00:02:23.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="481" reactiontime="+82" swimtime="00:05:48.99" resultid="4033" heatid="9050" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:23.05" />
                    <SPLIT distance="150" swimtime="00:02:07.97" />
                    <SPLIT distance="200" swimtime="00:02:53.61" />
                    <SPLIT distance="250" swimtime="00:03:39.77" />
                    <SPLIT distance="300" swimtime="00:04:24.88" />
                    <SPLIT distance="350" swimtime="00:05:09.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-03-21" firstname="Dariusz" gender="M" lastname="Wolny" nation="POL" athleteid="4034">
              <RESULTS>
                <RESULT eventid="1108" points="947" reactiontime="+79" swimtime="00:02:25.53" resultid="4035" heatid="7732" lane="8" entrytime="00:02:26.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:07.30" />
                    <SPLIT distance="150" swimtime="00:01:50.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="859" reactiontime="+69" swimtime="00:00:30.90" resultid="4036" heatid="7775" lane="4" entrytime="00:00:30.30" />
                <RESULT eventid="1286" points="931" reactiontime="+79" swimtime="00:01:07.05" resultid="4037" heatid="7853" lane="5" entrytime="00:01:07.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="927" reactiontime="+73" swimtime="00:01:06.50" resultid="4038" heatid="7941" lane="5" entrytime="00:01:07.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="995" reactiontime="+70" swimtime="00:02:25.19" resultid="4039" heatid="8019" lane="2" entrytime="00:02:26.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:09.18" />
                    <SPLIT distance="150" swimtime="00:01:46.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-23" firstname="Agnieszka" gender="F" lastname="Bystrzycka" nation="POL" athleteid="4040">
              <RESULTS>
                <RESULT eventid="1059" points="834" reactiontime="+81" swimtime="00:00:27.76" resultid="4041" heatid="7683" lane="3" entrytime="00:00:28.49" />
                <RESULT eventid="1206" points="865" reactiontime="+82" swimtime="00:02:43.91" resultid="4042" heatid="7783" lane="4" entrytime="00:02:44.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:17.99" />
                    <SPLIT distance="150" swimtime="00:02:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="922" reactiontime="+83" swimtime="00:01:14.66" resultid="4043" heatid="7880" lane="4" entrytime="00:01:14.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="882" reactiontime="+80" swimtime="00:00:30.30" resultid="4044" heatid="7905" lane="3" entrytime="00:00:31.49" />
                <RESULT eventid="1639" points="818" reactiontime="+78" swimtime="00:00:33.94" resultid="4045" heatid="8028" lane="4" entrytime="00:00:33.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-02-28" firstname="Magdalena" gender="F" lastname="Mongiało" nation="POL" athleteid="4046">
              <RESULTS>
                <RESULT eventid="1059" points="815" reactiontime="+76" swimtime="00:00:28.39" resultid="4047" heatid="7683" lane="6" entrytime="00:00:28.49" />
                <RESULT eventid="1140" points="675" reactiontime="+91" swimtime="00:10:34.27" resultid="4048" heatid="8712" lane="5" entrytime="00:10:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:50.04" />
                    <SPLIT distance="200" swimtime="00:02:29.61" />
                    <SPLIT distance="250" swimtime="00:03:09.12" />
                    <SPLIT distance="300" swimtime="00:03:49.23" />
                    <SPLIT distance="350" swimtime="00:04:29.41" />
                    <SPLIT distance="400" swimtime="00:05:09.75" />
                    <SPLIT distance="450" swimtime="00:05:50.21" />
                    <SPLIT distance="500" swimtime="00:06:30.74" />
                    <SPLIT distance="550" swimtime="00:07:11.63" />
                    <SPLIT distance="600" swimtime="00:07:53.03" />
                    <SPLIT distance="650" swimtime="00:08:34.53" />
                    <SPLIT distance="700" swimtime="00:09:15.11" />
                    <SPLIT distance="750" swimtime="00:09:55.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="808" reactiontime="+81" swimtime="00:01:02.68" resultid="4049" heatid="7805" lane="7" entrytime="00:01:03.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="747" reactiontime="+89" swimtime="00:02:18.94" resultid="4050" heatid="7951" lane="5" entrytime="00:02:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="613" reactiontime="+88" swimtime="00:05:15.21" resultid="4051" heatid="9047" lane="7" entrytime="00:05:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:51.90" />
                    <SPLIT distance="200" swimtime="00:02:32.75" />
                    <SPLIT distance="250" swimtime="00:03:16.03" />
                    <SPLIT distance="300" swimtime="00:03:57.46" />
                    <SPLIT distance="350" swimtime="00:04:36.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-13" firstname="Kazimiera" gender="F" lastname="Syguła" nation="POL" athleteid="4052">
              <RESULTS>
                <RESULT eventid="1059" points="341" reactiontime="+115" swimtime="00:00:46.16" resultid="4053" heatid="7672" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1173" points="436" reactiontime="+77" swimtime="00:00:52.78" resultid="4054" heatid="7755" lane="8" entrytime="00:00:54.20" />
                <RESULT eventid="1238" points="287" reactiontime="+116" swimtime="00:01:47.51" resultid="4055" heatid="7797" lane="3" entrytime="00:01:49.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="464" reactiontime="+82" swimtime="00:01:54.64" resultid="4056" heatid="7927" lane="7" entrytime="00:01:57.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-03" firstname="Łukasz" gender="M" lastname="Hałada" nation="POL" athleteid="4057">
              <RESULTS>
                <RESULT eventid="1076" points="540" reactiontime="+76" swimtime="00:00:27.17" resultid="4058" heatid="7706" lane="2" entrytime="00:00:27.30" />
                <RESULT eventid="1190" points="588" reactiontime="+73" swimtime="00:00:31.63" resultid="4059" heatid="7774" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1254" points="500" reactiontime="+80" swimtime="00:01:01.75" resultid="4060" heatid="7820" lane="8" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="575" reactiontime="+73" swimtime="00:01:09.21" resultid="4061" heatid="7941" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="415" reactiontime="+71" swimtime="00:02:36.27" resultid="4062" heatid="8017" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:55.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-01" firstname="Wojciech" gender="M" lastname="Dobrowolski" nation="POL" athleteid="4063">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4064" heatid="7698" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="4065" heatid="7818" lane="8" entrytime="00:01:04.85" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="4066" heatid="7915" lane="3" entrytime="00:00:32.99" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="4067" heatid="7997" lane="1" entrytime="00:01:21.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-26" firstname="Wojciech" gender="M" lastname="Urban" nation="POL" athleteid="4068">
              <RESULTS>
                <RESULT eventid="1076" points="650" reactiontime="+71" swimtime="00:00:25.54" resultid="4069" heatid="7711" lane="4" entrytime="00:00:25.40" />
                <RESULT eventid="1254" points="602" reactiontime="+75" swimtime="00:00:58.06" resultid="4070" heatid="7824" lane="2" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="498" reactiontime="+78" swimtime="00:00:28.84" resultid="4071" heatid="7923" lane="3" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-28" firstname="Maciej" gender="M" lastname="Kownacki" nation="POL" athleteid="4072">
              <RESULTS>
                <RESULT eventid="1076" points="692" reactiontime="+88" swimtime="00:00:25.82" resultid="4073" heatid="7711" lane="2" entrytime="00:00:25.80" />
                <RESULT eventid="1254" points="630" reactiontime="+85" swimtime="00:00:56.66" resultid="4074" heatid="7823" lane="3" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="607" reactiontime="+88" swimtime="00:00:27.98" resultid="4075" heatid="7923" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1479" points="682" reactiontime="+85" swimtime="00:02:07.86" resultid="4076" heatid="7965" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                    <SPLIT distance="100" swimtime="00:01:01.55" />
                    <SPLIT distance="150" swimtime="00:01:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="614" reactiontime="+88" swimtime="00:01:03.43" resultid="4077" heatid="8000" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-28" firstname="Przemek" gender="M" lastname="Marek" nation="POL" athleteid="4078">
              <RESULTS>
                <RESULT eventid="1076" points="527" reactiontime="+79" swimtime="00:00:27.39" resultid="4079" heatid="7705" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="1254" points="494" reactiontime="+77" swimtime="00:01:02.03" resultid="4080" heatid="7818" lane="1" entrytime="00:01:04.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="425" reactiontime="+79" swimtime="00:00:30.40" resultid="4081" heatid="7919" lane="7" entrytime="00:00:30.30" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="4082" heatid="7961" lane="6" entrytime="00:02:28.00" />
                <RESULT eventid="1591" points="421" reactiontime="+75" swimtime="00:01:10.21" resultid="4083" heatid="7998" lane="4" entrytime="00:01:14.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-07" firstname="Łukasz" gender="M" lastname="Ptak" nation="POL" athleteid="4084">
              <RESULTS>
                <RESULT eventid="1222" points="801" reactiontime="+83" swimtime="00:02:31.30" resultid="4085" heatid="7795" lane="3" entrytime="00:02:32.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:52.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="578" reactiontime="+84" swimtime="00:01:06.00" resultid="4086" heatid="7856" lane="1" entrytime="00:01:03.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="734" reactiontime="+86" swimtime="00:01:07.99" resultid="4087" heatid="7896" lane="3" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="738" reactiontime="+82" swimtime="00:00:30.77" resultid="4088" heatid="8048" lane="5" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Dariusz" gender="M" lastname="Patrzałek" nation="POL" athleteid="4089">
              <RESULTS>
                <RESULT eventid="1222" points="206" reactiontime="+109" swimtime="00:04:35.23" resultid="4090" heatid="7787" lane="8" entrytime="00:03:55.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.69" />
                    <SPLIT distance="100" swimtime="00:01:57.90" />
                    <SPLIT distance="150" swimtime="00:03:11.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="234" reactiontime="+112" swimtime="00:01:34.04" resultid="4091" heatid="7810" lane="8" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="4092" heatid="7883" lane="8" entrytime="00:01:50.00" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="4093" heatid="7908" lane="2" entrytime="00:00:44.63" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="4094" heatid="8031" lane="5" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Małgorzata" gender="F" lastname="Garbarek" nation="POL" athleteid="4095">
              <RESULTS>
                <RESULT eventid="1059" points="420" reactiontime="+82" swimtime="00:00:34.88" resultid="4096" heatid="7678" lane="4" entrytime="00:00:34.50" />
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="4097" heatid="7803" lane="3" entrytime="00:01:09.09" />
                <RESULT eventid="1366" status="DNS" swimtime="00:00:00.00" resultid="4098" heatid="7876" lane="4" entrytime="00:01:45.00" />
                <RESULT eventid="1399" status="DNS" swimtime="00:00:00.00" resultid="4099" heatid="7901" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1639" points="332" reactiontime="+77" swimtime="00:00:45.85" resultid="4100" heatid="8026" lane="1" entrytime="00:00:44.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-16" firstname="Mariusz" gender="M" lastname="Bazanowski" nation="POL" athleteid="4101">
              <RESULTS>
                <RESULT eventid="1076" points="535" reactiontime="+85" swimtime="00:00:29.21" resultid="4102" heatid="7700" lane="6" entrytime="00:00:29.29" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="4103" heatid="7816" lane="3" entrytime="00:01:05.55" />
                <RESULT eventid="1415" points="436" reactiontime="+82" swimtime="00:00:33.84" resultid="4104" heatid="7914" lane="7" entrytime="00:00:34.34" />
                <RESULT eventid="1655" points="412" reactiontime="+79" swimtime="00:00:38.77" resultid="4105" heatid="8039" lane="3" entrytime="00:00:38.38" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-17" firstname="Jakub" gender="M" lastname="Piątkowski" nation="POL" athleteid="4106">
              <RESULTS>
                <RESULT eventid="1076" points="593" reactiontime="+72" swimtime="00:00:26.34" resultid="4107" heatid="7711" lane="6" entrytime="00:00:25.55" />
                <RESULT eventid="1190" points="695" reactiontime="+68" swimtime="00:00:29.91" resultid="4108" heatid="7776" lane="5" entrytime="00:00:29.99" />
                <RESULT eventid="1286" points="580" reactiontime="+71" swimtime="00:01:05.94" resultid="4109" heatid="7855" lane="1" entrytime="00:01:05.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="538" reactiontime="+79" swimtime="00:01:15.40" resultid="4110" heatid="7895" lane="4" entrytime="00:01:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="452" reactiontime="+75" swimtime="00:00:29.80" resultid="4111" heatid="7922" lane="2" entrytime="00:00:28.55" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="4112" heatid="8046" lane="5" entrytime="00:00:32.88" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Redeco Wrocław B" number="1">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+83" swimtime="00:01:45.41" resultid="4119" heatid="7973" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                    <SPLIT distance="100" swimtime="00:00:53.92" />
                    <SPLIT distance="150" swimtime="00:01:19.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4057" number="1" />
                    <RELAYPOSITION athleteid="4084" number="2" />
                    <RELAYPOSITION athleteid="4106" number="3" />
                    <RELAYPOSITION athleteid="4068" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1357" reactiontime="+69" swimtime="00:01:55.73" resultid="4120" heatid="7871" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="100" swimtime="00:01:00.40" />
                    <SPLIT distance="150" swimtime="00:01:30.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4106" number="1" />
                    <RELAYPOSITION athleteid="4084" number="2" />
                    <RELAYPOSITION athleteid="4078" number="3" />
                    <RELAYPOSITION athleteid="4068" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Redeco Wrocław B" number="2">
              <RESULTS>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="4121" heatid="7972" lane="2" entrytime="00:01:59.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4034" number="1" />
                    <RELAYPOSITION athleteid="4078" number="2" />
                    <RELAYPOSITION athleteid="4072" number="3" />
                    <RELAYPOSITION athleteid="4101" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1357" reactiontime="+69" swimtime="00:02:03.66" resultid="4122" heatid="7870" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                    <SPLIT distance="150" swimtime="00:01:35.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4057" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4063" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4072" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4101" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Redeco Wrocław B" number="1">
              <RESULTS>
                <RESULT eventid="1495" status="DNS" swimtime="00:00:00.00" resultid="4117" heatid="7969" lane="3" entrytime="00:02:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4040" number="1" />
                    <RELAYPOSITION athleteid="4095" number="2" />
                    <RELAYPOSITION athleteid="4046" number="3" />
                    <RELAYPOSITION athleteid="4026" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" reactiontime="+73" swimtime="00:02:29.20" resultid="4118" heatid="7867" lane="3" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:01:22.96" />
                    <SPLIT distance="150" swimtime="00:01:53.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4046" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4095" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4040" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="4026" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="Redeco Wrocław A" number="1">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+73" swimtime="00:02:02.47" resultid="4113" heatid="8052" lane="5" entrytime="00:02:02.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:06.67" />
                    <SPLIT distance="150" swimtime="00:01:34.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4057" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4040" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4072" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="4046" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1124" reactiontime="+77" swimtime="00:01:47.05" resultid="4114" heatid="7737" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                    <SPLIT distance="100" swimtime="00:00:55.71" />
                    <SPLIT distance="150" swimtime="00:01:21.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4040" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4106" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="4072" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4046" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Redeco Wrocław C" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+76" swimtime="00:02:04.17" resultid="4115" heatid="7737" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                    <SPLIT distance="100" swimtime="00:00:54.54" />
                    <SPLIT distance="150" swimtime="00:01:28.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4034" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4078" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="4026" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="4017" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" status="DNS" swimtime="00:00:00.00" resultid="4116" heatid="8051" lane="1" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4034" number="1" />
                    <RELAYPOSITION athleteid="4017" number="2" />
                    <RELAYPOSITION athleteid="4026" number="3" />
                    <RELAYPOSITION athleteid="4078" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SGGWA" nation="POL" region="14" clubid="2204" name="SGGW Warszawa">
          <CONTACT city="Warszawa" email="olszewski.krzysiek.pl@gmail.com" name="Olszewski Krzysztof" phone="512828406" state="MAZOW" street="Nowoursynowska 166" zip="02-787" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-28" firstname="Krzysztof" gender="M" lastname="Olszewski" nation="POL" athleteid="2205">
              <RESULTS>
                <RESULT eventid="1108" points="555" reactiontime="+75" swimtime="00:02:34.50" resultid="2206" heatid="7729" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="150" swimtime="00:01:54.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="589" reactiontime="+75" swimtime="00:02:46.43" resultid="2207" heatid="7793" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:01:20.93" />
                    <SPLIT distance="150" swimtime="00:02:03.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="668" reactiontime="+75" swimtime="00:01:05.69" resultid="2208" heatid="7853" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="571" reactiontime="+78" swimtime="00:01:14.43" resultid="2209" heatid="7894" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="633" reactiontime="+73" swimtime="00:00:32.90" resultid="2210" heatid="8044" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1703" points="459" reactiontime="+73" swimtime="00:05:18.16" resultid="2211" heatid="9063" lane="4" entrytime="00:05:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:08.75" />
                    <SPLIT distance="150" swimtime="00:01:47.52" />
                    <SPLIT distance="200" swimtime="00:02:27.58" />
                    <SPLIT distance="250" swimtime="00:03:08.80" />
                    <SPLIT distance="300" swimtime="00:03:51.77" />
                    <SPLIT distance="350" swimtime="00:04:36.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="F" lastname="Nawrocka" nation="POL" athleteid="2212">
              <RESULTS>
                <RESULT eventid="1092" points="696" reactiontime="+91" swimtime="00:02:41.39" resultid="2213" heatid="7718" lane="7" entrytime="00:02:47.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:16.94" />
                    <SPLIT distance="150" swimtime="00:02:04.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="584" reactiontime="+75" swimtime="00:00:36.25" resultid="2214" heatid="7761" lane="1" entrytime="00:00:34.40" />
                <RESULT eventid="1270" points="669" reactiontime="+88" swimtime="00:01:14.42" resultid="2215" heatid="7837" lane="8" entrytime="00:01:13.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="565" reactiontime="+94" swimtime="00:01:26.53" resultid="2216" heatid="7879" lane="6" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="550" reactiontime="+93" swimtime="00:00:34.94" resultid="2217" heatid="7903" lane="3" entrytime="00:00:34.90" />
                <RESULT eventid="1574" points="493" reactiontime="+92" swimtime="00:01:20.40" resultid="2218" heatid="7990" lane="8" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="548" reactiontime="+97" swimtime="00:00:40.12" resultid="2219" heatid="8027" lane="4" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCHU" nation="CZE" clubid="2509" name="SK Spolchemie Usti nad Labem" shortname="Spolchemie Usti n/L">
          <CONTACT city="Praha" email="benova.dana@seznam.cz" name="SK Spolchemie Usti nad Labem" phone="+420728212656" street="Tupolevova 466" zip="199 00" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-26" firstname="Dana" gender="F" lastname="Benova" nation="CZE" license="565126" athleteid="2529">
              <RESULTS>
                <RESULT eventid="1206" points="235" reactiontime="+86" swimtime="00:05:00.16" resultid="2530" heatid="7778" lane="4" entrytime="00:05:05.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.71" />
                    <SPLIT distance="100" swimtime="00:02:20.51" />
                    <SPLIT distance="150" swimtime="00:03:42.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="199" reactiontime="+72" swimtime="00:02:12.71" resultid="2531" heatid="7827" lane="2" entrytime="00:02:10.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="228" reactiontime="+83" swimtime="00:02:16.81" resultid="2532" heatid="7874" lane="2" entrytime="00:02:18.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" status="DNS" swimtime="00:00:00.00" resultid="2533" heatid="7926" lane="4" entrytime="00:02:06.30" entrycourse="SCM" />
                <RESULT eventid="1527" points="184" reactiontime="+84" swimtime="00:10:49.43" resultid="2534" heatid="8804" lane="4" entrytime="00:10:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.97" />
                    <SPLIT distance="100" swimtime="00:03:23.57" />
                    <SPLIT distance="150" swimtime="00:04:45.32" />
                    <SPLIT distance="200" swimtime="00:06:01.42" />
                    <SPLIT distance="250" swimtime="00:07:15.49" />
                    <SPLIT distance="300" swimtime="00:08:30.97" />
                    <SPLIT distance="350" swimtime="00:09:41.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-10" firstname="Vaclav" gender="M" lastname="Valtr" nation="CZE" license="560710" athleteid="2535">
              <RESULTS>
                <RESULT comment="K16 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu  (Czas: 11:03)" eventid="1222" reactiontime="+82" status="DSQ" swimtime="00:03:05.16" resultid="2536" heatid="7791" lane="5" entrytime="00:03:10.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:28.13" />
                    <SPLIT distance="150" swimtime="00:02:16.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="840" reactiontime="+83" swimtime="00:01:13.30" resultid="2537" heatid="7848" lane="1" entrytime="00:01:15.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="739" reactiontime="+83" swimtime="00:00:31.54" resultid="2538" heatid="7915" lane="4" entrytime="00:00:32.20" entrycourse="SCM" />
                <RESULT eventid="1447" points="740" reactiontime="+77" swimtime="00:01:15.87" resultid="2539" heatid="7939" lane="2" entrytime="00:01:15.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="640" reactiontime="+90" status="EXH" swimtime="00:06:16.08" resultid="2540" heatid="8809" lane="2" entrytime="00:06:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                    <SPLIT distance="100" swimtime="00:01:29.78" />
                    <SPLIT distance="150" swimtime="00:02:17.82" />
                    <SPLIT distance="200" swimtime="00:03:05.24" />
                    <SPLIT distance="250" swimtime="00:03:57.82" />
                    <SPLIT distance="300" swimtime="00:04:50.86" />
                    <SPLIT distance="350" swimtime="00:05:34.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LEWAR" nation="POL" region="14" clubid="5719" name="SKP Legia Warszawa" shortname="Legia Warszawa">
          <CONTACT email="janek@plywanielegia.pl" name="Drzewiński" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1987-04-27" firstname="Jan" gender="M" lastname="Peńsko" nation="POL" athleteid="5727">
              <RESULTS>
                <RESULT eventid="1254" points="716" reactiontime="+76" swimtime="00:00:54.30" resultid="5728" heatid="7825" lane="7" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="828" reactiontime="+79" swimtime="00:00:57.43" resultid="5729" heatid="8003" lane="5" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-23" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" athleteid="5730">
              <RESULTS>
                <RESULT eventid="1076" points="589" reactiontime="+72" swimtime="00:00:26.40" resultid="5731" heatid="7709" lane="3" entrytime="00:00:26.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-26" firstname="Tomasz" gender="M" lastname="Wilczęga" nation="POL" athleteid="5732">
              <RESULTS>
                <RESULT eventid="1076" points="634" reactiontime="+72" swimtime="00:00:26.58" resultid="5733" heatid="7707" lane="2" entrytime="00:00:27.00" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="5734" heatid="7922" lane="5" entrytime="00:00:28.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-10" firstname="Krzysztof" gender="M" lastname="Spyra" nation="POL" athleteid="5735">
              <RESULTS>
                <RESULT eventid="1076" points="673" reactiontime="+78" swimtime="00:00:27.10" resultid="5736" heatid="7707" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1254" points="668" reactiontime="+77" swimtime="00:00:59.56" resultid="5737" heatid="7823" lane="8" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="5738" heatid="7966" lane="6" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-05" firstname="Maciej" gender="M" lastname="Grzelak" nation="POL" athleteid="5739">
              <RESULTS>
                <RESULT eventid="1076" points="445" reactiontime="+79" swimtime="00:00:31.11" resultid="5740" heatid="7694" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="1108" points="349" reactiontime="+77" swimtime="00:03:01.59" resultid="5741" heatid="7726" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:25.08" />
                    <SPLIT distance="150" swimtime="00:02:19.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="432" reactiontime="+71" swimtime="00:01:19.09" resultid="5742" heatid="7844" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="269" reactiontime="+96" swimtime="00:03:15.16" resultid="5743" heatid="7863" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:01:26.28" />
                    <SPLIT distance="150" swimtime="00:02:19.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="452" reactiontime="+82" swimtime="00:00:32.73" resultid="5744" heatid="7913" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1543" status="WDR" swimtime="00:00:00.00" resultid="5745" entrytime="00:07:00.00" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="5746" heatid="7997" lane="4" entrytime="00:01:17.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-09" firstname="Łukasz" gender="M" lastname="Drzewiński" nation="POL" athleteid="5747">
              <RESULTS>
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="5748" heatid="8003" lane="3" entrytime="00:00:57.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-06-23" firstname="Krzysztof" gender="M" lastname="Micorek" nation="POL" athleteid="5749">
              <RESULTS>
                <RESULT eventid="1254" points="757" reactiontime="+79" swimtime="00:00:55.85" resultid="5750" heatid="7824" lane="4" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="761" reactiontime="+80" swimtime="00:00:27.37" resultid="5751" heatid="7923" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="1591" points="624" reactiontime="+81" swimtime="00:01:04.49" resultid="5752" heatid="8003" lane="8" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="6324" heatid="8047" lane="1" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-09-03" firstname="Urszula" gender="F" lastname="Pawlikowska" nation="POL" athleteid="6691">
              <RESULTS>
                <RESULT eventid="1059" points="490" reactiontime="+78" swimtime="00:00:34.45" resultid="6692" heatid="7679" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="6693" heatid="7801" lane="7" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Legia Warszawa B">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+74" swimtime="00:01:43.13" resultid="5753" heatid="7974" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.07" />
                    <SPLIT distance="100" swimtime="00:00:53.00" />
                    <SPLIT distance="150" swimtime="00:01:18.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5735" number="1" />
                    <RELAYPOSITION athleteid="5732" number="2" />
                    <RELAYPOSITION athleteid="5730" number="3" />
                    <RELAYPOSITION athleteid="5727" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1357" reactiontime="+80" swimtime="00:01:56.25" resultid="5754" heatid="7872" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                    <SPLIT distance="100" swimtime="00:01:01.62" />
                    <SPLIT distance="150" swimtime="00:01:29.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5727" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5730" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="5732" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="5735" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KUPI" nation="SVK" region="BAO" clubid="6348" name="SPK Kupele Piestany">
          <ATHLETES>
            <ATHLETE birthdate="1987-01-15" firstname="Lucia" gender="F" lastname="Vachanova" nation="SVK" athleteid="6349">
              <RESULTS>
                <RESULT eventid="1173" points="708" reactiontime="+71" swimtime="00:00:34.63" resultid="6350" heatid="7759" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1238" points="738" reactiontime="+86" swimtime="00:01:04.59" resultid="6351" heatid="7804" lane="7" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="637" reactiontime="+75" swimtime="00:01:14.08" resultid="6352" heatid="7931" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="661" reactiontime="+84" swimtime="00:02:24.69" resultid="6353" heatid="7951" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:08.91" />
                    <SPLIT distance="150" swimtime="00:01:46.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="594" reactiontime="+73" swimtime="00:02:42.27" resultid="6354" heatid="8008" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:02.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="660" reactiontime="+85" swimtime="00:05:07.54" resultid="6355" heatid="9048" lane="5" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:47.69" />
                    <SPLIT distance="200" swimtime="00:02:26.80" />
                    <SPLIT distance="250" swimtime="00:03:06.40" />
                    <SPLIT distance="300" swimtime="00:03:46.49" />
                    <SPLIT distance="350" swimtime="00:04:27.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-04-03" firstname="Juraj" gender="M" lastname="Horil" nation="SVK" athleteid="6356">
              <RESULTS>
                <RESULT eventid="1222" points="448" reactiontime="+83" swimtime="00:03:06.71" resultid="6357" heatid="7792" lane="7" entrytime="00:03:09.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                    <SPLIT distance="100" swimtime="00:01:25.98" />
                    <SPLIT distance="150" swimtime="00:02:15.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="378" reactiontime="+76" swimtime="00:01:12.01" resultid="6358" heatid="7812" lane="1" entrytime="00:01:12.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="491" reactiontime="+79" swimtime="00:01:23.17" resultid="6359" heatid="7890" lane="5" entrytime="00:01:24.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="352" reactiontime="+86" swimtime="00:00:35.58" resultid="6360" heatid="7912" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1655" points="507" reactiontime="+79" swimtime="00:00:36.97" resultid="6361" heatid="8040" lane="5" entrytime="00:00:37.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-04-20" firstname="Anna" gender="F" lastname="Kicinova" nation="SVK" athleteid="6362">
              <RESULTS>
                <RESULT eventid="1206" points="575" reactiontime="+94" swimtime="00:03:33.37" resultid="6363" heatid="7781" lane="6" entrytime="00:03:33.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:42.60" />
                    <SPLIT distance="150" swimtime="00:02:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="479" reactiontime="+97" swimtime="00:01:32.75" resultid="6364" heatid="7831" lane="8" entrytime="00:01:31.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="533" reactiontime="+105" swimtime="00:01:38.92" resultid="6365" heatid="7878" lane="7" entrytime="00:01:37.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="379" reactiontime="+98" swimtime="00:03:06.24" resultid="6366" heatid="7947" lane="2" entrytime="00:03:05.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="100" swimtime="00:01:28.06" />
                    <SPLIT distance="150" swimtime="00:02:17.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="537" reactiontime="+86" swimtime="00:00:45.07" resultid="6367" heatid="8025" lane="6" entrytime="00:00:45.40" />
                <RESULT eventid="1687" points="358" reactiontime="+91" swimtime="00:06:43.20" resultid="6368" heatid="9051" lane="5" entrytime="00:06:24.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:01:31.22" />
                    <SPLIT distance="150" swimtime="00:02:22.42" />
                    <SPLIT distance="200" swimtime="00:03:14.59" />
                    <SPLIT distance="250" swimtime="00:04:07.36" />
                    <SPLIT distance="300" swimtime="00:04:59.52" />
                    <SPLIT distance="350" swimtime="00:05:52.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-10-27" firstname="Pavol" gender="M" lastname="Skodny" nation="SVK" athleteid="6369">
              <RESULTS>
                <RESULT eventid="1190" points="496" reactiontime="+71" swimtime="00:00:34.28" resultid="6370" heatid="7774" lane="7" entrytime="00:00:33.30" />
                <RESULT eventid="1286" points="592" reactiontime="+78" swimtime="00:01:11.24" resultid="6371" heatid="7851" lane="2" entrytime="00:01:11.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="530" reactiontime="+75" swimtime="00:01:12.94" resultid="6372" heatid="7940" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="497" reactiontime="+87" swimtime="00:05:42.05" resultid="6373" heatid="8807" lane="4" entrytime="00:05:38.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:01:17.59" />
                    <SPLIT distance="150" swimtime="00:02:01.32" />
                    <SPLIT distance="200" swimtime="00:02:44.52" />
                    <SPLIT distance="250" swimtime="00:03:34.48" />
                    <SPLIT distance="300" swimtime="00:04:24.19" />
                    <SPLIT distance="350" swimtime="00:05:03.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="570" reactiontime="+72" swimtime="00:02:38.52" resultid="6374" heatid="8018" lane="1" entrytime="00:02:37.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                    <SPLIT distance="150" swimtime="00:01:57.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="483" reactiontime="+85" swimtime="00:05:06.54" resultid="6375" heatid="9062" lane="2" entrytime="00:05:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:49.06" />
                    <SPLIT distance="200" swimtime="00:02:28.26" />
                    <SPLIT distance="250" swimtime="00:03:07.78" />
                    <SPLIT distance="300" swimtime="00:03:48.28" />
                    <SPLIT distance="350" swimtime="00:04:28.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SPNI" nation="SVK" region="SSO" clubid="6222" name="SPU Nitra">
          <ATHLETES>
            <ATHLETE birthdate="1947-10-01" firstname="Jozef" gender="M" lastname="Kral" nation="POL" athleteid="6221">
              <RESULTS>
                <RESULT comment="M8 - Przenoszenie ramion do przodu pod powierzchnią wody podczas ostatniego cyklu pracy ramion przed nawrotem lub na zakończenie wyścigu  (Czas: 13:54)" eventid="1318" reactiontime="+102" status="DSQ" swimtime="00:03:31.45" resultid="6223" heatid="7861" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                    <SPLIT distance="100" swimtime="00:01:40.65" />
                    <SPLIT distance="150" swimtime="00:02:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="557" reactiontime="+110" swimtime="00:00:37.14" resultid="6224" heatid="7910" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1591" points="496" reactiontime="+110" swimtime="00:01:30.46" resultid="6225" heatid="7996" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASZC" nation="POL" region="16" clubid="2011" name="STP Masters Szczecinek">
          <ATHLETES>
            <ATHLETE birthdate="1933-02-19" firstname="Zbigniew" gender="M" lastname="Ludwiczak" nation="POL" athleteid="2012">
              <RESULTS>
                <RESULT eventid="1190" points="353" reactiontime="+116" swimtime="00:01:01.82" resultid="2013" heatid="7764" lane="1" entrytime="00:00:57.00" />
                <RESULT eventid="1254" points="360" swimtime="00:01:50.50" resultid="2014" heatid="7807" lane="1" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="410" reactiontime="+117" swimtime="00:02:09.38" resultid="2015" heatid="7933" lane="2" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="426" swimtime="00:03:59.49" resultid="2016" heatid="7952" lane="4" entrytime="00:04:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.20" />
                    <SPLIT distance="100" swimtime="00:01:57.02" />
                    <SPLIT distance="150" swimtime="00:02:59.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="430" reactiontime="+108" swimtime="00:04:38.15" resultid="2017" heatid="8010" lane="5" entrytime="00:04:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.50" />
                    <SPLIT distance="100" swimtime="00:02:16.92" />
                    <SPLIT distance="150" swimtime="00:03:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="454" swimtime="00:08:27.54" resultid="2018" heatid="9070" lane="3" entrytime="00:08:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                    <SPLIT distance="100" swimtime="00:01:57.79" />
                    <SPLIT distance="150" swimtime="00:03:01.68" />
                    <SPLIT distance="200" swimtime="00:04:05.11" />
                    <SPLIT distance="250" swimtime="00:05:09.37" />
                    <SPLIT distance="300" swimtime="00:06:14.58" />
                    <SPLIT distance="350" swimtime="00:07:18.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SAKIE" nation="POL" region="12" clubid="6084" name="Salos Kielce">
          <CONTACT name="Kijewska Iwona" phone="606 760 616" />
          <ATHLETES>
            <ATHLETE birthdate="1970-05-17" firstname="Iwona" gender="F" lastname="Kijewska" nation="POL" athleteid="6097">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="6098" heatid="7676" lane="3" entrytime="00:00:36.81" />
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="6099" heatid="7715" lane="6" entrytime="00:03:15.24" />
                <RESULT eventid="1206" status="DNS" swimtime="00:00:00.00" resultid="6100" heatid="7782" lane="6" entrytime="00:03:20.46" />
                <RESULT eventid="1270" status="DNS" swimtime="00:00:00.00" resultid="6101" heatid="7832" lane="8" entrytime="00:01:28.56" />
                <RESULT eventid="1366" status="DNS" swimtime="00:00:00.00" resultid="6102" heatid="7877" lane="4" entrytime="00:01:38.21" />
                <RESULT eventid="1399" status="DNS" swimtime="00:00:00.00" resultid="6103" heatid="7901" lane="1" entrytime="00:00:39.78" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="6104" heatid="7988" lane="4" entrytime="00:01:35.11" />
                <RESULT eventid="1639" status="DNS" swimtime="00:00:00.00" resultid="6105" heatid="8025" lane="2" entrytime="00:00:45.81" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIGLI" nation="POL" region="11" clubid="2245" name="SiKReT Masters Gliwice">
          <CONTACT city="Gliwice" email="joannaeco@wp.pl" name="Joanna Zagała" phone="601427257" street="Jagielońska 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1962-05-15" firstname="Mietek" gender="M" lastname="Mydłowski" nation="POL" athleteid="2246">
              <RESULTS>
                <RESULT eventid="1076" points="605" reactiontime="+94" swimtime="00:00:30.04" resultid="2247" heatid="7694" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1108" points="525" reactiontime="+87" swimtime="00:02:57.17" resultid="2248" heatid="7727" lane="6" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:15.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="547" reactiontime="+88" swimtime="00:03:09.20" resultid="2249" heatid="7791" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                    <SPLIT distance="100" swimtime="00:01:30.35" />
                    <SPLIT distance="150" swimtime="00:02:20.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="563" reactiontime="+87" swimtime="00:01:19.28" resultid="2250" heatid="7847" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="529" reactiontime="+86" swimtime="00:01:25.95" resultid="2251" heatid="7889" lane="7" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="495" reactiontime="+91" swimtime="00:01:21.95" resultid="2252" heatid="7937" lane="5" entrytime="00:01:21.37" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="2253">
              <RESULTS>
                <RESULT eventid="1092" points="301" reactiontime="+90" swimtime="00:04:15.14" resultid="2254" heatid="7714" lane="2" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.38" />
                    <SPLIT distance="100" swimtime="00:02:12.35" />
                    <SPLIT distance="150" swimtime="00:03:16.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="404" reactiontime="+94" swimtime="00:04:10.47" resultid="2255" heatid="7779" lane="6" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.71" />
                    <SPLIT distance="100" swimtime="00:02:03.75" />
                    <SPLIT distance="150" swimtime="00:03:08.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="305" reactiontime="+91" swimtime="00:01:55.04" resultid="2256" heatid="7828" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="431" reactiontime="+87" swimtime="00:01:50.78" resultid="2257" heatid="7876" lane="8" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="331" reactiontime="+78" swimtime="00:03:40.54" resultid="2258" heatid="7945" lane="8" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                    <SPLIT distance="100" swimtime="00:01:46.72" />
                    <SPLIT distance="150" swimtime="00:02:45.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="240" reactiontime="+77" swimtime="00:02:06.42" resultid="2259" heatid="7987" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="466" reactiontime="+79" swimtime="00:00:48.42" resultid="2260" heatid="8022" lane="4" entrytime="00:00:51.00" />
                <RESULT eventid="1059" points="378" reactiontime="+83" swimtime="00:00:41.81" resultid="3559" heatid="7674" lane="6" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="2261">
              <RESULTS>
                <RESULT eventid="1059" points="380" reactiontime="+72" swimtime="00:00:39.32" resultid="2262" heatid="7673" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1092" points="338" reactiontime="+85" swimtime="00:03:42.94" resultid="2263" heatid="7714" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.62" />
                    <SPLIT distance="100" swimtime="00:01:47.46" />
                    <SPLIT distance="150" swimtime="00:02:50.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="395" reactiontime="+80" swimtime="00:04:01.76" resultid="2264" heatid="7779" lane="3" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.22" />
                    <SPLIT distance="100" swimtime="00:01:56.82" />
                    <SPLIT distance="150" swimtime="00:03:00.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="364" reactiontime="+77" swimtime="00:01:41.62" resultid="2265" heatid="7828" lane="4" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="383" reactiontime="+77" swimtime="00:01:50.43" resultid="2266" heatid="7875" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="307" reactiontime="+77" swimtime="00:03:19.92" resultid="2267" heatid="7945" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                    <SPLIT distance="100" swimtime="00:01:36.92" />
                    <SPLIT distance="150" swimtime="00:02:30.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="313" reactiontime="+86" swimtime="00:03:51.87" resultid="2268" heatid="8005" lane="5" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.13" />
                    <SPLIT distance="100" swimtime="00:02:55.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="408" reactiontime="+71" swimtime="00:00:49.38" resultid="2269" heatid="8022" lane="8" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIWAR" nation="POL" region="14" clubid="5120" name="Sinnet Warszawa">
          <CONTACT email="piotrbarski@uw.edu.pl" name="barski" />
          <ATHLETES>
            <ATHLETE birthdate="1965-02-17" firstname="Piotr" gender="M" lastname="Barski" nation="POL" athleteid="5121">
              <RESULTS>
                <RESULT eventid="1076" points="802" reactiontime="+78" swimtime="00:00:26.02" resultid="5122" heatid="7710" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1222" points="787" reactiontime="+82" swimtime="00:02:41.63" resultid="5123" heatid="7789" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                    <SPLIT distance="100" swimtime="00:01:17.72" />
                    <SPLIT distance="150" swimtime="00:02:00.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="796" reactiontime="+82" swimtime="00:00:57.09" resultid="5124" heatid="7824" lane="8" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="779" reactiontime="+84" swimtime="00:01:13.05" resultid="5125" heatid="7895" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="5126" heatid="7967" lane="8" entrytime="00:02:08.00" />
                <RESULT eventid="1655" points="879" reactiontime="+79" swimtime="00:00:32.02" resultid="5127" heatid="8047" lane="2" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-25" firstname="Agnieszka" gender="F" lastname="Besler" nation="POL" athleteid="5128">
              <RESULTS>
                <RESULT eventid="1059" points="601" reactiontime="+101" swimtime="00:00:32.18" resultid="5129" heatid="7681" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1206" points="504" reactiontime="+82" swimtime="00:03:24.45" resultid="5130" heatid="7782" lane="8" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                    <SPLIT distance="100" swimtime="00:01:35.97" />
                    <SPLIT distance="150" swimtime="00:02:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="504" reactiontime="+78" swimtime="00:01:32.74" resultid="5131" heatid="7878" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="473" reactiontime="+82" swimtime="00:00:43.49" resultid="5132" heatid="8026" lane="6" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="FIWAR" nation="POL" region="14" clubid="6106" name="Sport Figielski Warszawa">
          <CONTACT city="Warszawa" email="grzegorz.figielski@sport-figielski.pl" fax="224032788" internet="www.sport-figielski.pl" name="Grzegorz Figielski" phone="501294477" state="MAZ" street="Sarmacka 21 m. 41" zip="02-972" />
          <ATHLETES>
            <ATHLETE birthdate="1959-04-28" firstname="Joanna" gender="F" lastname="Szczepańska" nation="POL" athleteid="6107">
              <RESULTS>
                <RESULT eventid="1140" points="150" swimtime="00:18:19.83" resultid="6108" heatid="8715" lane="2" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                    <SPLIT distance="100" swimtime="00:01:58.12" />
                    <SPLIT distance="200" swimtime="00:04:17.49" />
                    <SPLIT distance="300" swimtime="00:06:25.83" />
                    <SPLIT distance="400" swimtime="00:08:56.11" />
                    <SPLIT distance="500" swimtime="00:11:18.97" />
                    <SPLIT distance="600" swimtime="00:13:38.91" />
                    <SPLIT distance="700" swimtime="00:16:06.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-03-04" firstname="Wiktor" gender="M" lastname="Dębski" nation="POL" athleteid="6111">
              <RESULTS>
                <RESULT eventid="1076" points="665" reactiontime="+87" swimtime="00:00:27.21" resultid="6112" heatid="7698" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1286" points="660" reactiontime="+90" swimtime="00:01:08.68" resultid="6113" heatid="7848" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="6114" heatid="7890" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="1415" points="598" reactiontime="+88" swimtime="00:00:29.82" resultid="6115" heatid="7916" lane="1" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SBKRA" nation="POL" region="06" clubid="6273" name="Sport and Body Kraków">
          <ATHLETES>
            <ATHLETE birthdate="1987-12-13" firstname="Mateusz" gender="M" lastname="Miłek" nation="POL" athleteid="6272">
              <RESULTS>
                <RESULT eventid="1076" points="711" reactiontime="+70" swimtime="00:00:25.58" resultid="6274" heatid="7709" lane="5" entrytime="00:00:26.20" />
                <RESULT eventid="1108" points="576" reactiontime="+65" swimtime="00:02:24.86" resultid="6275" heatid="7729" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="100" swimtime="00:01:09.06" />
                    <SPLIT distance="150" swimtime="00:01:51.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="669" reactiontime="+55" swimtime="00:00:28.64" resultid="6276" heatid="7777" lane="1" entrytime="00:00:29.90" />
                <RESULT eventid="1318" points="588" reactiontime="+67" swimtime="00:02:31.91" resultid="6277" heatid="7865" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:52.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="690" reactiontime="+71" swimtime="00:00:26.82" resultid="6278" heatid="7923" lane="7" entrytime="00:00:27.90" />
                <RESULT eventid="1447" points="649" reactiontime="+62" swimtime="00:01:03.54" resultid="6279" heatid="7941" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="691" reactiontime="+69" swimtime="00:01:01.00" resultid="6280" heatid="8001" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="564" reactiontime="+71" swimtime="00:00:34.20" resultid="6281" heatid="8041" lane="5" entrytime="00:00:36.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SQOST" nation="POL" region="14" clubid="6142" name="Squatina Ostrołęka">
          <CONTACT city="Ostrołęka" email="biezunskamaja@gmail.com" name="Bieżuńska Maja" phone="666-353-028" state="MAZ" street="ul. Łęczysk 10/14/26" zip="07-410" />
          <ATHLETES>
            <ATHLETE birthdate="1979-06-26" firstname="Maja" gender="F" lastname="Bieżuńska" nation="POL" athleteid="6164">
              <RESULTS>
                <RESULT eventid="1639" points="567" reactiontime="+84" swimtime="00:00:38.36" resultid="6165" heatid="8028" lane="3" entrytime="00:00:36.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWWAR" nation="POL" region="14" clubid="5546" name="St. Pływackie Swimmers Warszawa" shortname="Swimmers Warszawa">
          <CONTACT city="WARSZAWA" email="remog@swimmersteam.pl" internet="www.swimmersteam.pl" name="GOŁĘBIOWSKI" phone="601333782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1976-07-07" firstname="Remigiusz" gender="M" lastname="Gołębiowski" nation="POL" athleteid="5554">
              <RESULTS>
                <RESULT eventid="1156" points="756" reactiontime="+94" swimtime="00:18:28.81" resultid="5555" heatid="8717" lane="5" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:06.91" />
                    <SPLIT distance="150" swimtime="00:01:42.54" />
                    <SPLIT distance="200" swimtime="00:02:18.66" />
                    <SPLIT distance="250" swimtime="00:02:55.20" />
                    <SPLIT distance="300" swimtime="00:03:31.62" />
                    <SPLIT distance="350" swimtime="00:04:07.96" />
                    <SPLIT distance="400" swimtime="00:04:44.79" />
                    <SPLIT distance="450" swimtime="00:05:21.37" />
                    <SPLIT distance="500" swimtime="00:05:57.81" />
                    <SPLIT distance="550" swimtime="00:06:34.80" />
                    <SPLIT distance="600" swimtime="00:07:11.93" />
                    <SPLIT distance="650" swimtime="00:07:48.94" />
                    <SPLIT distance="700" swimtime="00:08:26.40" />
                    <SPLIT distance="750" swimtime="00:09:03.98" />
                    <SPLIT distance="800" swimtime="00:09:41.82" />
                    <SPLIT distance="850" swimtime="00:10:19.86" />
                    <SPLIT distance="900" swimtime="00:10:57.76" />
                    <SPLIT distance="950" swimtime="00:11:35.66" />
                    <SPLIT distance="1000" swimtime="00:12:13.77" />
                    <SPLIT distance="1050" swimtime="00:12:51.19" />
                    <SPLIT distance="1100" swimtime="00:13:28.82" />
                    <SPLIT distance="1150" swimtime="00:14:06.52" />
                    <SPLIT distance="1200" swimtime="00:14:44.24" />
                    <SPLIT distance="1250" swimtime="00:15:21.97" />
                    <SPLIT distance="1300" swimtime="00:15:59.60" />
                    <SPLIT distance="1350" swimtime="00:16:37.63" />
                    <SPLIT distance="1400" swimtime="00:17:15.02" />
                    <SPLIT distance="1450" swimtime="00:17:52.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="768" reactiontime="+83" swimtime="00:00:28.01" resultid="5556" heatid="7924" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1479" points="664" reactiontime="+84" swimtime="00:02:07.71" resultid="5557" heatid="7967" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                    <SPLIT distance="100" swimtime="00:01:00.45" />
                    <SPLIT distance="150" swimtime="00:01:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="748" reactiontime="+74" swimtime="00:01:02.62" resultid="5558" heatid="8002" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="668" reactiontime="+83" swimtime="00:04:37.15" resultid="5559" heatid="9059" lane="5" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:04.70" />
                    <SPLIT distance="150" swimtime="00:01:39.71" />
                    <SPLIT distance="200" swimtime="00:02:15.36" />
                    <SPLIT distance="250" swimtime="00:02:50.94" />
                    <SPLIT distance="300" swimtime="00:03:26.73" />
                    <SPLIT distance="350" swimtime="00:04:02.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-03" firstname="Bolesław" gender="M" lastname="Porolniczak" nation="POL" athleteid="5560">
              <RESULTS>
                <RESULT eventid="1076" points="570" reactiontime="+88" swimtime="00:00:26.69" resultid="5561" heatid="7708" lane="4" entrytime="00:00:26.50" />
                <RESULT eventid="1254" points="512" reactiontime="+85" swimtime="00:01:01.28" resultid="5562" heatid="7821" lane="6" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="5563" heatid="7920" lane="8" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STPOZ" nation="POL" region="15" clubid="3575" name="Start Poznań">
          <ATHLETES>
            <ATHLETE birthdate="1969-02-26" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="3574">
              <RESULTS>
                <RESULT eventid="1076" points="684" reactiontime="+83" swimtime="00:00:26.96" resultid="3576" heatid="7707" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1254" points="661" reactiontime="+85" swimtime="00:00:59.76" resultid="3577" heatid="7816" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="635" reactiontime="+85" swimtime="00:01:09.58" resultid="3578" heatid="7852" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="619" reactiontime="+79" swimtime="00:01:09.27" resultid="3579" heatid="7940" lane="3" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="685" reactiontime="+76" swimtime="00:02:29.16" resultid="3580" heatid="8018" lane="4" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:12.42" />
                    <SPLIT distance="150" swimtime="00:01:50.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-02" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="6190">
              <RESULTS>
                <RESULT eventid="1076" points="747" reactiontime="+73" swimtime="00:00:26.64" resultid="6191" heatid="7708" lane="1" entrytime="00:00:26.80" />
                <RESULT eventid="1108" points="776" reactiontime="+77" swimtime="00:02:28.63" resultid="6192" heatid="7731" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:10.62" />
                    <SPLIT distance="150" swimtime="00:01:54.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="791" reactiontime="+66" swimtime="00:00:57.22" resultid="6193" heatid="7823" lane="2" entrytime="00:00:58.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="720" reactiontime="+73" swimtime="00:01:07.48" resultid="6194" heatid="7853" lane="3" entrytime="00:01:07.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="694" reactiontime="+73" swimtime="00:02:09.57" resultid="6195" heatid="7953" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                    <SPLIT distance="150" swimtime="00:01:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K4 - Cykl ruchowy inny niż jeden ruch ramion i jedno kopnięcie nogami  (Czas: 21:31)" eventid="1543" reactiontime="+84" status="DSQ" swimtime="00:05:24.48" resultid="6196" heatid="8806" lane="7" entrytime="00:05:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:13.40" />
                    <SPLIT distance="150" swimtime="00:01:55.03" />
                    <SPLIT distance="200" swimtime="00:02:36.77" />
                    <SPLIT distance="250" swimtime="00:03:24.60" />
                    <SPLIT distance="300" swimtime="00:04:13.24" />
                    <SPLIT distance="350" swimtime="00:04:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="654" reactiontime="+76" swimtime="00:04:43.26" resultid="6197" heatid="9060" lane="5" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:09.01" />
                    <SPLIT distance="150" swimtime="00:01:44.88" />
                    <SPLIT distance="200" swimtime="00:02:21.29" />
                    <SPLIT distance="250" swimtime="00:02:57.34" />
                    <SPLIT distance="300" swimtime="00:03:33.12" />
                    <SPLIT distance="350" swimtime="00:04:08.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STWRO" nation="POL" region="01" clubid="2889" name="Start Wrocław">
          <CONTACT city="Wrocław" email="WZSSTART@POST.PL" fax="0713437281" internet="www.start.wroclaw.pl" name="Sajdel" phone="0713430231" state="DOL" street="Notecka 12" zip="54-128" />
          <ATHLETES>
            <ATHLETE birthdate="1974-04-30" firstname="Sebastian" gender="M" lastname="Szymański" nation="POL" athleteid="2913">
              <RESULTS>
                <RESULT eventid="1076" points="620" reactiontime="+95" swimtime="00:00:27.81" resultid="2914" heatid="7703" lane="7" entrytime="00:00:28.05" entrycourse="SCM" />
                <RESULT eventid="1190" points="527" reactiontime="+83" swimtime="00:00:33.60" resultid="2915" heatid="7773" lane="1" entrytime="00:00:34.34" entrycourse="SCM" />
                <RESULT eventid="1254" points="594" reactiontime="+94" swimtime="00:01:01.18" resultid="2916" heatid="7820" lane="2" entrytime="00:01:01.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="657" reactiontime="+97" swimtime="00:00:29.51" resultid="2917" heatid="7920" lane="7" entrytime="00:00:29.88" entrycourse="SCM" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="2918" heatid="7962" lane="4" entrytime="00:02:22.22" entrycourse="SCM" />
                <RESULT eventid="1591" points="594" reactiontime="+99" swimtime="00:01:07.63" resultid="2919" heatid="7999" lane="4" entrytime="00:01:10.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWTAK" nation="LTU" clubid="4636" name="Swimming Masters Club Takas Kaunas" shortname="SMC Takas Kaunas">
          <CONTACT city="Kaunas" email="abicka@takas.lt" internet="www.klubastakas.lt" name="Romaldas Bickauskas" phone="+37068687934" street="Lentvario g. 19-1" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1964-10-18" firstname="Ramune" gender="F" lastname="Ivanauskaite" nation="LTU" athleteid="4650">
              <RESULTS>
                <RESULT eventid="1092" points="485" reactiontime="+84" swimtime="00:03:14.63" resultid="4651" heatid="7715" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                    <SPLIT distance="100" swimtime="00:01:32.03" />
                    <SPLIT distance="150" swimtime="00:02:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="426" reactiontime="+85" swimtime="00:01:20.23" resultid="4652" heatid="7802" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="490" reactiontime="+95" swimtime="00:01:29.96" resultid="4653" heatid="7928" lane="6" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="439" reactiontime="+90" swimtime="00:02:55.86" resultid="4654" heatid="7948" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                    <SPLIT distance="150" swimtime="00:02:11.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="509" reactiontime="+90" swimtime="00:03:12.46" resultid="4655" heatid="8007" lane="3" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                    <SPLIT distance="100" swimtime="00:01:34.41" />
                    <SPLIT distance="150" swimtime="00:02:23.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-12-26" firstname="Arlandas Antanas" gender="M" lastname="Juodeska" nation="LTU" athleteid="4656">
              <RESULTS>
                <RESULT eventid="1076" points="702" reactiontime="+76" swimtime="00:00:28.58" resultid="4657" heatid="7701" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1190" points="700" reactiontime="+64" swimtime="00:00:33.08" resultid="4658" heatid="7773" lane="2" entrytime="00:00:34.06" />
                <RESULT eventid="1222" points="600" reactiontime="+81" swimtime="00:03:03.45" resultid="4659" heatid="7792" lane="2" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:28.78" />
                    <SPLIT distance="150" swimtime="00:02:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="4660" heatid="7849" lane="2" entrytime="00:01:14.57" />
                <RESULT eventid="1383" points="631" reactiontime="+79" swimtime="00:01:21.06" resultid="4661" heatid="7891" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="657" reactiontime="+71" swimtime="00:01:14.58" resultid="4662" heatid="7939" lane="5" entrytime="00:01:14.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="4663" heatid="8017" lane="2" entrytime="00:02:42.00" />
                <RESULT eventid="1655" points="690" reactiontime="+79" swimtime="00:00:35.51" resultid="4664" heatid="8043" lane="8" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-06-18" firstname="Linas" gender="M" lastname="Kersevicius" nation="LTU" athleteid="4665">
              <RESULTS>
                <RESULT eventid="1076" points="614" reactiontime="+81" swimtime="00:00:27.95" resultid="4666" heatid="7704" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="1190" points="683" reactiontime="+74" swimtime="00:00:30.82" resultid="4667" heatid="7775" lane="3" entrytime="00:00:30.80" />
                <RESULT eventid="1447" points="699" reactiontime="+73" swimtime="00:01:06.53" resultid="4668" heatid="7942" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="730" reactiontime="+80" swimtime="00:02:26.00" resultid="4669" heatid="8019" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:47.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-04-12" firstname="Aleksandra" gender="F" lastname="Yliene" nation="LTU" athleteid="4670">
              <RESULTS>
                <RESULT eventid="1059" points="420" reactiontime="+99" swimtime="00:00:43.04" resultid="4671" heatid="7674" lane="1" entrytime="00:00:43.50" />
                <RESULT eventid="1173" points="506" reactiontime="+83" swimtime="00:00:50.22" resultid="4672" heatid="7755" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1238" points="364" reactiontime="+121" swimtime="00:01:39.32" resultid="4673" heatid="7798" lane="1" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="431" reactiontime="+82" swimtime="00:01:57.52" resultid="4674" heatid="7927" lane="1" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="374" reactiontime="+79" swimtime="00:04:21.40" resultid="4675" heatid="8005" lane="6" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.07" />
                    <SPLIT distance="100" swimtime="00:02:03.47" />
                    <SPLIT distance="150" swimtime="00:03:14.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMSZC" nation="POL" region="16" clubid="2050" name="Swimming Masters Team Szczecin">
          <CONTACT email="teczowy.dyndol@gmail.com" name="Brodacki Maciej" phone="608396939" />
          <ATHLETES>
            <ATHLETE birthdate="1987-02-27" firstname="Szymon" gender="M" lastname="Kluczyk" nation="POL" athleteid="2051">
              <RESULTS>
                <RESULT eventid="1108" points="559" reactiontime="+86" swimtime="00:02:26.30" resultid="2052" heatid="7731" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:51.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="657" reactiontime="+95" swimtime="00:05:13.89" resultid="2053" heatid="8806" lane="8" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:11.45" />
                    <SPLIT distance="150" swimtime="00:01:52.10" />
                    <SPLIT distance="200" swimtime="00:02:32.27" />
                    <SPLIT distance="250" swimtime="00:03:17.82" />
                    <SPLIT distance="300" swimtime="00:04:03.59" />
                    <SPLIT distance="350" swimtime="00:04:39.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="715" reactiontime="+90" swimtime="00:04:33.30" resultid="2054" heatid="9061" lane="3" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:05.13" />
                    <SPLIT distance="150" swimtime="00:01:39.34" />
                    <SPLIT distance="200" swimtime="00:02:13.98" />
                    <SPLIT distance="250" swimtime="00:02:48.77" />
                    <SPLIT distance="300" swimtime="00:03:23.76" />
                    <SPLIT distance="350" swimtime="00:03:58.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="Roenig" nation="POL" athleteid="2055">
              <RESULTS>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="2056" heatid="7848" lane="6" entrytime="00:01:15.00" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="2057" heatid="7893" lane="6" entrytime="00:01:18.00" />
                <RESULT eventid="1415" points="134" swimtime="00:00:46.29" resultid="2058" heatid="7919" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="2059" heatid="8044" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-04-17" firstname="Alicja" gender="F" lastname="Nowak" nation="POL" athleteid="2060">
              <RESULTS>
                <RESULT eventid="1059" points="672" reactiontime="+81" swimtime="00:00:30.22" resultid="2061" heatid="7682" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1173" points="689" reactiontime="+70" swimtime="00:00:34.29" resultid="2062" heatid="7761" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1270" points="656" reactiontime="+84" swimtime="00:01:14.92" resultid="2063" heatid="7836" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="715" reactiontime="+80" swimtime="00:00:32.01" resultid="2064" heatid="7905" lane="7" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="Brodacki" nation="POL" athleteid="2065">
              <RESULTS>
                <RESULT eventid="1076" points="666" reactiontime="+75" swimtime="00:00:25.34" resultid="2066" heatid="7710" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1108" points="540" reactiontime="+77" swimtime="00:02:25.00" resultid="2067" heatid="7730" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:51.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="677" reactiontime="+80" swimtime="00:00:55.85" resultid="2068" heatid="7823" lane="4" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="607" reactiontime="+80" swimtime="00:01:04.95" resultid="2069" heatid="7853" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="478" reactiontime="+81" swimtime="00:00:29.25" resultid="2070" heatid="7919" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1479" points="587" reactiontime="+84" swimtime="00:02:07.21" resultid="2071" heatid="7964" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                    <SPLIT distance="100" swimtime="00:01:00.02" />
                    <SPLIT distance="150" swimtime="00:01:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="607" reactiontime="+83" swimtime="00:04:43.68" resultid="2072" heatid="9061" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:06.80" />
                    <SPLIT distance="150" swimtime="00:01:42.71" />
                    <SPLIT distance="200" swimtime="00:02:18.54" />
                    <SPLIT distance="250" swimtime="00:02:54.26" />
                    <SPLIT distance="300" swimtime="00:03:31.28" />
                    <SPLIT distance="350" swimtime="00:04:08.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-27" firstname="Rafał" gender="M" lastname="Lisiecki" nation="POL" athleteid="2073">
              <RESULTS>
                <RESULT eventid="1076" points="601" reactiontime="+84" swimtime="00:00:27.06" resultid="2074" heatid="7707" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="1190" points="538" reactiontime="+73" swimtime="00:00:30.79" resultid="2075" heatid="7775" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="1447" points="541" reactiontime="+70" swimtime="00:01:07.51" resultid="2076" heatid="7941" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1357" status="WDR" swimtime="00:00:00.00" resultid="2077" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2073" number="1" />
                    <RELAYPOSITION athleteid="2055" number="2" />
                    <RELAYPOSITION athleteid="2051" number="3" />
                    <RELAYPOSITION athleteid="2065" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" status="WDR" swimtime="00:00:00.00" resultid="2078" entrytime="00:01:53.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2051" number="1" />
                    <RELAYPOSITION athleteid="2065" number="2" />
                    <RELAYPOSITION athleteid="2073" number="3" />
                    <RELAYPOSITION athleteid="2055" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TKKOS" nation="POL" region="16" clubid="4676" name="TKKF Koszalin">
          <CONTACT email="jakubkielar3@gmail.com" internet="www.k-swim.pl" name="Kielar Jakub" phone="693193137" />
          <ATHLETES>
            <ATHLETE birthdate="1988-02-16" firstname="Katarzyna" gender="F" lastname="Gudaniec" nation="POL" athleteid="4677">
              <RESULTS>
                <RESULT eventid="1463" points="567" reactiontime="+81" swimtime="00:02:32.30" resultid="4678" heatid="7950" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                    <SPLIT distance="150" swimtime="00:01:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="571" reactiontime="+83" swimtime="00:05:22.75" resultid="4679" heatid="9047" lane="1" entrytime="00:05:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:13.36" />
                    <SPLIT distance="150" swimtime="00:01:54.17" />
                    <SPLIT distance="200" swimtime="00:02:35.39" />
                    <SPLIT distance="250" swimtime="00:03:17.82" />
                    <SPLIT distance="300" swimtime="00:03:59.99" />
                    <SPLIT distance="350" swimtime="00:04:41.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-08-28" firstname="Dorota" gender="F" lastname="Gudaniec" nation="POL" athleteid="4680">
              <RESULTS>
                <RESULT eventid="1140" points="402" swimtime="00:13:12.80" resultid="4681" heatid="8714" lane="1" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                    <SPLIT distance="100" swimtime="00:01:28.98" />
                    <SPLIT distance="200" swimtime="00:03:09.02" />
                    <SPLIT distance="300" swimtime="00:04:50.05" />
                    <SPLIT distance="400" swimtime="00:06:31.19" />
                    <SPLIT distance="500" swimtime="00:08:12.46" />
                    <SPLIT distance="600" swimtime="00:09:53.66" />
                    <SPLIT distance="700" swimtime="00:11:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="499" reactiontime="+99" swimtime="00:03:43.77" resultid="4682" heatid="7781" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.76" />
                    <SPLIT distance="100" swimtime="00:01:45.58" />
                    <SPLIT distance="150" swimtime="00:02:44.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="478" reactiontime="+102" swimtime="00:01:32.87" resultid="4683" heatid="7830" lane="3" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="477" reactiontime="+106" swimtime="00:01:42.64" resultid="4684" heatid="7877" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" status="DNS" swimtime="00:00:00.00" resultid="4685" heatid="8803" lane="4" entrytime="00:07:10.00" />
                <RESULT eventid="1687" points="412" reactiontime="+101" swimtime="00:06:24.74" resultid="4686" heatid="9051" lane="4" entrytime="00:06:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:27.56" />
                    <SPLIT distance="150" swimtime="00:02:16.57" />
                    <SPLIT distance="200" swimtime="00:03:06.42" />
                    <SPLIT distance="250" swimtime="00:03:56.82" />
                    <SPLIT distance="300" swimtime="00:04:46.80" />
                    <SPLIT distance="350" swimtime="00:05:36.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-02-03" firstname="Andrzej" gender="M" lastname="Michałkowski" nation="POL" athleteid="4687">
              <RESULTS>
                <RESULT eventid="1076" points="320" reactiontime="+95" swimtime="00:00:39.46" resultid="4688" heatid="7702" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="1286" points="364" reactiontime="+95" swimtime="00:01:41.39" resultid="4689" heatid="7840" lane="4" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="493" reactiontime="+115" swimtime="00:01:38.87" resultid="4690" heatid="7885" lane="7" entrytime="00:01:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="261" reactiontime="+111" swimtime="00:03:35.48" resultid="4691" heatid="7953" lane="2" entrytime="00:03:41.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.37" />
                    <SPLIT distance="100" swimtime="00:01:40.56" />
                    <SPLIT distance="150" swimtime="00:02:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="566" reactiontime="+97" swimtime="00:00:40.85" resultid="4692" heatid="8035" lane="7" entrytime="00:00:42.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-06" firstname="Joanna" gender="F" lastname="Stankiewicz-Majkowska" nation="POL" athleteid="4693">
              <RESULTS>
                <RESULT eventid="1059" points="328" reactiontime="+105" swimtime="00:00:39.39" resultid="4694" heatid="7675" lane="6" entrytime="00:00:39.38" />
                <RESULT eventid="1173" points="324" reactiontime="+80" swimtime="00:00:46.03" resultid="4695" heatid="7755" lane="5" entrytime="00:00:47.40" />
                <RESULT eventid="1270" points="347" reactiontime="+102" swimtime="00:01:36.95" resultid="4696" heatid="7829" lane="2" entrytime="00:01:39.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="387" reactiontime="+105" swimtime="00:01:43.84" resultid="4697" heatid="7877" lane="1" entrytime="00:01:44.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="354" reactiontime="+112" swimtime="00:00:48.51" resultid="4698" heatid="8024" lane="8" entrytime="00:00:49.06" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-07-05" firstname="Krzysztof" gender="M" lastname="Stefański" nation="POL" athleteid="4699">
              <RESULTS>
                <RESULT eventid="1076" points="578" reactiontime="+74" swimtime="00:00:28.52" resultid="4700" heatid="7701" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1254" points="505" reactiontime="+91" swimtime="00:01:05.37" resultid="4701" heatid="7816" lane="5" entrytime="00:01:05.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="422" reactiontime="+87" swimtime="00:00:33.48" resultid="4702" heatid="7915" lane="1" entrytime="00:00:33.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-21" firstname="Jakub" gender="M" lastname="Kielar" nation="POL" athleteid="4703">
              <RESULTS>
                <RESULT eventid="1076" points="623" reactiontime="+80" swimtime="00:00:27.77" resultid="4704" heatid="7708" lane="8" entrytime="00:00:26.94" />
                <RESULT eventid="1254" points="575" reactiontime="+85" swimtime="00:01:01.84" resultid="4705" heatid="7806" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.30" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G8 - Ukończenie wyścigu nie w położeniu na plecach  (Czas: 13:22)" eventid="1286" reactiontime="+83" status="DSQ" swimtime="00:01:11.74" resultid="4706" heatid="7853" lane="6" entrytime="00:01:07.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="662" reactiontime="+82" swimtime="00:00:29.43" resultid="4707" heatid="7921" lane="1" entrytime="00:00:29.47" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="4708" heatid="7966" lane="5" entrytime="00:02:09.00" />
                <RESULT eventid="1623" points="492" reactiontime="+71" swimtime="00:02:44.63" resultid="4709" heatid="8017" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:18.48" />
                    <SPLIT distance="150" swimtime="00:02:02.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="4710" entrytime="00:04:49.70" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="TKKF Koszalin C" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+89" swimtime="00:02:18.34" resultid="4711" heatid="7735" lane="4" entrytime="00:02:12.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:17.03" />
                    <SPLIT distance="150" swimtime="00:01:49.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4693" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="4687" number="2" reactiontime="+5" />
                    <RELAYPOSITION athleteid="4677" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4699" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" reactiontime="+85" swimtime="00:02:29.47" resultid="4712" heatid="8050" lane="3" entrytime="00:02:33.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:32.13" />
                    <SPLIT distance="150" swimtime="00:02:01.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4680" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="4693" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="4703" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4699" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00607" nation="POL" region="07" clubid="4445" name="TP Masters Opole" shortname="Masters Opole">
          <CONTACT email="opolbud@onet.eu" name="KRASNODĘBSKI" phone="694402057" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Janusz" gender="M" lastname="Garbarczuk" nation="POL" athleteid="4446">
              <RESULTS>
                <RESULT eventid="1076" points="376" reactiontime="+90" swimtime="00:00:37.38" resultid="4447" heatid="7688" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1190" points="324" reactiontime="+94" swimtime="00:00:48.22" resultid="4448" heatid="7768" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1447" points="294" reactiontime="+73" swimtime="00:01:49.32" resultid="4449" heatid="7935" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="315" reactiontime="+70" swimtime="00:04:03.07" resultid="4450" heatid="8011" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.99" />
                    <SPLIT distance="100" swimtime="00:01:56.30" />
                    <SPLIT distance="150" swimtime="00:02:59.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Witkowski" nation="POL" athleteid="4451">
              <RESULTS>
                <RESULT eventid="1076" points="751" reactiontime="+107" swimtime="00:00:35.19" resultid="4452" heatid="7689" lane="1" entrytime="00:00:35.50" />
                <RESULT eventid="1108" points="412" reactiontime="+113" swimtime="00:04:15.23" resultid="4453" heatid="7720" lane="2" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.30" />
                    <SPLIT distance="100" swimtime="00:02:08.46" />
                    <SPLIT distance="150" swimtime="00:03:28.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="591" reactiontime="+89" swimtime="00:00:47.53" resultid="4454" heatid="7765" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1254" points="598" reactiontime="+117" swimtime="00:01:25.57" resultid="4455" heatid="7808" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="262" reactiontime="+116" swimtime="00:00:58.05" resultid="4456" heatid="7906" lane="5" entrytime="00:00:58.00" />
                <RESULT eventid="1447" points="621" reactiontime="+72" swimtime="00:01:47.11" resultid="4457" heatid="7934" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="547" reactiontime="+97" swimtime="00:04:01.35" resultid="4458" heatid="8011" lane="3" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.37" />
                    <SPLIT distance="150" swimtime="00:03:00.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="478" reactiontime="+112" swimtime="00:00:50.11" resultid="4459" heatid="8031" lane="6" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Roman" gender="M" lastname="Birecki" nation="POL" athleteid="4460">
              <RESULTS>
                <RESULT eventid="1076" points="575" reactiontime="+92" swimtime="00:00:31.35" resultid="4461" heatid="7691" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="4462" heatid="8722" lane="8" entrytime="00:26:54.00" />
                <RESULT eventid="1190" points="533" reactiontime="+75" swimtime="00:00:38.80" resultid="4463" heatid="7768" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1318" points="478" reactiontime="+99" swimtime="00:03:08.72" resultid="4464" heatid="7863" lane="8" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:01:28.76" />
                    <SPLIT distance="150" swimtime="00:02:19.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="482" reactiontime="+93" swimtime="00:00:36.37" resultid="4465" heatid="7912" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1479" points="570" reactiontime="+96" swimtime="00:02:40.80" resultid="4466" heatid="7959" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:15.64" />
                    <SPLIT distance="150" swimtime="00:01:58.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="484" reactiontime="+98" swimtime="00:01:22.46" resultid="4467" heatid="7995" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="4468">
              <RESULTS>
                <RESULT eventid="1076" points="787" reactiontime="+80" swimtime="00:00:27.52" resultid="4469" heatid="7698" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1190" points="809" reactiontime="+68" swimtime="00:00:31.52" resultid="4470" heatid="7775" lane="7" entrytime="00:00:31.20" />
                <RESULT eventid="1254" points="816" reactiontime="+87" swimtime="00:01:00.38" resultid="4471" heatid="7817" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="794" reactiontime="+80" swimtime="00:00:29.75" resultid="4472" heatid="7918" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1447" points="830" reactiontime="+63" swimtime="00:01:08.99" resultid="4473" heatid="7941" lane="1" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="859" reactiontime="+68" swimtime="00:02:32.47" resultid="4474" heatid="8018" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                    <SPLIT distance="150" swimtime="00:01:52.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Jan" gender="M" lastname="Bryniak" nation="POL" athleteid="4475">
              <RESULTS>
                <RESULT eventid="1222" points="664" reactiontime="+99" swimtime="00:03:20.50" resultid="4476" heatid="7788" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:36.04" />
                    <SPLIT distance="150" swimtime="00:02:28.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="478" reactiontime="+105" swimtime="00:03:24.24" resultid="4477" heatid="7861" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                    <SPLIT distance="100" swimtime="00:01:36.22" />
                    <SPLIT distance="150" swimtime="00:02:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="635" reactiontime="+100" swimtime="00:01:30.91" resultid="4478" heatid="7884" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="575" reactiontime="+97" swimtime="00:06:59.45" resultid="4479" heatid="8811" lane="6" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="100" swimtime="00:01:35.54" />
                    <SPLIT distance="150" swimtime="00:02:32.62" />
                    <SPLIT distance="200" swimtime="00:03:30.23" />
                    <SPLIT distance="250" swimtime="00:04:24.42" />
                    <SPLIT distance="300" swimtime="00:05:19.77" />
                    <SPLIT distance="350" swimtime="00:06:09.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="408" reactiontime="+102" swimtime="00:01:32.08" resultid="4480" heatid="7995" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="545" reactiontime="+104" swimtime="00:00:41.38" resultid="4481" heatid="8033" lane="7" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Jerzy" gender="M" lastname="Minkiewicz" nation="POL" athleteid="4482">
              <RESULTS>
                <RESULT eventid="1076" points="589" reactiontime="+86" swimtime="00:00:31.11" resultid="4483" heatid="7695" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1108" points="457" reactiontime="+97" swimtime="00:03:12.33" resultid="4484" heatid="7724" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:30.96" />
                    <SPLIT distance="150" swimtime="00:02:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="549" reactiontime="+100" swimtime="00:01:10.83" resultid="4485" heatid="7814" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="534" reactiontime="+95" swimtime="00:01:25.24" resultid="4486" heatid="7843" lane="6" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="467" reactiontime="+102" swimtime="00:00:36.74" resultid="4487" heatid="7912" lane="5" entrytime="00:00:35.50" />
                <RESULT eventid="1479" points="474" reactiontime="+104" swimtime="00:02:50.91" resultid="4488" heatid="7957" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:19.69" />
                    <SPLIT distance="150" swimtime="00:02:05.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="462" reactiontime="+81" swimtime="00:03:20.48" resultid="4489" heatid="8013" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.13" />
                    <SPLIT distance="100" swimtime="00:01:37.94" />
                    <SPLIT distance="150" swimtime="00:02:31.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Oskar" gender="M" lastname="Orski" nation="POL" athleteid="4490">
              <RESULTS>
                <RESULT eventid="1076" points="547" reactiontime="+105" swimtime="00:00:29.55" resultid="4491" heatid="7699" lane="6" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1933-01-01" firstname="Bronisław" gender="M" lastname="Pichurski" nation="POL" athleteid="4492">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4493" heatid="7684" lane="3" entrytime="00:01:30.00" />
                <RESULT eventid="1222" points="57" swimtime="00:09:31.58" resultid="4494" heatid="7785" lane="8" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:02.07" />
                    <SPLIT distance="100" swimtime="00:04:30.80" />
                    <SPLIT distance="150" swimtime="00:07:03.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="45" swimtime="00:04:31.31" resultid="4495" heatid="7882" lane="1" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:01.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="59" swimtime="00:01:54.92" resultid="4496" heatid="8030" lane="1" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Zbigniew" gender="M" lastname="Krasnodębski" nation="POL" athleteid="4497">
              <RESULTS>
                <RESULT eventid="1222" points="519" reactiontime="+80" swimtime="00:03:22.34" resultid="4498" heatid="7790" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.23" />
                    <SPLIT distance="100" swimtime="00:01:38.12" />
                    <SPLIT distance="150" swimtime="00:02:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="427" reactiontime="+87" swimtime="00:01:30.44" resultid="4499" heatid="7888" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="453" reactiontime="+80" swimtime="00:00:39.69" resultid="4500" heatid="8038" lane="7" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Janusz" gender="M" lastname="Szpala" nation="POL" athleteid="4501">
              <RESULTS>
                <RESULT eventid="1076" points="394" reactiontime="+103" swimtime="00:00:38.42" resultid="4502" heatid="7687" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1108" points="303" reactiontime="+101" swimtime="00:04:00.46" resultid="4503" heatid="7721" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.36" />
                    <SPLIT distance="100" swimtime="00:01:56.01" />
                    <SPLIT distance="150" swimtime="00:03:07.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="342" reactiontime="+104" swimtime="00:01:45.59" resultid="4504" heatid="7839" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="271" reactiontime="+103" swimtime="00:00:47.22" resultid="4505" heatid="7907" lane="1" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Józef" gender="M" lastname="Ciupek" nation="POL" athleteid="4506">
              <RESULTS>
                <RESULT eventid="1076" points="343" reactiontime="+107" swimtime="00:00:40.21" resultid="4507" heatid="7686" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1190" points="343" reactiontime="+85" swimtime="00:00:47.56" resultid="4508" heatid="7767" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1415" points="433" reactiontime="+97" swimtime="00:00:40.39" resultid="4509" heatid="7910" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1655" points="586" reactiontime="+99" swimtime="00:00:42.21" resultid="4510" heatid="8035" lane="3" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Robert" gender="M" lastname="Brysz" nation="POL" athleteid="4511">
              <RESULTS>
                <RESULT eventid="1190" points="536" reactiontime="+69" swimtime="00:00:30.82" resultid="4512" heatid="7776" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1286" points="522" reactiontime="+70" swimtime="00:01:08.54" resultid="4513" heatid="7854" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="472" reactiontime="+72" swimtime="00:01:09.24" resultid="4514" heatid="8001" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Masters Opole  D">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+88" swimtime="00:02:04.68" resultid="4517" heatid="7971" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                    <SPLIT distance="100" swimtime="00:00:59.96" />
                    <SPLIT distance="150" swimtime="00:01:33.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4468" number="1" />
                    <RELAYPOSITION athleteid="4460" number="2" />
                    <RELAYPOSITION athleteid="4497" number="3" />
                    <RELAYPOSITION athleteid="4482" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Masters Opole C">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+63" swimtime="00:02:10.81" resultid="4518" heatid="7870" lane="3" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:41.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4468" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4497" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4511" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="4490" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Masters Opole E">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+106" swimtime="00:02:30.85" resultid="4515" heatid="7970" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:14.80" />
                    <SPLIT distance="150" swimtime="00:01:52.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4501" number="1" />
                    <RELAYPOSITION athleteid="4475" number="2" />
                    <RELAYPOSITION athleteid="4446" number="3" />
                    <RELAYPOSITION athleteid="4451" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1357" reactiontime="+84" swimtime="00:02:36.27" resultid="4516" heatid="7869" lane="8" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="100" swimtime="00:01:24.74" />
                    <SPLIT distance="150" swimtime="00:02:01.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4460" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="4506" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4482" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4451" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02611" nation="POL" clubid="4249" name="TP Weteran  Zabrze" shortname="Weteran  Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW.JANA  4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="502611100002" athleteid="4268">
              <RESULTS>
                <RESULT eventid="1092" points="516" reactiontime="+108" swimtime="00:03:59.55" resultid="4269" heatid="7714" lane="7" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.56" />
                    <SPLIT distance="100" swimtime="00:02:03.76" />
                    <SPLIT distance="150" swimtime="00:03:06.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="586" swimtime="00:15:36.29" resultid="4270" heatid="8715" lane="7" entrytime="00:16:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                    <SPLIT distance="100" swimtime="00:01:47.38" />
                    <SPLIT distance="200" swimtime="00:03:47.59" />
                    <SPLIT distance="300" swimtime="00:05:45.20" />
                    <SPLIT distance="400" swimtime="00:07:43.60" />
                    <SPLIT distance="500" swimtime="00:09:40.84" />
                    <SPLIT distance="600" swimtime="00:11:42.17" />
                    <SPLIT distance="700" swimtime="00:13:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="732" reactiontime="+113" swimtime="00:03:56.56" resultid="4271" heatid="7780" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.91" />
                    <SPLIT distance="100" swimtime="00:01:56.38" />
                    <SPLIT distance="150" swimtime="00:02:58.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="643" reactiontime="+112" swimtime="00:01:52.50" resultid="4272" heatid="7876" lane="2" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="641" reactiontime="+104" swimtime="00:01:49.98" resultid="4273" heatid="7988" lane="6" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="626" reactiontime="+105" swimtime="00:00:50.47" resultid="4274" heatid="8023" lane="2" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="502611200002" athleteid="4275">
              <RESULTS>
                <RESULT eventid="1222" points="701" reactiontime="+92" swimtime="00:03:28.51" resultid="4276" heatid="7789" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.75" />
                    <SPLIT distance="100" swimtime="00:01:40.44" />
                    <SPLIT distance="150" swimtime="00:02:35.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="683" reactiontime="+96" swimtime="00:01:35.01" resultid="4277" heatid="7885" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="460" reactiontime="+96" swimtime="00:00:42.39" resultid="4278" heatid="7909" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1655" points="615" reactiontime="+94" swimtime="00:00:44.01" resultid="4279" heatid="8035" lane="6" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" license="502611200004" athleteid="4280">
              <RESULTS>
                <RESULT eventid="1190" points="475" reactiontime="+72" swimtime="00:00:42.70" resultid="4281" heatid="7768" lane="2" entrytime="00:00:42.27" />
                <RESULT eventid="1447" points="401" reactiontime="+74" swimtime="00:01:38.06" resultid="4282" heatid="7935" lane="2" entrytime="00:01:35.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="363" reactiontime="+73" swimtime="00:03:40.93" resultid="4283" heatid="8012" lane="2" entrytime="00:03:38.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.78" />
                    <SPLIT distance="100" swimtime="00:01:44.97" />
                    <SPLIT distance="150" swimtime="00:02:42.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-05" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" license="502611100005" athleteid="4284">
              <RESULTS>
                <RESULT eventid="1059" points="561" reactiontime="+99" swimtime="00:00:38.97" resultid="4285" heatid="7675" lane="8" entrytime="00:00:40.30" />
                <RESULT eventid="1238" points="512" reactiontime="+94" swimtime="00:01:29.26" resultid="4286" heatid="7798" lane="5" entrytime="00:01:33.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="438" reactiontime="+97" swimtime="00:03:29.14" resultid="4287" heatid="7945" lane="3" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:39.01" />
                    <SPLIT distance="150" swimtime="00:02:34.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="502611100001" athleteid="4288">
              <RESULTS>
                <RESULT eventid="1059" points="831" reactiontime="+79" swimtime="00:00:35.45" resultid="4289" heatid="7677" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1173" points="894" reactiontime="+65" swimtime="00:00:43.41" resultid="4290" heatid="7757" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="1270" points="774" reactiontime="+79" swimtime="00:01:35.15" resultid="4291" heatid="7828" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="639" reactiontime="+81" swimtime="00:00:45.29" resultid="4292" heatid="7899" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1607" points="736" reactiontime="+72" swimtime="00:03:39.12" resultid="4293" heatid="8005" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.70" />
                    <SPLIT distance="100" swimtime="00:01:47.50" />
                    <SPLIT distance="150" swimtime="00:02:45.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-07-16" firstname="Ewald" gender="M" lastname="Bastek" nation="POL" license="502611200001" athleteid="4294">
              <RESULTS>
                <RESULT eventid="1108" points="628" reactiontime="+100" swimtime="00:03:27.53" resultid="4295" heatid="7722" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.77" />
                    <SPLIT distance="100" swimtime="00:01:46.34" />
                    <SPLIT distance="150" swimtime="00:02:44.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="620" reactiontime="+96" swimtime="00:01:31.98" resultid="4296" heatid="7841" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="527" reactiontime="+99" swimtime="00:00:40.50" resultid="4297" heatid="7909" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1703" points="655" reactiontime="+96" swimtime="00:06:25.40" resultid="4298" heatid="9068" lane="7" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                    <SPLIT distance="100" swimtime="00:01:30.51" />
                    <SPLIT distance="150" swimtime="00:02:21.06" />
                    <SPLIT distance="200" swimtime="00:03:10.95" />
                    <SPLIT distance="250" swimtime="00:04:00.42" />
                    <SPLIT distance="300" swimtime="00:04:50.70" />
                    <SPLIT distance="350" swimtime="00:05:40.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-28" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="502611200007" athleteid="4299">
              <RESULTS>
                <RESULT eventid="1076" points="667" reactiontime="+80" swimtime="00:00:30.90" resultid="4300" heatid="7694" lane="6" entrytime="00:00:31.50" />
                <RESULT eventid="1254" points="525" reactiontime="+92" swimtime="00:01:14.20" resultid="4301" heatid="7812" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="636" reactiontime="+83" swimtime="00:00:34.81" resultid="4302" heatid="7913" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="502611100009" athleteid="4303">
              <RESULTS>
                <RESULT eventid="1092" points="721" reactiontime="+81" swimtime="00:02:43.64" resultid="4304" heatid="7718" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:20.19" />
                    <SPLIT distance="150" swimtime="00:02:06.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="736" reactiontime="+86" swimtime="00:03:03.95" resultid="4305" heatid="7783" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                    <SPLIT distance="100" swimtime="00:01:29.01" />
                    <SPLIT distance="150" swimtime="00:02:16.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="631" reactiontime="+91" swimtime="00:01:09.28" resultid="4306" heatid="7803" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="686" reactiontime="+82" swimtime="00:01:25.80" resultid="4307" heatid="7880" lane="7" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="685" reactiontime="+84" swimtime="00:02:27.66" resultid="4308" heatid="7951" lane="8" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:11.84" />
                    <SPLIT distance="150" swimtime="00:01:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="598" reactiontime="+81" swimtime="00:01:18.43" resultid="4309" heatid="7990" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="707" reactiontime="+83" swimtime="00:05:10.84" resultid="4310" heatid="9047" lane="6" entrytime="00:05:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:13.80" />
                    <SPLIT distance="150" swimtime="00:01:53.27" />
                    <SPLIT distance="200" swimtime="00:02:33.01" />
                    <SPLIT distance="250" swimtime="00:03:12.79" />
                    <SPLIT distance="300" swimtime="00:03:52.75" />
                    <SPLIT distance="350" swimtime="00:04:32.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-02" firstname="Władysław" gender="M" lastname="Buczkowski" nation="POL" license="502611200003" athleteid="4311">
              <RESULTS>
                <RESULT eventid="1076" points="611" reactiontime="+83" swimtime="00:00:34.17" resultid="4312" heatid="7688" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1190" points="462" reactiontime="+79" swimtime="00:00:44.83" resultid="4313" heatid="7766" lane="3" entrytime="00:00:46.00" />
                <RESULT eventid="1254" points="678" reactiontime="+101" swimtime="00:01:17.21" resultid="4314" heatid="7810" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="687" reactiontime="+85" swimtime="00:01:34.84" resultid="4315" heatid="7885" lane="3" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="541" reactiontime="+105" swimtime="00:03:04.84" resultid="4316" heatid="7954" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:01:30.45" />
                    <SPLIT distance="150" swimtime="00:02:19.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="779" reactiontime="+77" swimtime="00:00:40.69" resultid="4317" heatid="8033" lane="5" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-14" firstname="Maciej" gender="M" lastname="Kunicki" nation="POL" license="502611200011" athleteid="4318">
              <RESULTS>
                <RESULT eventid="1108" points="429" reactiontime="+88" swimtime="00:02:49.50" resultid="4319" heatid="7729" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:18.46" />
                    <SPLIT distance="150" swimtime="00:02:11.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="407" reactiontime="+84" swimtime="00:02:50.08" resultid="4320" heatid="7863" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:21.72" />
                    <SPLIT distance="150" swimtime="00:02:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="521" reactiontime="+89" swimtime="00:00:31.22" resultid="4321" heatid="7916" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1591" points="488" reactiontime="+87" swimtime="00:01:11.89" resultid="4322" heatid="7999" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-02-24" firstname="Maria" gender="F" lastname="Buczkowska" nation="POL" license="502611100003" athleteid="4323">
              <RESULTS>
                <RESULT eventid="1206" points="573" reactiontime="+114" swimtime="00:04:01.66" resultid="4324" heatid="7779" lane="5" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.34" />
                    <SPLIT distance="100" swimtime="00:02:01.18" />
                    <SPLIT distance="150" swimtime="00:03:04.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="379" reactiontime="+126" swimtime="00:01:53.08" resultid="4325" heatid="7827" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="565" reactiontime="+114" swimtime="00:01:50.23" resultid="4326" heatid="7876" lane="1" entrytime="00:01:51.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="627" reactiontime="+107" swimtime="00:00:48.17" resultid="4327" heatid="8022" lane="1" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-08-16" firstname="Tadeusz" gender="M" lastname="Stuchlik" nation="POL" license="502611200010" athleteid="4328">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="4329" heatid="7732" lane="5" entrytime="00:02:24.00" />
                <RESULT eventid="1190" points="767" reactiontime="+72" swimtime="00:00:29.66" resultid="4330" heatid="7776" lane="3" entrytime="00:00:30.00" />
                <RESULT comment="G8 - Ukończenie wyścigu nie w położeniu na plecach  (Czas: 13:26)" eventid="1286" reactiontime="+79" status="DSQ" swimtime="00:01:05.43" resultid="4331" heatid="7855" lane="8" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="675" reactiontime="+78" swimtime="00:00:28.64" resultid="4332" heatid="7922" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1447" points="779" reactiontime="+82" swimtime="00:01:04.17" resultid="4333" heatid="7942" lane="2" entrytime="00:01:04.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="789" reactiontime="+76" swimtime="00:02:22.25" resultid="4334" heatid="8019" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:09.82" />
                    <SPLIT distance="150" swimtime="00:01:47.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="502611200011" athleteid="4335">
              <RESULTS>
                <RESULT eventid="1190" points="422" reactiontime="+71" swimtime="00:00:39.16" resultid="4336" heatid="7770" lane="1" entrytime="00:00:39.30" />
                <RESULT eventid="1447" points="402" reactiontime="+78" swimtime="00:01:27.81" resultid="4337" heatid="7936" lane="5" entrytime="00:01:28.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="426" reactiontime="+64" swimtime="00:03:12.59" resultid="4338" heatid="8014" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:28.49" />
                    <SPLIT distance="150" swimtime="00:02:17.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-02-18" firstname="Grażyna" gender="F" lastname="Kiszczak" nation="POL" license="502611100006" athleteid="4339">
              <RESULTS>
                <RESULT eventid="1059" points="735" reactiontime="+71" swimtime="00:00:35.62" resultid="4340" heatid="7677" lane="4" entrytime="00:00:35.20" />
                <RESULT eventid="1173" points="977" reactiontime="+71" swimtime="00:00:39.99" resultid="4341" heatid="7758" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1270" points="644" reactiontime="+72" swimtime="00:01:31.55" resultid="4342" heatid="7832" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="688" reactiontime="+74" swimtime="00:00:40.77" resultid="4343" heatid="7900" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1431" points="833" reactiontime="+64" swimtime="00:01:29.13" resultid="4344" heatid="7929" lane="1" entrytime="00:01:28.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="567" reactiontime="+82" swimtime="00:00:46.62" resultid="4345" heatid="8025" lane="4" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-05" firstname="Stanisław" gender="M" lastname="Kiszczak" nation="POL" license="502611200006" athleteid="4346">
              <RESULTS>
                <RESULT eventid="1076" points="562" reactiontime="+92" swimtime="00:00:34.13" resultid="4347" heatid="7692" lane="3" entrytime="00:00:32.50" />
                <RESULT eventid="1190" points="434" reactiontime="+79" swimtime="00:00:44.00" resultid="4348" heatid="7767" lane="5" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-08" firstname="Aurelia" gender="F" lastname="Wrona" nation="POL" license="502611100007" athleteid="4349">
              <RESULTS>
                <RESULT eventid="1059" points="451" reactiontime="+80" swimtime="00:00:39.42" resultid="4350" heatid="7676" lane="8" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-09" firstname="Anna" gender="F" lastname="Karlsson" nation="POL" athleteid="4351">
              <RESULTS>
                <RESULT eventid="1059" points="516" reactiontime="+91" swimtime="00:00:32.57" resultid="4352" heatid="7680" lane="8" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-23" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" license="502611100004" athleteid="4353">
              <RESULTS>
                <RESULT eventid="1059" points="374" reactiontime="+91" swimtime="00:00:44.75" resultid="4354" heatid="7673" lane="8" entrytime="00:00:46.00" />
                <RESULT eventid="1173" points="413" reactiontime="+111" swimtime="00:00:53.75" resultid="4355" heatid="7755" lane="1" entrytime="00:00:53.00" />
                <RESULT eventid="1270" points="321" reactiontime="+87" swimtime="00:01:59.52" resultid="4356" heatid="7827" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="285" reactiontime="+88" swimtime="00:00:56.11" resultid="4357" heatid="7898" lane="1" entrytime="00:00:57.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="502611200005" athleteid="4358">
              <RESULTS>
                <RESULT eventid="1076" points="418" reactiontime="+108" swimtime="00:00:37.66" resultid="4359" heatid="7687" lane="4" entrytime="00:00:36.50" />
                <RESULT eventid="1286" points="305" reactiontime="+110" swimtime="00:01:49.71" resultid="4360" heatid="7840" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="329" reactiontime="+103" swimtime="00:00:44.26" resultid="4361" heatid="7909" lane="7" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-04" firstname="Ulasz" gender="M" lastname="Szanli" nation="POL" athleteid="4362">
              <RESULTS>
                <RESULT eventid="1076" points="255" reactiontime="+106" swimtime="00:00:34.86" resultid="4363" heatid="7689" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1254" points="172" reactiontime="+115" swimtime="00:01:28.18" resultid="4364" heatid="7807" lane="5" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-03" firstname="Marta" gender="F" lastname="Frank" nation="POL" license="502611100008" athleteid="4365">
              <RESULTS>
                <RESULT eventid="1059" points="701" reactiontime="+80" swimtime="00:00:31.26" resultid="4366" heatid="7680" lane="5" entrytime="00:00:32.20" />
                <RESULT eventid="1173" points="840" reactiontime="+68" swimtime="00:00:34.54" resultid="4367" heatid="7760" lane="2" entrytime="00:00:35.90" />
                <RESULT eventid="1270" points="729" reactiontime="+78" swimtime="00:01:18.39" resultid="4368" heatid="7835" lane="6" entrytime="00:01:19.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="661" reactiontime="+84" swimtime="00:00:34.46" resultid="4369" heatid="7900" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1431" points="809" reactiontime="+73" swimtime="00:01:16.12" resultid="4370" heatid="7930" lane="3" entrytime="00:01:17.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="699" reactiontime="+79" swimtime="00:02:53.24" resultid="4371" heatid="8008" lane="6" entrytime="00:02:53.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="150" swimtime="00:02:09.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-21" firstname="Marek" gender="M" lastname="Rother" nation="POL" license="502611200009" athleteid="4372">
              <RESULTS>
                <RESULT eventid="1190" points="917" reactiontime="+64" swimtime="00:00:29.49" resultid="4373" heatid="7776" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1286" points="766" reactiontime="+72" swimtime="00:01:06.10" resultid="4374" heatid="7852" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="761" reactiontime="+78" swimtime="00:00:28.95" resultid="4375" heatid="7911" lane="4" entrytime="00:00:36.50" />
                <RESULT eventid="1447" points="916" reactiontime="+71" swimtime="00:01:03.99" resultid="4376" heatid="7942" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="926" reactiontime="+67" swimtime="00:02:19.83" resultid="4377" heatid="8019" lane="3" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:07.82" />
                    <SPLIT distance="150" swimtime="00:01:43.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="M" name="Weteran Zabrze  F" number="4">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+70" swimtime="00:02:43.25" resultid="4381" heatid="7868" lane="3" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                    <SPLIT distance="100" swimtime="00:01:29.00" />
                    <SPLIT distance="150" swimtime="00:02:08.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4280" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4275" number="2" reactiontime="+12" />
                    <RELAYPOSITION athleteid="4294" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4311" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Weteran Zabrze D" number="5">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+67" swimtime="00:02:09.20" resultid="4382" heatid="7869" lane="1" entrytime="00:02:31.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="100" swimtime="00:01:02.74" />
                    <SPLIT distance="150" swimtime="00:01:38.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4372" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="4328" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4299" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="4335" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="M" name="Weteran Zabrze F" number="7">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+105" swimtime="00:02:19.30" resultid="4384" heatid="7970" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:10.52" />
                    <SPLIT distance="150" swimtime="00:01:47.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4311" number="1" />
                    <RELAYPOSITION athleteid="4275" number="2" />
                    <RELAYPOSITION athleteid="4294" number="3" />
                    <RELAYPOSITION athleteid="4346" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Weteran Zabrze E" number="8">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+87" swimtime="00:02:15.19" resultid="4385" heatid="7970" lane="4" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:10.25" />
                    <SPLIT distance="150" swimtime="00:01:47.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4299" number="1" />
                    <RELAYPOSITION athleteid="4358" number="2" />
                    <RELAYPOSITION athleteid="4280" number="3" />
                    <RELAYPOSITION athleteid="4372" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" name="Weteran Zabrze E" number="3">
              <RESULTS>
                <RESULT eventid="1334" reactiontime="+67" swimtime="00:02:38.33" resultid="4380" heatid="7866" lane="3" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                    <SPLIT distance="100" swimtime="00:01:28.70" />
                    <SPLIT distance="150" swimtime="00:02:03.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4339" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="4323" number="2" reactiontime="+105" />
                    <RELAYPOSITION athleteid="4365" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="4288" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" name="Weteran Zabrze E" number="6">
              <RESULTS>
                <RESULT eventid="1495" reactiontime="+82" swimtime="00:02:31.50" resultid="4383" heatid="7968" lane="6" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:00.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4288" number="1" />
                    <RELAYPOSITION athleteid="4353" number="2" />
                    <RELAYPOSITION athleteid="4284" number="3" />
                    <RELAYPOSITION athleteid="4365" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="X" name="Weteran Zabrze F" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+79" swimtime="00:02:24.32" resultid="4378" heatid="7735" lane="1" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:47.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4288" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4294" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4275" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4339" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Weteran Zabrze E" number="2">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+99" swimtime="00:02:19.64" resultid="4379" heatid="7735" lane="7" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:01:48.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4284" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="4349" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="4299" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="4346" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="X" name="Weteran Zabrze F" number="9">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+74" swimtime="00:02:45.22" resultid="4386" heatid="8050" lane="2" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:01:25.46" />
                    <SPLIT distance="150" swimtime="00:02:09.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4339" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4275" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="4294" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="4288" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Weteran Zabrze E" number="10">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+67" swimtime="00:02:48.11" resultid="4387" heatid="8050" lane="1" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:01:33.50" />
                    <SPLIT distance="150" swimtime="00:02:08.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4280" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="4268" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4299" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="4284" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Weteran Zabrze D" number="11">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+71" swimtime="00:02:16.94" resultid="4388" heatid="8052" lane="8" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:01:17.58" />
                    <SPLIT distance="150" swimtime="00:01:45.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4372" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4323" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4328" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="4365" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00215" nation="POL" region="15" clubid="5497" name="TS Olimpia Poznań" shortname="Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="5498">
              <RESULTS>
                <RESULT eventid="1059" points="567" reactiontime="+94" swimtime="00:00:38.83" resultid="5499" heatid="7676" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1238" points="517" reactiontime="+94" swimtime="00:01:28.93" resultid="5500" heatid="7798" lane="3" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="475" reactiontime="+102" swimtime="00:01:41.32" resultid="5501" heatid="7828" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="382" reactiontime="+101" swimtime="00:00:49.60" resultid="5502" heatid="7898" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1463" points="512" reactiontime="+96" swimtime="00:03:18.63" resultid="5503" heatid="7945" lane="5" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.44" />
                    <SPLIT distance="100" swimtime="00:01:37.51" />
                    <SPLIT distance="150" swimtime="00:02:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="485" reactiontime="+94" swimtime="00:00:49.12" resultid="5504" heatid="8022" lane="5" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Janusz" gender="M" lastname="Woch" nation="POL" athleteid="5505">
              <RESULTS>
                <RESULT eventid="1108" points="409" reactiontime="+77" swimtime="00:03:37.62" resultid="5506" heatid="7722" lane="8" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                    <SPLIT distance="100" swimtime="00:01:42.93" />
                    <SPLIT distance="150" swimtime="00:02:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="482" reactiontime="+89" swimtime="00:03:52.21" resultid="5507" heatid="7788" lane="5" entrytime="00:03:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                    <SPLIT distance="100" swimtime="00:01:51.24" />
                    <SPLIT distance="150" swimtime="00:02:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="479" reactiontime="+81" swimtime="00:01:34.43" resultid="5508" heatid="7841" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="448" reactiontime="+79" swimtime="00:01:43.73" resultid="5509" heatid="7884" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="383" reactiontime="+106" swimtime="00:01:39.64" resultid="5510" heatid="7935" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="407" reactiontime="+82" swimtime="00:03:32.59" resultid="5511" heatid="8012" lane="5" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.43" />
                    <SPLIT distance="100" swimtime="00:01:42.60" />
                    <SPLIT distance="150" swimtime="00:02:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="525" reactiontime="+85" swimtime="00:00:43.79" resultid="5512" heatid="8034" lane="3" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="5513">
              <RESULTS>
                <RESULT eventid="1156" points="427" swimtime="00:28:22.50" resultid="5514" heatid="8724" lane="5" entrytime="00:28:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:43.48" />
                    <SPLIT distance="200" swimtime="00:03:34.77" />
                    <SPLIT distance="300" swimtime="00:05:25.76" />
                    <SPLIT distance="400" swimtime="00:07:19.31" />
                    <SPLIT distance="500" swimtime="00:09:14.92" />
                    <SPLIT distance="600" swimtime="00:11:11.60" />
                    <SPLIT distance="700" swimtime="00:13:05.75" />
                    <SPLIT distance="800" swimtime="00:15:01.05" />
                    <SPLIT distance="900" swimtime="00:16:56.04" />
                    <SPLIT distance="1000" swimtime="00:18:52.88" />
                    <SPLIT distance="1100" swimtime="00:20:48.07" />
                    <SPLIT distance="1200" swimtime="00:22:43.15" />
                    <SPLIT distance="1300" swimtime="00:24:37.95" />
                    <SPLIT distance="1400" swimtime="00:26:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="450" reactiontime="+79" swimtime="00:00:43.23" resultid="5515" heatid="7768" lane="1" entrytime="00:00:42.50" />
                <RESULT eventid="1447" points="418" reactiontime="+78" swimtime="00:01:37.23" resultid="5516" heatid="7935" lane="4" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="5517" heatid="8012" lane="6" entrytime="00:03:35.00" />
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="5518" heatid="9069" lane="6" entrytime="00:06:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="5519">
              <RESULTS>
                <RESULT eventid="1108" points="512" reactiontime="+93" swimtime="00:03:05.23" resultid="5520" heatid="7725" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:31.00" />
                    <SPLIT distance="150" swimtime="00:02:22.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="448" reactiontime="+81" swimtime="00:00:41.11" resultid="5521" heatid="7769" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1286" points="550" reactiontime="+89" swimtime="00:01:24.41" resultid="5522" heatid="7845" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="482" reactiontime="+82" swimtime="00:01:27.54" resultid="5523" heatid="7937" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="553" reactiontime="+102" swimtime="00:06:34.77" resultid="5524" heatid="8809" lane="7" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.18" />
                    <SPLIT distance="100" swimtime="00:01:41.51" />
                    <SPLIT distance="150" swimtime="00:02:30.82" />
                    <SPLIT distance="200" swimtime="00:03:18.83" />
                    <SPLIT distance="250" swimtime="00:04:12.38" />
                    <SPLIT distance="300" swimtime="00:05:06.00" />
                    <SPLIT distance="350" swimtime="00:05:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="586" reactiontime="+89" swimtime="00:03:05.17" resultid="5525" heatid="8014" lane="5" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:01:30.10" />
                    <SPLIT distance="150" swimtime="00:02:17.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="413" reactiontime="+89" swimtime="00:00:40.94" resultid="5526" heatid="8038" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="5527">
              <RESULTS>
                <RESULT eventid="1108" points="565" reactiontime="+76" swimtime="00:02:45.18" resultid="5528" heatid="7728" lane="7" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                    <SPLIT distance="150" swimtime="00:02:06.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="600" reactiontime="+83" swimtime="00:02:56.89" resultid="5529" heatid="7793" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:10.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="622" reactiontime="+84" swimtime="00:01:18.71" resultid="5530" heatid="7892" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="511" reactiontime="+84" swimtime="00:02:23.48" resultid="5531" heatid="7963" lane="7" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:08.74" />
                    <SPLIT distance="150" swimtime="00:01:46.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="462" reactiontime="+81" swimtime="00:01:16.02" resultid="5532" heatid="7998" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="646" reactiontime="+80" swimtime="00:00:35.48" resultid="5533" heatid="8043" lane="4" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Ryszard" gender="M" lastname="Krzyżanowski" nation="POL" athleteid="5534">
              <RESULTS>
                <RESULT eventid="1076" points="556" reactiontime="+104" swimtime="00:00:32.82" resultid="5535" heatid="7693" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1254" points="437" reactiontime="+99" swimtime="00:01:18.85" resultid="5536" heatid="7812" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="350" reactiontime="+121" swimtime="00:00:42.48" resultid="5537" heatid="7912" lane="6" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Bartłomiej" gender="M" lastname="Zadorożny" nation="POL" athleteid="5538">
              <RESULTS>
                <RESULT eventid="1076" points="628" reactiontime="+85" swimtime="00:00:27.69" resultid="5539" heatid="7703" lane="2" entrytime="00:00:28.04" />
                <RESULT eventid="1254" points="580" reactiontime="+83" swimtime="00:01:01.66" resultid="5540" heatid="7818" lane="4" entrytime="00:01:03.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="540" reactiontime="+84" swimtime="00:01:18.60" resultid="5541" heatid="7892" lane="8" entrytime="00:01:21.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="428" reactiontime="+86" swimtime="00:02:27.90" resultid="5542" heatid="7965" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="100" swimtime="00:01:07.08" />
                    <SPLIT distance="150" swimtime="00:01:46.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="563" reactiontime="+80" swimtime="00:00:34.95" resultid="5543" heatid="8043" lane="6" entrytime="00:00:35.73" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Olimpia Poznań D">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+80" swimtime="00:02:04.58" resultid="5545" heatid="7972" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:01:02.21" />
                    <SPLIT distance="150" swimtime="00:01:36.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5527" number="1" />
                    <RELAYPOSITION athleteid="5519" number="2" />
                    <RELAYPOSITION athleteid="5534" number="3" />
                    <RELAYPOSITION athleteid="5538" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Olimpia Poznań E">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+74" swimtime="00:02:31.66" resultid="5544" heatid="7869" lane="7" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:01:24.81" />
                    <SPLIT distance="150" swimtime="00:01:57.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5513" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="5505" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="5527" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="5534" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01806" nation="POL" region="06" clubid="2611" name="TS Wisła Masters Kraków" shortname="Wisła Masters Kraków">
          <ATHLETES>
            <ATHLETE birthdate="1930-01-01" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="2612">
              <RESULTS>
                <RESULT eventid="1076" points="559" reactiontime="+114" swimtime="00:00:40.33" resultid="2613" heatid="7687" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1108" points="626" reactiontime="+124" swimtime="00:04:01.29" resultid="2614" heatid="7721" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.49" />
                    <SPLIT distance="100" swimtime="00:02:02.03" />
                    <SPLIT distance="150" swimtime="00:03:09.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="601" reactiontime="+80" swimtime="00:00:51.77" resultid="2615" heatid="7763" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1286" points="620" reactiontime="+118" swimtime="00:01:48.18" resultid="2616" heatid="7840" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="432" reactiontime="+115" swimtime="00:00:58.73" resultid="2617" heatid="7906" lane="4" entrytime="00:00:57.00" />
                <RESULT eventid="1543" points="551" reactiontime="+124" swimtime="00:09:04.08" resultid="2618" heatid="8811" lane="8" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.98" />
                    <SPLIT distance="100" swimtime="00:02:25.60" />
                    <SPLIT distance="150" swimtime="00:03:35.33" />
                    <SPLIT distance="200" swimtime="00:04:47.22" />
                    <SPLIT distance="250" swimtime="00:06:00.19" />
                    <SPLIT distance="300" swimtime="00:07:13.64" />
                    <SPLIT distance="350" swimtime="00:08:08.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="583" reactiontime="+109" swimtime="00:00:53.83" resultid="2619" heatid="8030" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1703" points="665" reactiontime="+113" swimtime="00:07:26.87" resultid="2620" heatid="9069" lane="7" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:38.09" />
                    <SPLIT distance="150" swimtime="00:02:33.87" />
                    <SPLIT distance="200" swimtime="00:03:30.66" />
                    <SPLIT distance="250" swimtime="00:04:28.67" />
                    <SPLIT distance="300" swimtime="00:05:26.99" />
                    <SPLIT distance="350" swimtime="00:06:27.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Janusz" gender="M" lastname="Konstanty" nation="POL" athleteid="2621">
              <RESULTS>
                <RESULT eventid="1108" points="573" reactiontime="+89" swimtime="00:02:58.35" resultid="2622" heatid="7726" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:01:20.56" />
                    <SPLIT distance="150" swimtime="00:02:15.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="658" reactiontime="+79" swimtime="00:00:36.18" resultid="2623" heatid="7770" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1286" points="643" reactiontime="+93" swimtime="00:01:20.15" resultid="2624" heatid="7844" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="646" reactiontime="+80" swimtime="00:01:19.39" resultid="2625" heatid="7938" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="682" reactiontime="+89" swimtime="00:02:56.11" resultid="2626" heatid="8014" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:24.82" />
                    <SPLIT distance="150" swimtime="00:02:11.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Paulina" gender="F" lastname="Palka" nation="POL" athleteid="2627">
              <RESULTS>
                <RESULT eventid="1173" points="721" reactiontime="+65" swimtime="00:00:33.79" resultid="2628" heatid="7761" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1270" points="593" reactiontime="+68" swimtime="00:01:17.48" resultid="2629" heatid="7835" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="721" reactiontime="+58" swimtime="00:01:12.69" resultid="2630" heatid="7931" lane="3" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="754" reactiontime="+58" swimtime="00:02:38.02" resultid="2631" heatid="8009" lane="2" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:16.48" />
                    <SPLIT distance="150" swimtime="00:01:57.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Wojciech" gender="M" lastname="Wolski" nation="POL" athleteid="2632">
              <RESULTS>
                <RESULT eventid="1655" points="482" reactiontime="+90" swimtime="00:00:39.13" resultid="2633" heatid="8029" lane="4" />
                <RESULT eventid="1286" points="360" reactiontime="+90" swimtime="00:01:25.01" resultid="6205" heatid="7838" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Piotr Krzysztof" gender="M" lastname="Dąbski" nation="POL" athleteid="2634">
              <RESULTS>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="2635" heatid="7859" lane="1" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="2636" heatid="7906" lane="2" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="2637" heatid="7992" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Stanisław" gender="M" lastname="Trzaska" nation="POL" athleteid="2638">
              <RESULTS>
                <RESULT eventid="1156" points="609" swimtime="00:22:46.42" resultid="2639" heatid="8721" lane="3" entrytime="00:23:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.87" />
                    <SPLIT distance="100" swimtime="00:01:24.07" />
                    <SPLIT distance="200" swimtime="00:02:52.90" />
                    <SPLIT distance="300" swimtime="00:04:22.95" />
                    <SPLIT distance="400" swimtime="00:05:53.67" />
                    <SPLIT distance="500" swimtime="00:07:24.89" />
                    <SPLIT distance="600" swimtime="00:08:56.17" />
                    <SPLIT distance="700" swimtime="00:10:26.53" />
                    <SPLIT distance="800" swimtime="00:11:57.69" />
                    <SPLIT distance="900" swimtime="00:13:29.46" />
                    <SPLIT distance="1000" swimtime="00:15:01.61" />
                    <SPLIT distance="1100" swimtime="00:16:34.65" />
                    <SPLIT distance="1200" swimtime="00:18:07.35" />
                    <SPLIT distance="1300" swimtime="00:19:41.02" />
                    <SPLIT distance="1400" swimtime="00:21:14.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" status="WDR" swimtime="00:00:00.00" resultid="2640" heatid="7809" lane="4" entrytime="00:01:20.00" />
                <RESULT eventid="1623" points="436" reactiontime="+131" swimtime="00:03:24.40" resultid="2641" heatid="8014" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.89" />
                    <SPLIT distance="100" swimtime="00:02:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="548" reactiontime="+122" swimtime="00:05:53.04" resultid="2642" heatid="9067" lane="6" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="100" swimtime="00:01:23.84" />
                    <SPLIT distance="150" swimtime="00:02:08.76" />
                    <SPLIT distance="200" swimtime="00:02:53.53" />
                    <SPLIT distance="250" swimtime="00:03:38.52" />
                    <SPLIT distance="300" swimtime="00:04:24.05" />
                    <SPLIT distance="350" swimtime="00:05:09.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Michał" gender="M" lastname="Syryca" nation="POL" athleteid="2643">
              <RESULTS>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="2644" heatid="7906" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Mateusz" gender="M" lastname="Dybek" nation="POL" athleteid="3581">
              <RESULTS>
                <RESULT eventid="1076" points="589" reactiontime="+76" swimtime="00:00:26.40" resultid="3582" heatid="7707" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1254" points="588" reactiontime="+77" swimtime="00:00:58.53" resultid="3583" heatid="7822" lane="8" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="486" reactiontime="+83" swimtime="00:02:15.41" resultid="3584" heatid="7962" lane="1" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:05.61" />
                    <SPLIT distance="150" swimtime="00:01:41.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="472" reactiontime="+82" swimtime="00:05:08.43" resultid="3585" heatid="9064" lane="3" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                    <SPLIT distance="150" swimtime="00:01:52.08" />
                    <SPLIT distance="200" swimtime="00:02:32.20" />
                    <SPLIT distance="250" swimtime="00:03:12.22" />
                    <SPLIT distance="300" swimtime="00:03:52.33" />
                    <SPLIT distance="350" swimtime="00:04:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="425" swimtime="00:22:20.84" resultid="3586" heatid="8720" lane="8" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                    <SPLIT distance="100" swimtime="00:01:20.35" />
                    <SPLIT distance="200" swimtime="00:02:49.08" />
                    <SPLIT distance="300" swimtime="00:04:19.22" />
                    <SPLIT distance="400" swimtime="00:05:47.92" />
                    <SPLIT distance="500" swimtime="00:07:20.73" />
                    <SPLIT distance="600" swimtime="00:08:53.30" />
                    <SPLIT distance="700" swimtime="00:10:25.30" />
                    <SPLIT distance="800" swimtime="00:11:56.79" />
                    <SPLIT distance="900" swimtime="00:13:29.26" />
                    <SPLIT distance="1000" swimtime="00:15:01.38" />
                    <SPLIT distance="1100" swimtime="00:16:33.40" />
                    <SPLIT distance="1200" swimtime="00:18:03.60" />
                    <SPLIT distance="1300" swimtime="00:19:34.04" />
                    <SPLIT distance="1400" swimtime="00:21:00.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Agnieszka" gender="F" lastname="Leńczowska" nation="POL" athleteid="3587">
              <RESULTS>
                <RESULT eventid="1059" points="626" reactiontime="+81" swimtime="00:00:30.55" resultid="3589" heatid="7682" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1092" points="586" reactiontime="+86" swimtime="00:02:50.92" resultid="3590" heatid="7718" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:19.08" />
                    <SPLIT distance="150" swimtime="00:02:09.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="609" reactiontime="+62" swimtime="00:00:35.81" resultid="3591" heatid="7759" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1270" points="589" reactiontime="+80" swimtime="00:01:17.65" resultid="3592" heatid="7836" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="600" reactiontime="+65" swimtime="00:02:47.82" resultid="3593" heatid="8008" lane="5" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                    <SPLIT distance="100" swimtime="00:01:20.46" />
                    <SPLIT distance="150" swimtime="00:02:04.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-10" firstname="Dariusz" gender="M" lastname="Wesołowski" nation="POL" athleteid="6206">
              <RESULTS>
                <RESULT eventid="1254" points="451" reactiontime="+88" swimtime="00:01:07.86" resultid="6207" heatid="7816" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="370" reactiontime="+85" swimtime="00:02:37.40" resultid="6208" heatid="7961" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:02:00.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Ewa" gender="F" lastname="Macierzewska" nation="POL" athleteid="6341">
              <RESULTS>
                <RESULT eventid="1059" points="76" reactiontime="+131" swimtime="00:01:18.58" resultid="6342" heatid="7671" lane="3" />
                <RESULT eventid="1173" points="165" reactiontime="+101" swimtime="00:01:16.20" resultid="6343" heatid="7753" lane="3" />
                <RESULT eventid="1206" status="DNS" swimtime="00:00:00.00" resultid="6344" heatid="7778" lane="3" />
                <RESULT eventid="1366" points="159" reactiontime="+140" swimtime="00:02:59.21" resultid="6345" heatid="7873" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.73" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K15 - Brak dotknięcia ściany obydwoma rozłączonymi dłońmi przy nawrocie lub na zakończenie wyścigu" eventid="1639" reactiontime="+118" status="DSQ" swimtime="00:01:18.42" resultid="6346" heatid="8020" lane="3" />
                <RESULT eventid="1431" status="DNS" swimtime="00:00:00.00" resultid="6347" heatid="7926" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Wisła Kraków Masters E">
              <RESULTS>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="8782" heatid="7868" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2612" number="1" />
                    <RELAYPOSITION athleteid="2621" number="2" />
                    <RELAYPOSITION athleteid="2638" number="3" />
                    <RELAYPOSITION athleteid="2632" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Wisa Masters  Kraków E" number="1">
              <RESULTS>
                <RESULT eventid="1357" status="WDR" swimtime="00:00:00.00" resultid="2645">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2612" number="1" />
                    <RELAYPOSITION athleteid="2621" number="2" />
                    <RELAYPOSITION athleteid="2638" number="3" />
                    <RELAYPOSITION athleteid="2632" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WOTAR" nation="POL" region="06" clubid="4713" name="Tarnowskie WOPR Masters">
          <CONTACT city="tarnów" email="przemoju@gmail.com" name="przemek jurek" phone="533633523" state="MAŁ" street="bat. chłopskich 2" zip="33-101" />
          <ATHLETES>
            <ATHLETE birthdate="1983-04-24" firstname="Radosław" gender="M" lastname="Jurek" nation="POL" athleteid="4714">
              <RESULTS>
                <RESULT eventid="1108" points="305" reactiontime="+88" swimtime="00:02:55.41" resultid="4715" heatid="7730" lane="8" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:19.90" />
                    <SPLIT distance="150" swimtime="00:02:14.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="398" reactiontime="+82" swimtime="00:00:36.00" resultid="4716" heatid="7771" lane="5" entrytime="00:00:35.20" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="4717" heatid="7864" lane="4" entrytime="00:02:45.00" />
                <RESULT eventid="1415" points="394" reactiontime="+85" swimtime="00:00:31.19" resultid="4718" heatid="7920" lane="4" entrytime="00:00:29.50" />
                <RESULT eventid="1591" points="349" reactiontime="+89" swimtime="00:01:14.73" resultid="4719" heatid="8000" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="433" reactiontime="+85" swimtime="00:00:36.76" resultid="4720" heatid="8042" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-07-08" firstname="Andrzej" gender="M" lastname="Maciejczak" nation="POL" athleteid="4721">
              <RESULTS>
                <RESULT eventid="1076" points="439" reactiontime="+88" swimtime="00:00:33.41" resultid="4722" heatid="7691" lane="8" entrytime="00:00:33.30" />
                <RESULT eventid="1156" points="316" swimtime="00:26:07.90" resultid="4723" heatid="8722" lane="7" entrytime="00:26:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:24.45" />
                    <SPLIT distance="200" swimtime="00:03:03.72" />
                    <SPLIT distance="300" swimtime="00:04:46.05" />
                    <SPLIT distance="400" swimtime="00:06:29.50" />
                    <SPLIT distance="500" swimtime="00:08:14.43" />
                    <SPLIT distance="600" swimtime="00:09:59.61" />
                    <SPLIT distance="700" swimtime="00:11:45.42" />
                    <SPLIT distance="800" swimtime="00:13:32.37" />
                    <SPLIT distance="900" swimtime="00:15:19.21" />
                    <SPLIT distance="1000" swimtime="00:17:06.36" />
                    <SPLIT distance="1100" swimtime="00:18:54.11" />
                    <SPLIT distance="1200" swimtime="00:20:42.25" />
                    <SPLIT distance="1300" swimtime="00:22:31.27" />
                    <SPLIT distance="1400" swimtime="00:24:21.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="377" reactiontime="+108" swimtime="00:01:18.06" resultid="4724" heatid="7810" lane="1" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="4725" heatid="7839" lane="6" entrytime="00:01:57.00" />
                <RESULT eventid="1415" points="252" reactiontime="+110" swimtime="00:00:43.60" resultid="4726" heatid="7908" lane="6" entrytime="00:00:43.50" />
                <RESULT eventid="1479" points="346" reactiontime="+103" swimtime="00:02:59.09" resultid="4727" heatid="7955" lane="6" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:25.12" />
                    <SPLIT distance="150" swimtime="00:02:12.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="337" reactiontime="+105" swimtime="00:06:22.76" resultid="4728" heatid="9068" lane="4" entrytime="00:06:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:24.59" />
                    <SPLIT distance="150" swimtime="00:02:15.54" />
                    <SPLIT distance="200" swimtime="00:03:05.91" />
                    <SPLIT distance="250" swimtime="00:03:56.01" />
                    <SPLIT distance="300" swimtime="00:04:46.15" />
                    <SPLIT distance="350" swimtime="00:05:35.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-23" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" athleteid="4729">
              <RESULTS>
                <RESULT eventid="1092" points="604" reactiontime="+93" swimtime="00:02:49.33" resultid="4730" heatid="7717" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:02:08.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="692" reactiontime="+75" swimtime="00:00:34.90" resultid="4731" heatid="7761" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1270" points="580" reactiontime="+88" swimtime="00:01:18.43" resultid="4732" heatid="7836" lane="7" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="624" reactiontime="+76" swimtime="00:01:14.61" resultid="4733" heatid="7931" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="607" reactiontime="+77" swimtime="00:02:41.07" resultid="4734" heatid="8009" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:18.83" />
                    <SPLIT distance="150" swimtime="00:02:00.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-07" firstname="Łukasz" gender="M" lastname="Litwora" nation="POL" athleteid="4735">
              <RESULTS>
                <RESULT eventid="1076" points="611" reactiontime="+75" swimtime="00:00:27.94" resultid="4736" heatid="7708" lane="7" entrytime="00:00:26.80" />
                <RESULT eventid="1254" points="477" reactiontime="+78" swimtime="00:01:05.78" resultid="4737" heatid="7821" lane="2" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-14" firstname="Agnieszka" gender="F" lastname="Opitz" nation="POL" athleteid="4738">
              <RESULTS>
                <RESULT eventid="1092" points="574" reactiontime="+82" swimtime="00:02:52.02" resultid="4739" heatid="7717" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:23.11" />
                    <SPLIT distance="150" swimtime="00:02:12.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="542" reactiontime="+93" swimtime="00:03:11.55" resultid="4740" heatid="7783" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.42" />
                    <SPLIT distance="100" swimtime="00:01:32.20" />
                    <SPLIT distance="150" swimtime="00:02:22.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="572" reactiontime="+81" swimtime="00:01:18.41" resultid="4741" heatid="7837" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="633" reactiontime="+76" swimtime="00:00:33.84" resultid="4742" heatid="7904" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1463" points="549" reactiontime="+91" swimtime="00:02:33.74" resultid="4743" heatid="7950" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="150" swimtime="00:01:54.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="544" reactiontime="+81" swimtime="00:01:18.11" resultid="4744" heatid="7991" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="553" reactiontime="+86" swimtime="00:00:38.67" resultid="4745" heatid="8028" lane="1" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-25" firstname="Adam" gender="M" lastname="Wytrwał" nation="POL" athleteid="4746">
              <RESULTS>
                <RESULT eventid="1156" points="303" swimtime="00:24:44.21" resultid="4747" heatid="8722" lane="2" entrytime="00:26:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:26.21" />
                    <SPLIT distance="200" swimtime="00:03:01.50" />
                    <SPLIT distance="300" swimtime="00:04:40.65" />
                    <SPLIT distance="400" swimtime="00:06:20.44" />
                    <SPLIT distance="500" swimtime="00:08:00.61" />
                    <SPLIT distance="600" swimtime="00:09:41.62" />
                    <SPLIT distance="700" swimtime="00:11:21.83" />
                    <SPLIT distance="800" swimtime="00:13:03.39" />
                    <SPLIT distance="900" swimtime="00:14:43.69" />
                    <SPLIT distance="1000" swimtime="00:16:24.67" />
                    <SPLIT distance="1100" swimtime="00:18:06.83" />
                    <SPLIT distance="1200" swimtime="00:19:47.61" />
                    <SPLIT distance="1300" swimtime="00:21:27.91" />
                    <SPLIT distance="1400" swimtime="00:23:10.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="382" reactiontime="+75" swimtime="00:01:11.74" resultid="4748" heatid="7814" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="349" reactiontime="+80" swimtime="00:01:24.94" resultid="4749" heatid="7847" lane="4" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="285" reactiontime="+82" swimtime="00:02:51.57" resultid="4750" heatid="7960" lane="6" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:21.86" />
                    <SPLIT distance="150" swimtime="00:02:07.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="255" reactiontime="+91" swimtime="00:06:19.39" resultid="4751" heatid="9063" lane="1" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:25.15" />
                    <SPLIT distance="150" swimtime="00:02:12.74" />
                    <SPLIT distance="200" swimtime="00:03:02.76" />
                    <SPLIT distance="250" swimtime="00:03:52.46" />
                    <SPLIT distance="300" swimtime="00:04:42.93" />
                    <SPLIT distance="350" swimtime="00:05:32.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-11-13" firstname="Barbara" gender="F" lastname="Wytrwał" nation="POL" athleteid="4752">
              <RESULTS>
                <RESULT eventid="1059" points="104" reactiontime="+120" swimtime="00:00:57.68" resultid="4753" heatid="7672" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="1270" points="58" reactiontime="+121" swimtime="00:02:55.26" resultid="4754" heatid="7826" lane="4" entrytime="00:02:22.00" />
                <RESULT eventid="1463" reactiontime="+139" status="DNF" swimtime="00:00:00.00" resultid="4755" heatid="7944" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.20" />
                    <SPLIT distance="100" swimtime="00:03:43.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" status="DNS" swimtime="00:00:00.00" resultid="4756" heatid="8022" lane="7" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-27" firstname="Miłosz" gender="M" lastname="Pagacz" nation="POL" athleteid="4757">
              <RESULTS>
                <RESULT eventid="1076" points="210" reactiontime="+141" swimtime="00:00:38.67" resultid="4758" heatid="7684" lane="7" />
                <RESULT eventid="1254" points="167" reactiontime="+84" swimtime="00:01:32.34" resultid="4759" heatid="7806" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="139" reactiontime="+191" swimtime="00:03:32.11" resultid="4760" heatid="7952" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                    <SPLIT distance="100" swimtime="00:01:35.02" />
                    <SPLIT distance="150" swimtime="00:02:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="156" reactiontime="+134" swimtime="00:07:35.02" resultid="4761" heatid="9070" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                    <SPLIT distance="100" swimtime="00:01:35.98" />
                    <SPLIT distance="150" swimtime="00:02:33.37" />
                    <SPLIT distance="200" swimtime="00:03:33.00" />
                    <SPLIT distance="250" swimtime="00:04:32.86" />
                    <SPLIT distance="300" swimtime="00:05:36.19" />
                    <SPLIT distance="350" swimtime="00:06:36.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-08-30" firstname="Norbert" gender="M" lastname="Charchouli" nation="POL" athleteid="4762">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="4763" heatid="7722" lane="5" entrytime="00:03:30.00" />
                <RESULT eventid="1190" points="217" reactiontime="+77" swimtime="00:00:45.15" resultid="4764" heatid="7769" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1254" points="274" reactiontime="+82" swimtime="00:01:19.12" resultid="4765" heatid="7809" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="243" reactiontime="+77" swimtime="00:01:34.65" resultid="4766" heatid="7935" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="219" reactiontime="+90" swimtime="00:03:04.91" resultid="4767" heatid="7957" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:22.64" />
                    <SPLIT distance="150" swimtime="00:02:13.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="240" reactiontime="+78" swimtime="00:03:29.01" resultid="4768" heatid="8014" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.87" />
                    <SPLIT distance="100" swimtime="00:01:41.09" />
                    <SPLIT distance="150" swimtime="00:02:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="316" reactiontime="+86" swimtime="00:00:42.38" resultid="4769" heatid="8034" lane="6" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-16" firstname="Maciej" gender="M" lastname="Kacer" nation="POL" athleteid="4770">
              <RESULTS>
                <RESULT eventid="1415" points="682" reactiontime="+68" swimtime="00:00:25.98" resultid="4771" heatid="7925" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1655" points="816" reactiontime="+70" swimtime="00:00:29.75" resultid="4772" heatid="8048" lane="3" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-23" firstname="Mateusz" gender="M" lastname="Dymiter" nation="POL" athleteid="4773">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4774" heatid="7705" lane="2" entrytime="00:00:27.70" />
                <RESULT eventid="1108" points="401" reactiontime="+84" swimtime="00:02:43.40" resultid="4775" heatid="7729" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:02:04.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="448" reactiontime="+100" swimtime="00:01:03.47" resultid="4776" heatid="7817" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="423" reactiontime="+88" swimtime="00:01:13.52" resultid="4777" heatid="7850" lane="7" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="467" reactiontime="+90" swimtime="00:05:51.55" resultid="4778" heatid="8807" lane="1" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:14.16" />
                    <SPLIT distance="150" swimtime="00:02:02.64" />
                    <SPLIT distance="200" swimtime="00:02:49.73" />
                    <SPLIT distance="250" swimtime="00:03:40.77" />
                    <SPLIT distance="300" swimtime="00:04:30.30" />
                    <SPLIT distance="350" swimtime="00:05:12.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="4779" heatid="9063" lane="2" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-06-18" firstname="Paweł" gender="M" lastname="Pasryszko" nation="POL" athleteid="4780">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4781" heatid="7687" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="4782" heatid="7790" lane="5" entrytime="00:03:20.00" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="4783" heatid="7808" lane="8" entrytime="00:01:29.00" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="4784" heatid="7885" lane="2" entrytime="00:01:39.00" />
                <RESULT eventid="1655" points="263" reactiontime="+115" swimtime="00:00:45.05" resultid="4785" heatid="8033" lane="4" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-05-18" firstname="Agata" gender="F" lastname="Rompała" nation="POL" athleteid="4786">
              <RESULTS>
                <RESULT eventid="1140" points="625" reactiontime="+87" swimtime="00:11:16.11" resultid="4787" heatid="8712" lane="4" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:13.83" />
                    <SPLIT distance="150" swimtime="00:01:54.94" />
                    <SPLIT distance="200" swimtime="00:02:37.50" />
                    <SPLIT distance="250" swimtime="00:03:20.44" />
                    <SPLIT distance="300" swimtime="00:04:04.02" />
                    <SPLIT distance="350" swimtime="00:04:47.79" />
                    <SPLIT distance="400" swimtime="00:05:31.98" />
                    <SPLIT distance="450" swimtime="00:06:15.63" />
                    <SPLIT distance="500" swimtime="00:06:59.20" />
                    <SPLIT distance="550" swimtime="00:07:43.42" />
                    <SPLIT distance="600" swimtime="00:08:26.49" />
                    <SPLIT distance="650" swimtime="00:09:09.63" />
                    <SPLIT distance="700" swimtime="00:09:52.79" />
                    <SPLIT distance="750" swimtime="00:10:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" status="DNS" swimtime="00:00:00.00" resultid="4788" heatid="7760" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="4789" heatid="7804" lane="4" entrytime="00:01:05.00" />
                <RESULT eventid="1463" points="559" reactiontime="+90" swimtime="00:02:32.88" resultid="4790" heatid="7950" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="546" reactiontime="+92" swimtime="00:05:34.50" resultid="4791" heatid="9047" lane="3" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="150" swimtime="00:01:58.73" />
                    <SPLIT distance="200" swimtime="00:02:42.33" />
                    <SPLIT distance="250" swimtime="00:03:26.06" />
                    <SPLIT distance="300" swimtime="00:04:09.80" />
                    <SPLIT distance="350" swimtime="00:04:53.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-13" firstname="Karolina" gender="F" lastname="Rompała" nation="POL" athleteid="4792">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="4793" heatid="7717" lane="4" entrytime="00:02:50.00" />
                <RESULT eventid="1140" status="WDR" swimtime="00:00:00.00" resultid="4794" entrytime="00:10:50.00" />
                <RESULT eventid="1270" points="495" reactiontime="+78" swimtime="00:01:22.70" resultid="4795" heatid="7836" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="533" reactiontime="+82" swimtime="00:00:35.85" resultid="4796" heatid="7904" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="4797" heatid="7991" lane="7" entrytime="00:01:16.00" />
                <RESULT eventid="1687" points="530" reactiontime="+85" swimtime="00:05:30.83" resultid="4798" heatid="9048" lane="2" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                    <SPLIT distance="100" swimtime="00:01:15.43" />
                    <SPLIT distance="150" swimtime="00:01:56.42" />
                    <SPLIT distance="200" swimtime="00:02:39.00" />
                    <SPLIT distance="250" swimtime="00:03:22.28" />
                    <SPLIT distance="300" swimtime="00:04:05.81" />
                    <SPLIT distance="350" swimtime="00:04:49.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-11" firstname="Przemysław" gender="M" lastname="Jurek" nation="POL" athleteid="4799">
              <RESULTS>
                <RESULT eventid="1108" points="462" reactiontime="+77" swimtime="00:02:32.74" resultid="4800" heatid="7731" lane="8" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:09.83" />
                    <SPLIT distance="150" swimtime="00:01:57.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="576" swimtime="00:20:11.22" resultid="4801" heatid="8718" lane="1" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:13.37" />
                    <SPLIT distance="200" swimtime="00:02:30.98" />
                    <SPLIT distance="300" swimtime="00:03:50.77" />
                    <SPLIT distance="400" swimtime="00:05:12.71" />
                    <SPLIT distance="500" swimtime="00:06:33.58" />
                    <SPLIT distance="600" swimtime="00:07:54.10" />
                    <SPLIT distance="700" swimtime="00:09:16.02" />
                    <SPLIT distance="800" swimtime="00:10:38.45" />
                    <SPLIT distance="900" swimtime="00:12:00.63" />
                    <SPLIT distance="1000" swimtime="00:13:22.39" />
                    <SPLIT distance="1100" swimtime="00:14:34.34" />
                    <SPLIT distance="1200" swimtime="00:16:05.44" />
                    <SPLIT distance="1300" swimtime="00:17:28.03" />
                    <SPLIT distance="1400" swimtime="00:18:51.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="583" reactiontime="+68" swimtime="00:00:31.71" resultid="4802" heatid="7775" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1286" points="527" reactiontime="+79" swimtime="00:01:08.06" resultid="4803" heatid="7854" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="4804" heatid="8807" lane="6" entrytime="00:05:45.00" />
                <RESULT eventid="1703" points="552" reactiontime="+85" swimtime="00:04:52.87" resultid="4805" heatid="9060" lane="7" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:08.40" />
                    <SPLIT distance="150" swimtime="00:01:45.60" />
                    <SPLIT distance="200" swimtime="00:02:22.92" />
                    <SPLIT distance="250" swimtime="00:03:00.50" />
                    <SPLIT distance="300" swimtime="00:03:38.38" />
                    <SPLIT distance="350" swimtime="00:04:16.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Tarnowskie WOPR Masters B" number="1">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+73" swimtime="00:01:58.14" resultid="4812" heatid="7871" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:00.35" />
                    <SPLIT distance="150" swimtime="00:01:30.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4799" number="1" />
                    <RELAYPOSITION athleteid="4770" number="2" />
                    <RELAYPOSITION athleteid="4714" number="3" />
                    <RELAYPOSITION athleteid="4735" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" reactiontime="+89" swimtime="00:01:47.37" resultid="4813" heatid="7974" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.67" />
                    <SPLIT distance="100" swimtime="00:00:54.36" />
                    <SPLIT distance="150" swimtime="00:01:22.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4799" number="1" />
                    <RELAYPOSITION athleteid="4714" number="2" />
                    <RELAYPOSITION athleteid="4735" number="3" />
                    <RELAYPOSITION athleteid="4770" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Tarnowskie WOPR Masters C" number="2">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+64" swimtime="00:02:34.13" resultid="4814" heatid="7869" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                    <SPLIT distance="100" swimtime="00:01:28.63" />
                    <SPLIT distance="150" swimtime="00:01:59.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4762" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4746" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4773" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="4721" number="4" reactiontime="+93" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" reactiontime="+82" swimtime="00:02:11.83" resultid="4815" heatid="7971" lane="6" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:08.85" />
                    <SPLIT distance="150" swimtime="00:01:42.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4762" number="1" />
                    <RELAYPOSITION athleteid="4721" number="2" />
                    <RELAYPOSITION athleteid="4746" number="3" />
                    <RELAYPOSITION athleteid="4773" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" name="Tarnowskie WOPR Masters A" number="1">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)  (Czas: 14:21), na trzeciej zmianie" eventid="1334" reactiontime="+71" status="DSQ" swimtime="00:02:18.78" resultid="4810" heatid="7867" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:12.98" />
                    <SPLIT distance="150" swimtime="00:01:48.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4729" number="1" reactiontime="+71" status="DSQ" />
                    <RELAYPOSITION athleteid="4738" number="2" reactiontime="+80" status="DSQ" />
                    <RELAYPOSITION athleteid="4792" number="3" reactiontime="+64" status="DSQ" />
                    <RELAYPOSITION athleteid="4786" number="4" reactiontime="-7" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1495" reactiontime="+94" swimtime="00:02:04.66" resultid="4811" heatid="7969" lane="5" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:03.80" />
                    <SPLIT distance="150" swimtime="00:01:34.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4729" number="1" />
                    <RELAYPOSITION athleteid="4792" number="2" />
                    <RELAYPOSITION athleteid="4786" number="3" />
                    <RELAYPOSITION athleteid="4738" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="Tarnowskie WOPR Masters A" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+81" swimtime="00:01:59.80" resultid="4808" heatid="7736" lane="3" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="100" swimtime="00:00:59.75" />
                    <SPLIT distance="150" swimtime="00:01:32.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4773" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4729" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4792" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="4714" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" reactiontime="+75" swimtime="00:02:28.65" resultid="4809" heatid="8051" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:13.04" />
                    <SPLIT distance="150" swimtime="00:01:49.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4729" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4714" number="2" reactiontime="+89" />
                    <RELAYPOSITION athleteid="4792" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4757" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Tarnowskie WOPR Masters B" number="2">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+75" swimtime="00:01:56.45" resultid="4806" heatid="7736" lane="6" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="100" swimtime="00:00:58.96" />
                    <SPLIT distance="150" swimtime="00:01:29.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4735" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4738" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4786" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="4799" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" reactiontime="+78" swimtime="00:02:07.23" resultid="4807" heatid="8052" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:07.58" />
                    <SPLIT distance="150" swimtime="00:01:41.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4786" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4770" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="4738" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4799" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TOTOR" nation="POL" region="02" clubid="5564" name="Toruńczyk Masters Toruń">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1984-10-22" firstname="Magdalena" gender="F" lastname="Bolewska" nation="POL" athleteid="5565">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="5566" heatid="7683" lane="8" entrytime="00:00:29.56" />
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="5567" heatid="7718" lane="1" entrytime="00:02:48.50" />
                <RESULT eventid="1206" points="674" reactiontime="+90" swimtime="00:02:55.24" resultid="5568" heatid="7783" lane="5" entrytime="00:02:52.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:23.88" />
                    <SPLIT distance="150" swimtime="00:02:09.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="693" reactiontime="+88" swimtime="00:01:19.81" resultid="5569" heatid="7880" lane="3" entrytime="00:01:21.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="737" reactiontime="+88" swimtime="00:00:32.18" resultid="5570" heatid="7904" lane="3" entrytime="00:00:33.56" />
                <RESULT eventid="1574" points="605" reactiontime="+86" swimtime="00:01:15.62" resultid="5571" heatid="7990" lane="5" entrytime="00:01:18.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="648" reactiontime="+85" swimtime="00:00:36.49" resultid="5572" heatid="8028" lane="6" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="5573">
              <RESULTS>
                <RESULT eventid="1059" points="524" reactiontime="+78" swimtime="00:00:32.84" resultid="5574" heatid="7679" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1140" points="381" swimtime="00:12:35.51" resultid="5575" heatid="8713" lane="5" entrytime="00:12:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                    <SPLIT distance="100" swimtime="00:01:25.48" />
                    <SPLIT distance="200" swimtime="00:02:56.16" />
                    <SPLIT distance="300" swimtime="00:04:28.43" />
                    <SPLIT distance="400" swimtime="00:06:02.68" />
                    <SPLIT distance="500" swimtime="00:07:40.61" />
                    <SPLIT distance="600" swimtime="00:09:19.91" />
                    <SPLIT distance="700" swimtime="00:10:58.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="386" reactiontime="+84" swimtime="00:03:28.54" resultid="5576" heatid="7781" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.66" />
                    <SPLIT distance="100" swimtime="00:01:41.14" />
                    <SPLIT distance="150" swimtime="00:02:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="448" reactiontime="+78" swimtime="00:01:25.03" resultid="5577" heatid="7834" lane="1" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="395" reactiontime="+83" swimtime="00:01:37.46" resultid="5578" heatid="7875" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="400" reactiontime="+81" swimtime="00:02:47.14" resultid="5579" heatid="7949" lane="5" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:16.74" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="475" reactiontime="+86" swimtime="00:03:04.36" resultid="5580" heatid="8006" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:30.88" />
                    <SPLIT distance="150" swimtime="00:02:17.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" status="WDR" swimtime="00:00:00.00" resultid="5581" entrytime="00:05:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-14" firstname="Marta" gender="F" lastname="Lord" nation="POL" athleteid="5582">
              <RESULTS>
                <RESULT eventid="1092" points="691" reactiontime="+85" swimtime="00:02:41.77" resultid="5583" heatid="7717" lane="7" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:17.58" />
                    <SPLIT distance="150" swimtime="00:02:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="745" reactiontime="+75" swimtime="00:00:33.48" resultid="5584" heatid="7760" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1431" points="734" reactiontime="+84" swimtime="00:01:13.75" resultid="5585" heatid="7930" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="754" reactiontime="+85" swimtime="00:02:35.55" resultid="5586" heatid="8009" lane="4" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:16.37" />
                    <SPLIT distance="150" swimtime="00:01:56.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="5587">
              <RESULTS>
                <RESULT eventid="1108" points="335" reactiontime="+81" swimtime="00:02:50.06" resultid="5588" heatid="7725" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:21.68" />
                    <SPLIT distance="150" swimtime="00:02:11.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="5589" heatid="7863" lane="2" entrytime="00:03:05.00" />
                <RESULT eventid="1415" points="352" reactiontime="+77" swimtime="00:00:32.39" resultid="5590" heatid="7915" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1543" points="352" reactiontime="+96" swimtime="00:06:17.97" resultid="5591" heatid="8809" lane="8" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                    <SPLIT distance="100" swimtime="00:01:22.26" />
                    <SPLIT distance="200" swimtime="00:03:06.01" />
                    <SPLIT distance="250" swimtime="00:03:59.12" />
                    <SPLIT distance="300" swimtime="00:04:51.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="308" reactiontime="+90" swimtime="00:01:17.88" resultid="5592" heatid="7997" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="342" reactiontime="+88" swimtime="00:05:43.47" resultid="5593" heatid="9066" lane="4" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:19.70" />
                    <SPLIT distance="150" swimtime="00:02:02.81" />
                    <SPLIT distance="200" swimtime="00:02:46.22" />
                    <SPLIT distance="250" swimtime="00:03:31.39" />
                    <SPLIT distance="300" swimtime="00:04:15.75" />
                    <SPLIT distance="350" swimtime="00:05:00.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-03-24" firstname="Dariusz" gender="M" lastname="Pela" nation="POL" athleteid="5594">
              <RESULTS>
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="5595" heatid="7790" lane="1" entrytime="00:03:25.00" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="5596" heatid="7887" lane="6" entrytime="00:01:32.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="5597" heatid="8036" lane="7" entrytime="00:00:41.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-04" firstname="Karol" gender="M" lastname="Twarowski" nation="POL" athleteid="5598">
              <RESULTS>
                <RESULT eventid="1076" points="652" reactiontime="+74" swimtime="00:00:25.51" resultid="5599" heatid="7697" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1108" points="600" reactiontime="+81" swimtime="00:02:20.05" resultid="5600" heatid="7728" lane="1" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="657" reactiontime="+92" swimtime="00:02:41.64" resultid="5601" heatid="7784" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:02:00.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="667" reactiontime="+76" swimtime="00:00:56.12" resultid="5602" heatid="7817" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="723" reactiontime="+79" swimtime="00:01:04.13" resultid="5603" heatid="7937" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="678" reactiontime="+81" swimtime="00:05:03.93" resultid="5604" heatid="8812" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:09.18" />
                    <SPLIT distance="150" swimtime="00:01:48.61" />
                    <SPLIT distance="200" swimtime="00:02:27.62" />
                    <SPLIT distance="250" swimtime="00:03:11.14" />
                    <SPLIT distance="300" swimtime="00:03:54.64" />
                    <SPLIT distance="350" swimtime="00:04:31.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="568" reactiontime="+79" swimtime="00:02:20.79" resultid="5605" heatid="8010" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="150" swimtime="00:01:44.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="674" reactiontime="+81" swimtime="00:04:33.93" resultid="5606" heatid="9070" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                    <SPLIT distance="100" swimtime="00:01:02.24" />
                    <SPLIT distance="150" swimtime="00:01:35.70" />
                    <SPLIT distance="200" swimtime="00:02:10.16" />
                    <SPLIT distance="250" swimtime="00:02:45.29" />
                    <SPLIT distance="300" swimtime="00:03:21.68" />
                    <SPLIT distance="350" swimtime="00:03:58.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="5607">
              <RESULTS>
                <RESULT eventid="1190" points="96" reactiontime="+95" swimtime="00:01:12.30" resultid="5608" heatid="7763" lane="5" entrytime="00:01:06.41" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="5609" heatid="7839" lane="2" entrytime="00:01:57.54" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="5610" heatid="7859" lane="2" entrytime="00:05:19.20" />
                <RESULT eventid="1447" points="81" reactiontime="+93" swimtime="00:02:47.57" resultid="5611" heatid="7933" lane="8" entrytime="00:02:29.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="119" reactiontime="+117" swimtime="00:05:35.60" resultid="5612" heatid="8010" lane="2" entrytime="00:05:30.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.01" />
                    <SPLIT distance="100" swimtime="00:02:42.64" />
                    <SPLIT distance="150" swimtime="00:04:07.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="5613" entrytime="00:08:40.56" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="5614">
              <RESULTS>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="5615" heatid="7765" lane="7" entrytime="00:00:51.10" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="5616" heatid="7786" lane="1" entrytime="00:04:13.80" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="5617" heatid="7882" lane="6" entrytime="00:01:59.30" />
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="5618" heatid="7933" lane="6" entrytime="00:02:05.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="Osóbka" nation="POL" athleteid="5619">
              <RESULTS>
                <RESULT eventid="1254" points="91" reactiontime="+117" swimtime="00:02:39.89" resultid="5620" heatid="7806" lane="5" entrytime="00:02:50.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="5621" heatid="8030" lane="8" entrytime="00:01:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="5622">
              <RESULTS>
                <RESULT eventid="1190" points="174" reactiontime="+79" swimtime="00:01:02.04" resultid="5623" heatid="7764" lane="8" entrytime="00:00:58.52" />
                <RESULT eventid="1254" points="296" reactiontime="+125" swimtime="00:01:41.77" resultid="5624" heatid="7807" lane="2" entrytime="00:01:41.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="5625" heatid="7933" lane="7" entrytime="00:02:08.45" />
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="5626" heatid="8010" lane="3" entrytime="00:04:54.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-03" firstname="Artur" gender="M" lastname="Kłosiński" nation="POL" athleteid="5627">
              <RESULTS>
                <RESULT eventid="1076" points="555" reactiontime="+75" swimtime="00:00:26.92" resultid="5628" heatid="7689" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1108" points="427" reactiontime="+81" swimtime="00:02:36.78" resultid="5629" heatid="7729" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:58.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="484" reactiontime="+79" swimtime="00:02:58.90" resultid="5630" heatid="7793" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="150" swimtime="00:02:10.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="507" reactiontime="+77" swimtime="00:01:08.95" resultid="5631" heatid="7852" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="497" reactiontime="+71" swimtime="00:01:12.67" resultid="5632" heatid="7937" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="479" reactiontime="+83" swimtime="00:02:16.12" resultid="5633" heatid="7964" lane="8" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:05.95" />
                    <SPLIT distance="150" swimtime="00:01:41.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="401" reactiontime="+72" swimtime="00:02:38.13" resultid="5634" heatid="8015" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="5635" heatid="9062" lane="1" entrytime="00:05:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-16" firstname="Maciej" gender="M" lastname="Kujawa" nation="POL" athleteid="5636">
              <RESULTS>
                <RESULT eventid="1108" points="531" reactiontime="+97" swimtime="00:03:03.00" resultid="5637" heatid="7719" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:25.02" />
                    <SPLIT distance="150" swimtime="00:02:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="638" reactiontime="+88" swimtime="00:01:20.32" resultid="5638" heatid="7846" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="473" reactiontime="+93" swimtime="00:01:27.41" resultid="5639" heatid="7889" lane="2" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="475" reactiontime="+94" swimtime="00:00:39.09" resultid="5640" heatid="8038" lane="4" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Jarosław" gender="M" lastname="Wysocki" nation="POL" athleteid="5641">
              <RESULTS>
                <RESULT eventid="1222" points="571" reactiontime="+85" swimtime="00:03:30.84" resultid="5642" heatid="7788" lane="4" entrytime="00:03:32.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:39.77" />
                    <SPLIT distance="150" swimtime="00:02:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="549" reactiontime="+88" swimtime="00:01:35.41" resultid="5643" heatid="7887" lane="1" entrytime="00:01:33.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="537" reactiontime="+88" swimtime="00:00:41.58" resultid="5644" heatid="8036" lane="6" entrytime="00:00:41.37" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="5645">
              <RESULTS>
                <RESULT eventid="1076" points="646" reactiontime="+79" swimtime="00:00:31.22" resultid="5646" heatid="7695" lane="7" entrytime="00:00:31.08" />
                <RESULT eventid="1108" points="628" reactiontime="+91" swimtime="00:03:11.73" resultid="5647" heatid="7723" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="100" swimtime="00:01:35.10" />
                    <SPLIT distance="150" swimtime="00:02:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="569" reactiontime="+83" swimtime="00:01:12.23" resultid="5648" heatid="7811" lane="4" entrytime="00:01:12.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="654" reactiontime="+79" swimtime="00:01:23.43" resultid="5649" heatid="7845" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="602" reactiontime="+77" swimtime="00:00:35.45" resultid="5650" heatid="7914" lane="8" entrytime="00:00:34.50" />
                <RESULT eventid="1543" points="516" reactiontime="+88" swimtime="00:07:14.90" resultid="5651" heatid="8810" lane="7" entrytime="00:07:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:36.71" />
                    <SPLIT distance="150" swimtime="00:02:38.77" />
                    <SPLIT distance="200" swimtime="00:03:41.34" />
                    <SPLIT distance="250" swimtime="00:04:40.46" />
                    <SPLIT distance="300" swimtime="00:05:41.07" />
                    <SPLIT distance="350" swimtime="00:06:30.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="520" reactiontime="+83" swimtime="00:01:24.91" resultid="5652" heatid="7996" lane="7" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="Szufarski" nation="POL" athleteid="5653">
              <RESULTS>
                <RESULT eventid="1108" points="470" reactiontime="+105" swimtime="00:03:31.17" resultid="5654" heatid="7721" lane="5" entrytime="00:03:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:38.97" />
                    <SPLIT distance="150" swimtime="00:02:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="422" reactiontime="+109" swimtime="00:03:53.21" resultid="5655" heatid="7787" lane="7" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.89" />
                    <SPLIT distance="100" swimtime="00:01:50.06" />
                    <SPLIT distance="150" swimtime="00:02:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="438" reactiontime="+102" swimtime="00:01:35.39" resultid="5656" heatid="7841" lane="7" entrytime="00:01:37.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="418" reactiontime="+107" swimtime="00:01:44.46" resultid="5657" heatid="7885" lane="5" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="389" reactiontime="+106" swimtime="00:07:57.88" resultid="5658" heatid="8812" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:51.42" />
                    <SPLIT distance="150" swimtime="00:02:57.56" />
                    <SPLIT distance="200" swimtime="00:04:00.49" />
                    <SPLIT distance="250" swimtime="00:05:01.72" />
                    <SPLIT distance="300" swimtime="00:06:05.92" />
                    <SPLIT distance="350" swimtime="00:07:03.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="302" reactiontime="+108" swimtime="00:01:41.76" resultid="5659" heatid="7994" lane="2" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="391" reactiontime="+99" swimtime="00:00:46.20" resultid="5660" heatid="8032" lane="1" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="M" name="Toruńczyk Masters Toruń F" number="2">
              <RESULTS>
                <RESULT eventid="1357" status="WDR" swimtime="00:00:00.00" resultid="5665" entrytime="00:03:55.40">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5614" number="1" />
                    <RELAYPOSITION athleteid="5619" number="2" />
                    <RELAYPOSITION athleteid="5607" number="3" />
                    <RELAYPOSITION athleteid="5622" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="5666" heatid="7970" lane="7" entrytime="00:03:10.20">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5614" number="1" />
                    <RELAYPOSITION athleteid="5619" number="2" />
                    <RELAYPOSITION athleteid="5607" number="3" />
                    <RELAYPOSITION athleteid="5622" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Toruńczyk Masters Toruń E" number="3">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+88" swimtime="00:02:36.80" resultid="5663" heatid="7869" lane="5" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                    <SPLIT distance="100" swimtime="00:01:29.21" />
                    <SPLIT distance="150" swimtime="00:02:05.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5653" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="5641" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="5636" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="5645" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="5664" heatid="7970" lane="3" entrytime="00:02:19.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5636" number="1" />
                    <RELAYPOSITION athleteid="5641" number="2" />
                    <RELAYPOSITION athleteid="5653" number="3" />
                    <RELAYPOSITION athleteid="5645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Toruńczyk Masters Toruń B" number="4">
              <RESULTS>
                <RESULT eventid="1357" status="WDR" swimtime="00:00:00.00" resultid="5667" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5627" number="1" />
                    <RELAYPOSITION athleteid="5594" number="2" />
                    <RELAYPOSITION athleteid="5587" number="3" />
                    <RELAYPOSITION athleteid="5598" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Toruńczyk Masters Toruń B" number="1">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="5661" heatid="7737" lane="3" entrytime="00:01:56.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5565" number="1" />
                    <RELAYPOSITION athleteid="5582" number="2" />
                    <RELAYPOSITION athleteid="5627" number="3" />
                    <RELAYPOSITION athleteid="5598" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" reactiontime="+76" swimtime="00:02:05.26" resultid="5662" heatid="8052" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:10.32" />
                    <SPLIT distance="150" swimtime="00:01:38.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5582" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="5565" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="5627" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="5598" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="5455" name="UKP Masters Unia Oświęcim" shortname="Masters Unia Oświęcim">
          <ATHLETES>
            <ATHLETE birthdate="1961-03-16" firstname="Tomasz" gender="M" lastname="Dorywalski" nation="POL" athleteid="5476">
              <RESULTS>
                <RESULT eventid="1190" points="542" reactiontime="+65" swimtime="00:00:36.02" resultid="5477" heatid="7770" lane="3" entrytime="00:00:38.50" />
                <RESULT eventid="1447" points="549" reactiontime="+69" swimtime="00:01:19.16" resultid="5478" heatid="7938" lane="7" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="542" reactiontime="+71" swimtime="00:02:57.75" resultid="5479" heatid="8015" lane="8" entrytime="00:02:58.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:23.94" />
                    <SPLIT distance="150" swimtime="00:02:10.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-27" firstname="Robert" gender="M" lastname="Krulikowski" nation="POL" athleteid="5480">
              <RESULTS>
                <RESULT eventid="1286" points="612" reactiontime="+95" swimtime="00:01:10.44" resultid="5481" heatid="7854" lane="4" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="531" reactiontime="+93" swimtime="00:00:31.03" resultid="5482" heatid="7920" lane="5" entrytime="00:00:29.50" />
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5492" heatid="7703" lane="5" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-10" firstname="Jolanta" gender="F" lastname="Płatek" nation="POL" athleteid="5483">
              <RESULTS>
                <RESULT eventid="1270" points="488" reactiontime="+98" swimtime="00:01:26.54" resultid="5484" heatid="7829" lane="3" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="542" reactiontime="+78" swimtime="00:01:23.31" resultid="5485" heatid="7928" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="476" reactiontime="+96" swimtime="00:05:54.48" resultid="5486" heatid="9051" lane="6" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                    <SPLIT distance="150" swimtime="00:02:05.94" />
                    <SPLIT distance="200" swimtime="00:02:51.28" />
                    <SPLIT distance="250" swimtime="00:03:37.24" />
                    <SPLIT distance="300" swimtime="00:04:23.51" />
                    <SPLIT distance="350" swimtime="00:05:10.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="651" reactiontime="+75" swimtime="00:00:36.49" resultid="5493" heatid="7759" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-03" firstname="Ilona" gender="F" lastname="Szkudlarz" nation="POL" athleteid="5487">
              <RESULTS>
                <RESULT eventid="1059" points="496" reactiontime="+94" swimtime="00:00:35.08" resultid="5488" heatid="7678" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1173" points="478" reactiontime="+81" swimtime="00:00:41.67" resultid="5489" heatid="7757" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1639" points="528" reactiontime="+84" swimtime="00:00:43.83" resultid="5490" heatid="8026" lane="7" entrytime="00:00:44.10" />
                <RESULT eventid="1366" points="543" reactiontime="+91" swimtime="00:01:36.67" resultid="6469" heatid="7877" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Masters Unia Oświęcim C">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+77" swimtime="00:02:23.72" resultid="5491" heatid="8050" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:20.29" />
                    <SPLIT distance="150" swimtime="00:01:51.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5483" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="5487" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="5480" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="5476" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="04514" nation="POL" region="14" clubid="2380" name="UKS 307 Warszawa">
          <CONTACT name="Ilczyszyn" />
          <ATHLETES>
            <ATHLETE birthdate="1983-07-13" firstname="Krzysztof" gender="M" lastname="Ilczyszyn" nation="POL" athleteid="2388">
              <RESULTS>
                <RESULT eventid="1254" points="479" reactiontime="+88" swimtime="00:01:02.67" resultid="2389" heatid="7819" lane="7" entrytime="00:01:02.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="399" reactiontime="+86" swimtime="00:01:14.66" resultid="2390" heatid="7850" lane="3" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="403" reactiontime="+87" swimtime="00:00:30.96" resultid="2391" heatid="7919" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1479" points="385" reactiontime="+90" swimtime="00:02:26.39" resultid="2392" heatid="7961" lane="4" entrytime="00:02:27.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="150" swimtime="00:01:51.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="409" reactiontime="+87" swimtime="00:01:10.90" resultid="2393" heatid="7998" lane="1" entrytime="00:01:15.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="424" reactiontime="+84" swimtime="00:05:19.61" resultid="2394" heatid="9064" lane="8" entrytime="00:05:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:54.01" />
                    <SPLIT distance="200" swimtime="00:02:35.38" />
                    <SPLIT distance="250" swimtime="00:03:17.62" />
                    <SPLIT distance="300" swimtime="00:03:59.89" />
                    <SPLIT distance="350" swimtime="00:04:40.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-03" firstname="Damian" gender="M" lastname="Ziółkowski" nation="POL" athleteid="2395">
              <RESULTS>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="2396" heatid="7770" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="2397" heatid="7819" lane="2" entrytime="00:01:02.63" />
                <RESULT eventid="1415" points="594" reactiontime="+86" swimtime="00:00:30.52" resultid="2398" heatid="7919" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1479" points="505" reactiontime="+85" swimtime="00:02:19.96" resultid="2399" heatid="7961" lane="5" entrytime="00:02:27.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:44.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="413" reactiontime="+85" swimtime="00:01:16.34" resultid="2400" heatid="7998" lane="7" entrytime="00:01:15.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="483" reactiontime="+90" swimtime="00:05:08.81" resultid="2401" heatid="9064" lane="1" entrytime="00:05:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:12.38" />
                    <SPLIT distance="150" swimtime="00:01:52.42" />
                    <SPLIT distance="200" swimtime="00:02:33.34" />
                    <SPLIT distance="250" swimtime="00:03:13.79" />
                    <SPLIT distance="300" swimtime="00:03:54.95" />
                    <SPLIT distance="350" swimtime="00:04:33.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="08" clubid="2925" name="UKS Delfin Masters Tarnobrzeg" shortname="Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1977-04-24" firstname="Renata" gender="F" lastname="Osmala" nation="POL" athleteid="2926">
              <RESULTS>
                <RESULT eventid="1173" points="675" reactiontime="+62" swimtime="00:00:36.34" resultid="2927" heatid="7759" lane="2" entrytime="00:00:37.70" />
                <RESULT eventid="1270" points="635" reactiontime="+82" swimtime="00:01:18.99" resultid="2928" heatid="7834" lane="6" entrytime="00:01:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="649" reactiontime="+83" swimtime="00:01:25.28" resultid="2929" heatid="7879" lane="8" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="584" reactiontime="+65" swimtime="00:01:18.87" resultid="2930" heatid="7930" lane="2" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="592" reactiontime="+73" swimtime="00:02:49.99" resultid="2931" heatid="8008" lane="2" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                    <SPLIT distance="100" swimtime="00:01:22.59" />
                    <SPLIT distance="150" swimtime="00:02:06.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="629" reactiontime="+82" swimtime="00:00:39.55" resultid="2932" heatid="8027" lane="1" entrytime="00:00:41.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="2933">
              <RESULTS>
                <RESULT eventid="1059" points="627" reactiontime="+77" swimtime="00:00:31.73" resultid="2934" heatid="7680" lane="3" entrytime="00:00:32.34" />
                <RESULT eventid="1238" points="544" reactiontime="+77" swimtime="00:01:10.75" resultid="2935" heatid="7803" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="613" reactiontime="+79" swimtime="00:01:19.92" resultid="2936" heatid="7834" lane="5" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="510" reactiontime="+82" swimtime="00:00:36.94" resultid="2937" heatid="7902" lane="1" entrytime="00:00:37.23" />
                <RESULT eventid="1574" points="487" reactiontime="+84" swimtime="00:01:23.05" resultid="2938" heatid="7989" lane="4" entrytime="00:01:25.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="587" reactiontime="+83" swimtime="00:00:40.46" resultid="2939" heatid="8027" lane="8" entrytime="00:00:41.68" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="2940">
              <RESULTS>
                <RESULT eventid="1059" points="619" reactiontime="+79" swimtime="00:00:31.86" resultid="2941" heatid="7680" lane="4" entrytime="00:00:32.10" />
                <RESULT eventid="1238" points="536" reactiontime="+80" swimtime="00:01:11.11" resultid="2942" heatid="7803" lane="6" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="573" reactiontime="+80" swimtime="00:01:21.73" resultid="2943" heatid="7833" lane="4" entrytime="00:01:23.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="486" reactiontime="+85" swimtime="00:00:37.54" resultid="2944" heatid="7901" lane="7" entrytime="00:00:38.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-08-01" firstname="Monika" gender="F" lastname="Maciąg" nation="POL" athleteid="2945">
              <RESULTS>
                <RESULT eventid="1059" points="518" reactiontime="+92" swimtime="00:00:33.84" resultid="2946" heatid="7678" lane="3" entrytime="00:00:34.84" />
                <RESULT eventid="1173" points="477" reactiontime="+75" swimtime="00:00:40.48" resultid="2947" heatid="7757" lane="8" entrytime="00:00:43.89" />
                <RESULT eventid="1270" points="487" reactiontime="+93" swimtime="00:01:26.58" resultid="2948" heatid="7831" lane="3" entrytime="00:01:29.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="491" reactiontime="+83" swimtime="00:01:26.14" resultid="2949" heatid="7929" lane="8" entrytime="00:01:29.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="534" reactiontime="+79" swimtime="00:03:04.14" resultid="2950" heatid="8007" lane="7" entrytime="00:03:14.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                    <SPLIT distance="100" swimtime="00:01:31.15" />
                    <SPLIT distance="150" swimtime="00:02:18.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-06-15" firstname="Anna" gender="F" lastname="Buczek" nation="POL" athleteid="2951">
              <RESULTS>
                <RESULT eventid="1059" points="353" reactiontime="+109" swimtime="00:00:38.43" resultid="2952" heatid="7674" lane="4" entrytime="00:00:40.32" />
                <RESULT eventid="1366" points="414" reactiontime="+101" swimtime="00:01:41.55" resultid="2953" heatid="7876" lane="5" entrytime="00:01:47.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="396" reactiontime="+94" swimtime="00:00:46.74" resultid="2954" heatid="8025" lane="8" entrytime="00:00:46.30" />
                <RESULT eventid="1238" points="342" reactiontime="+104" swimtime="00:01:24.91" resultid="3525" heatid="7799" lane="8" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Beata" gender="F" lastname="Kaczmarczyk" nation="POL" athleteid="2955">
              <RESULTS>
                <RESULT eventid="1059" points="479" reactiontime="+92" swimtime="00:00:34.69" resultid="2956" heatid="7677" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1238" points="418" reactiontime="+85" swimtime="00:01:17.25" resultid="2957" heatid="7801" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="421" reactiontime="+88" swimtime="00:02:50.85" resultid="2958" heatid="7947" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:21.64" />
                    <SPLIT distance="150" swimtime="00:02:07.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-07" firstname="Albert" gender="M" lastname="Szwajkowski" nation="POL" athleteid="2959">
              <RESULTS>
                <RESULT eventid="1076" points="474" reactiontime="+105" swimtime="00:00:30.46" resultid="2960" heatid="7697" lane="8" entrytime="00:00:30.28" />
                <RESULT eventid="1286" points="427" reactiontime="+79" swimtime="00:01:19.43" resultid="2961" heatid="7847" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="413" reactiontime="+87" swimtime="00:00:33.74" resultid="2962" heatid="7914" lane="4" entrytime="00:00:33.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="2963">
              <RESULTS>
                <RESULT eventid="1076" points="653" reactiontime="+78" swimtime="00:00:27.34" resultid="2964" heatid="7706" lane="1" entrytime="00:00:27.45" />
                <RESULT eventid="1254" points="591" reactiontime="+79" swimtime="00:01:01.28" resultid="2965" heatid="7820" lane="6" entrytime="00:01:01.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="542" reactiontime="+79" swimtime="00:01:12.41" resultid="2966" heatid="7849" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="599" reactiontime="+74" swimtime="00:00:30.44" resultid="2967" heatid="7917" lane="1" entrytime="00:00:31.39" />
                <RESULT eventid="1479" points="489" reactiontime="+84" swimtime="00:02:21.48" resultid="2968" heatid="7962" lane="5" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:06.73" />
                    <SPLIT distance="150" swimtime="00:01:44.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-21" firstname="Piotr" gender="M" lastname="Zawół" nation="POL" athleteid="2969">
              <RESULTS>
                <RESULT eventid="1076" points="568" reactiontime="+82" swimtime="00:00:28.64" resultid="2970" heatid="7703" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1318" points="404" reactiontime="+85" swimtime="00:02:51.30" resultid="2971" heatid="7864" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:18.48" />
                    <SPLIT distance="150" swimtime="00:02:05.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="466" reactiontime="+86" swimtime="00:01:13.33" resultid="2972" heatid="8000" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="2973">
              <RESULTS>
                <RESULT eventid="1076" points="462" reactiontime="+83" swimtime="00:00:30.68" resultid="2974" heatid="7695" lane="8" entrytime="00:00:31.25" />
                <RESULT eventid="1254" points="409" reactiontime="+81" swimtime="00:01:09.28" resultid="2975" heatid="7811" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="385" reactiontime="+82" swimtime="00:02:33.22" resultid="2976" heatid="7959" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="150" swimtime="00:01:54.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="378" reactiontime="+84" swimtime="00:05:34.89" resultid="2977" heatid="9065" lane="7" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:01.48" />
                    <SPLIT distance="200" swimtime="00:02:43.83" />
                    <SPLIT distance="250" swimtime="00:03:26.59" />
                    <SPLIT distance="300" swimtime="00:04:09.88" />
                    <SPLIT distance="350" swimtime="00:04:53.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-13" firstname="Rafał" gender="M" lastname="Woźniak" nation="POL" athleteid="2978">
              <RESULTS>
                <RESULT eventid="1156" points="322" swimtime="00:24:13.96" resultid="2979" heatid="8722" lane="5" entrytime="00:25:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:23.61" />
                    <SPLIT distance="200" swimtime="00:02:58.00" />
                    <SPLIT distance="300" swimtime="00:04:32.31" />
                    <SPLIT distance="400" swimtime="00:06:08.14" />
                    <SPLIT distance="500" swimtime="00:07:45.93" />
                    <SPLIT distance="600" swimtime="00:09:24.37" />
                    <SPLIT distance="700" swimtime="00:11:03.69" />
                    <SPLIT distance="800" swimtime="00:12:42.51" />
                    <SPLIT distance="900" swimtime="00:14:21.34" />
                    <SPLIT distance="1000" swimtime="00:16:01.54" />
                    <SPLIT distance="1100" swimtime="00:17:42.08" />
                    <SPLIT distance="1200" swimtime="00:19:21.43" />
                    <SPLIT distance="1300" swimtime="00:21:01.09" />
                    <SPLIT distance="1400" swimtime="00:22:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="383" reactiontime="+99" swimtime="00:03:16.59" resultid="2980" heatid="7793" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.98" />
                    <SPLIT distance="100" swimtime="00:01:33.73" />
                    <SPLIT distance="150" swimtime="00:02:25.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="299" reactiontime="+95" swimtime="00:05:59.64" resultid="2981" heatid="9065" lane="1" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:06.36" />
                    <SPLIT distance="200" swimtime="00:02:52.94" />
                    <SPLIT distance="250" swimtime="00:03:40.08" />
                    <SPLIT distance="300" swimtime="00:04:28.04" />
                    <SPLIT distance="350" swimtime="00:05:15.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="Szklarz" nation="POL" athleteid="2982">
              <RESULTS>
                <RESULT eventid="1076" points="547" reactiontime="+73" swimtime="00:00:28.99" resultid="2983" heatid="7704" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1286" points="443" reactiontime="+70" swimtime="00:01:17.44" resultid="2984" heatid="7851" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="458" reactiontime="+74" swimtime="00:01:23.05" resultid="2985" heatid="7892" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="508" reactiontime="+73" swimtime="00:00:36.18" resultid="2986" heatid="8042" lane="6" entrytime="00:00:36.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-15" firstname="Paweł" gender="M" lastname="Nowak" nation="POL" athleteid="2987">
              <RESULTS>
                <RESULT eventid="1190" points="404" reactiontime="+63" swimtime="00:00:36.69" resultid="2988" heatid="7772" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1447" points="389" reactiontime="+65" swimtime="00:01:20.93" resultid="2989" heatid="7938" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-17" firstname="Sławek" gender="M" lastname="Kowalski" nation="POL" athleteid="2990">
              <RESULTS>
                <RESULT eventid="1286" points="486" reactiontime="+80" swimtime="00:01:16.05" resultid="2991" heatid="7846" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="568" reactiontime="+85" swimtime="00:00:35.60" resultid="2992" heatid="8042" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-09-08" firstname="Patrycja" gender="F" lastname="Urbaniak" nation="POL" athleteid="2993">
              <RESULTS>
                <RESULT eventid="1059" points="676" reactiontime="+74" swimtime="00:00:30.17" resultid="2994" heatid="7682" lane="4" entrytime="00:00:29.60" />
                <RESULT eventid="1238" points="649" reactiontime="+76" swimtime="00:01:06.83" resultid="2995" heatid="7804" lane="5" entrytime="00:01:05.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="606" reactiontime="+73" swimtime="00:01:16.90" resultid="2996" heatid="7836" lane="6" entrytime="00:01:16.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="620" reactiontime="+76" swimtime="00:00:33.57" resultid="2997" heatid="7904" lane="5" entrytime="00:00:33.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-15" firstname="Andrzej" gender="M" lastname="Brożyna" nation="POL" athleteid="3526">
              <RESULTS>
                <RESULT eventid="1076" points="507" reactiontime="+70" swimtime="00:00:27.74" resultid="3527" heatid="7697" lane="7" entrytime="00:00:30.15" />
                <RESULT eventid="1415" points="328" reactiontime="+82" swimtime="00:00:33.13" resultid="3528" heatid="7916" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1190" points="497" reactiontime="+57" swimtime="00:00:33.44" resultid="3529" heatid="7772" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="3530" heatid="8037" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Delfin Masters Tarnobrzeg C" number="1">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+76" swimtime="00:01:54.96" resultid="3003" heatid="7972" lane="6" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                    <SPLIT distance="100" swimtime="00:00:57.93" />
                    <SPLIT distance="150" swimtime="00:01:27.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2982" number="1" />
                    <RELAYPOSITION athleteid="2990" number="2" />
                    <RELAYPOSITION athleteid="2959" number="3" />
                    <RELAYPOSITION athleteid="2963" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Delfin Masters Tarnobrzeg B">
              <RESULTS>
                <RESULT eventid="1334" reactiontime="+81" swimtime="00:02:27.74" resultid="3001" heatid="7867" lane="7" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                    <SPLIT distance="150" swimtime="00:01:56.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2945" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2926" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2933" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2940" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1495" reactiontime="+76" swimtime="00:02:09.98" resultid="3002" heatid="7969" lane="2" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:04.42" />
                    <SPLIT distance="150" swimtime="00:01:38.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2933" number="1" />
                    <RELAYPOSITION athleteid="2926" number="2" />
                    <RELAYPOSITION athleteid="2945" number="3" />
                    <RELAYPOSITION athleteid="2940" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Delfin Masters Tarnobrzeg B">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+78" swimtime="00:01:58.27" resultid="2998" heatid="7737" lane="7" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                    <SPLIT distance="150" swimtime="00:01:26.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2933" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="2982" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="2963" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2940" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1671" reactiontime="+75" swimtime="00:02:16.29" resultid="3000" heatid="8051" lane="3" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                    <SPLIT distance="150" swimtime="00:01:48.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2926" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="2933" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2982" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="2963" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Delfin Masters Tarnobrzeg C" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+81" swimtime="00:02:04.99" resultid="2999" heatid="7736" lane="4" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:02.95" />
                    <SPLIT distance="150" swimtime="00:01:33.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2990" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2945" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="2959" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="2926" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="04111" nation="POL" region="11" clubid="2768" name="UKS Delfinek Częstochowa" shortname="Delfinek Częstochowa">
          <CONTACT city="Częstochowa" email="uksdelfinek@op.pl" internet="ww.uksdelinek.pl" name="Langier Wojciech" phone="504940294" state="ŚŁĄSK" street="Niepodległości 20/22" zip="42-200" />
          <ATHLETES>
            <ATHLETE birthdate="1969-06-21" firstname="Jacek" gender="M" lastname="Drzewiecki" nation="POL" athleteid="2769">
              <RESULTS>
                <RESULT eventid="1286" points="493" reactiontime="+84" swimtime="00:01:15.68" resultid="2770" heatid="7849" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03801" nation="POL" region="01" clubid="5079" name="UKS Delfinek Legnica" shortname="Delfinek Legnica">
          <CONTACT email="jmalchar@o2.pl" name="Malchar" phone="506034671" />
          <ATHLETES>
            <ATHLETE birthdate="1971-04-11" firstname="Sebastian" gender="M" lastname="Hudyka" nation="POL" athleteid="5094">
              <RESULTS>
                <RESULT eventid="1156" points="351" swimtime="00:23:32.58" resultid="5095" heatid="8721" lane="4" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="200" swimtime="00:02:55.14" />
                    <SPLIT distance="300" swimtime="00:04:27.14" />
                    <SPLIT distance="400" swimtime="00:05:59.79" />
                    <SPLIT distance="500" swimtime="00:07:34.28" />
                    <SPLIT distance="600" swimtime="00:09:09.09" />
                    <SPLIT distance="700" swimtime="00:10:43.98" />
                    <SPLIT distance="800" swimtime="00:12:19.96" />
                    <SPLIT distance="900" swimtime="00:13:56.47" />
                    <SPLIT distance="1000" swimtime="00:15:33.87" />
                    <SPLIT distance="1100" swimtime="00:17:10.41" />
                    <SPLIT distance="1200" swimtime="00:18:47.42" />
                    <SPLIT distance="1300" swimtime="00:20:23.49" />
                    <SPLIT distance="1400" swimtime="00:22:00.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="339" reactiontime="+91" swimtime="00:05:45.00" resultid="5096" heatid="9066" lane="3" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="150" swimtime="00:02:05.00" />
                    <SPLIT distance="200" swimtime="00:02:49.46" />
                    <SPLIT distance="250" swimtime="00:03:34.23" />
                    <SPLIT distance="300" swimtime="00:04:18.80" />
                    <SPLIT distance="350" swimtime="00:05:03.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-12-28" firstname="Jowita" gender="F" lastname="Malchar" nation="POL" athleteid="5097">
              <RESULTS>
                <RESULT eventid="1059" points="625" reactiontime="+83" swimtime="00:00:30.56" resultid="5098" heatid="7681" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1092" points="593" reactiontime="+80" swimtime="00:02:50.20" resultid="5099" heatid="7716" lane="4" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:18.49" />
                    <SPLIT distance="150" swimtime="00:02:08.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="553" reactiontime="+81" swimtime="00:03:10.25" resultid="5100" heatid="7782" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:01:28.93" />
                    <SPLIT distance="150" swimtime="00:02:19.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="579" reactiontime="+74" swimtime="00:01:18.10" resultid="5101" heatid="7835" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="586" reactiontime="+71" swimtime="00:01:26.84" resultid="5102" heatid="7879" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="577" reactiontime="+90" swimtime="00:06:05.65" resultid="5103" heatid="8802" lane="3" entrytime="00:06:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                    <SPLIT distance="100" swimtime="00:01:22.58" />
                    <SPLIT distance="150" swimtime="00:02:08.99" />
                    <SPLIT distance="200" swimtime="00:02:55.35" />
                    <SPLIT distance="250" swimtime="00:03:48.11" />
                    <SPLIT distance="300" swimtime="00:04:40.39" />
                    <SPLIT distance="350" swimtime="00:05:24.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="540" reactiontime="+79" swimtime="00:01:18.32" resultid="5104" heatid="7990" lane="1" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="518" reactiontime="+79" swimtime="00:05:40.39" resultid="5105" heatid="9048" lane="8" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:17.83" />
                    <SPLIT distance="150" swimtime="00:02:01.23" />
                    <SPLIT distance="200" swimtime="00:03:30.21" />
                    <SPLIT distance="250" swimtime="00:04:14.84" />
                    <SPLIT distance="300" swimtime="00:04:59.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-11-28" firstname="Anna" gender="F" lastname="Sołtys" nation="POL" athleteid="5106">
              <RESULTS>
                <RESULT eventid="1059" points="183" reactiontime="+132" swimtime="00:00:46.58" resultid="5107" heatid="7673" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1206" points="223" swimtime="00:04:10.21" resultid="5108" heatid="7780" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.95" />
                    <SPLIT distance="100" swimtime="00:01:56.40" />
                    <SPLIT distance="150" swimtime="00:03:02.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="161" reactiontime="+100" swimtime="00:01:46.16" resultid="5109" heatid="7798" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="187" reactiontime="+96" swimtime="00:02:04.97" resultid="5110" heatid="7875" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="130" reactiontime="+100" swimtime="00:04:02.62" resultid="5111" heatid="7945" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.40" />
                    <SPLIT distance="100" swimtime="00:01:53.04" />
                    <SPLIT distance="150" swimtime="00:03:00.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="215" reactiontime="+96" swimtime="00:00:54.81" resultid="5112" heatid="8024" lane="3" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-10" firstname="Radosław" gender="M" lastname="Wirszuło" nation="POL" athleteid="5113">
              <RESULTS>
                <RESULT eventid="1076" points="428" reactiontime="+104" swimtime="00:00:30.30" resultid="5114" heatid="7692" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1190" points="250" reactiontime="+76" swimtime="00:00:39.75" resultid="5115" heatid="7770" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1254" points="330" reactiontime="+96" swimtime="00:01:10.25" resultid="5116" heatid="7813" lane="8" entrytime="00:01:12.00" />
                <RESULT eventid="1415" points="255" reactiontime="+86" swimtime="00:00:37.34" resultid="5117" heatid="7911" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1447" points="246" reactiontime="+81" swimtime="00:01:27.82" resultid="5118" heatid="7937" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="307" reactiontime="+104" swimtime="00:06:02.37" resultid="5119" heatid="9067" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="150" swimtime="00:02:01.57" />
                    <SPLIT distance="200" swimtime="00:02:48.50" />
                    <SPLIT distance="250" swimtime="00:03:37.58" />
                    <SPLIT distance="300" swimtime="00:04:27.08" />
                    <SPLIT distance="350" swimtime="00:05:16.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="01" clubid="3273" name="UKS Energetyk Zgorzelec" shortname="Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="andrzejdaszynski@tlen.pl" name="Daszyński Andrzej" phone="607151541" state="DOL" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="3289">
              <RESULTS>
                <RESULT eventid="1108" points="322" reactiontime="+93" swimtime="00:03:55.59" resultid="3290" heatid="7720" lane="4" entrytime="00:04:03.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.16" />
                    <SPLIT distance="100" swimtime="00:01:53.51" />
                    <SPLIT distance="150" swimtime="00:03:03.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="3291" heatid="8724" lane="1" entrytime="00:35:00.00" entrycourse="SCM" />
                <RESULT eventid="1190" points="326" reactiontime="+79" swimtime="00:00:48.41" resultid="3292" heatid="7765" lane="4" entrytime="00:00:49.00" entrycourse="SCM" />
                <RESULT eventid="1318" points="264" reactiontime="+95" swimtime="00:04:20.73" resultid="3293" heatid="7860" lane="8" entrytime="00:04:29.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.29" />
                    <SPLIT distance="100" swimtime="00:02:01.98" />
                    <SPLIT distance="150" swimtime="00:03:12.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="321" reactiontime="+78" swimtime="00:01:45.68" resultid="3294" heatid="7934" lane="6" entrytime="00:01:50.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="384" reactiontime="+95" swimtime="00:08:26.43" resultid="3295" heatid="8811" lane="1" entrytime="00:08:38.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.87" />
                    <SPLIT distance="100" swimtime="00:02:01.85" />
                    <SPLIT distance="150" swimtime="00:03:05.38" />
                    <SPLIT distance="200" swimtime="00:04:06.01" />
                    <SPLIT distance="250" swimtime="00:05:18.26" />
                    <SPLIT distance="300" swimtime="00:06:28.71" />
                    <SPLIT distance="350" swimtime="00:07:26.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="316" reactiontime="+84" swimtime="00:03:51.38" resultid="3296" heatid="8012" lane="8" entrytime="00:03:55.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.64" />
                    <SPLIT distance="100" swimtime="00:01:54.30" />
                    <SPLIT distance="150" swimtime="00:02:54.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="292" reactiontime="+101" swimtime="00:07:42.69" resultid="3297" heatid="9070" lane="4" entrytime="00:07:38.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.88" />
                    <SPLIT distance="100" swimtime="00:01:48.35" />
                    <SPLIT distance="150" swimtime="00:02:50.30" />
                    <SPLIT distance="200" swimtime="00:03:51.42" />
                    <SPLIT distance="250" swimtime="00:04:50.42" />
                    <SPLIT distance="300" swimtime="00:05:48.44" />
                    <SPLIT distance="350" swimtime="00:06:47.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05114" nation="POL" region="14" clubid="6390" name="UKS G-8 Bielany Warszawa" shortname="G-8 Bielany Warszawa">
          <CONTACT name="Michał Choiński" phone="783753723" />
          <ATHLETES>
            <ATHLETE birthdate="1990-06-24" firstname="Michał" gender="M" lastname="Choiński" nation="POL" license="105114200075" athleteid="6391">
              <RESULTS>
                <RESULT eventid="1254" points="775" reactiontime="+69" swimtime="00:00:55.43" resultid="6392" heatid="7825" lane="3" entrytime="00:00:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="696" reactiontime="+74" swimtime="00:01:04.81" resultid="6393" heatid="7856" lane="3" entrytime="00:01:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="916" reactiontime="+71" swimtime="00:00:25.73" resultid="6394" heatid="7925" lane="5" entrytime="00:00:25.80" entrycourse="SCM" />
                <RESULT eventid="1591" points="690" reactiontime="+74" swimtime="00:01:02.37" resultid="6395" heatid="8003" lane="6" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00305" nation="POL" region="05" clubid="2281" name="UKS Nawa Skierniewice" shortname="Nawa Skierniewice">
          <CONTACT name="Marcin Sarna" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-11" firstname="Sebastian" gender="M" lastname="Krawczyk" nation="POL" license="S00305200017" athleteid="2282">
              <RESULTS>
                <RESULT eventid="1383" points="725" reactiontime="+89" swimtime="00:01:08.75" resultid="2283" heatid="7896" lane="5" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="767" reactiontime="+86" swimtime="00:00:30.86" resultid="2284" heatid="8048" lane="2" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01305" nation="POL" region="05" clubid="4151" name="UKS Piątka Konstantynów Ł." shortname="Piątka Konstantynów Ł.">
          <CONTACT name="Kotus Tomasz" phone="603820602" />
          <ATHLETES>
            <ATHLETE birthdate="1979-10-05" firstname="Marcin" gender="M" lastname="Grabarczyk" nation="POL" athleteid="4152">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="4153" heatid="7728" lane="2" entrytime="00:02:47.77" />
                <RESULT eventid="1156" status="WDR" swimtime="00:00:00.00" resultid="4154" entrytime="00:19:57.77" />
                <RESULT eventid="1222" points="472" reactiontime="+83" swimtime="00:03:00.41" resultid="4155" heatid="7789" lane="4" entrytime="00:03:27.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="150" swimtime="00:02:12.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="506" reactiontime="+78" swimtime="00:01:09.02" resultid="4156" heatid="7850" lane="2" entrytime="00:01:13.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="481" reactiontime="+85" swimtime="00:02:15.93" resultid="4157" heatid="7959" lane="3" entrytime="00:02:37.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                    <SPLIT distance="150" swimtime="00:01:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="4158" heatid="8808" lane="8" entrytime="00:06:17.00" />
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="4159" heatid="8015" lane="1" entrytime="00:02:57.77" />
                <RESULT eventid="1703" points="533" reactiontime="+87" swimtime="00:04:56.30" resultid="4160" heatid="9061" lane="5" entrytime="00:04:57.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:08.31" />
                    <SPLIT distance="150" swimtime="00:01:44.89" />
                    <SPLIT distance="200" swimtime="00:02:22.67" />
                    <SPLIT distance="250" swimtime="00:03:00.20" />
                    <SPLIT distance="300" swimtime="00:03:39.19" />
                    <SPLIT distance="350" swimtime="00:04:18.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="4161">
              <RESULTS>
                <RESULT eventid="1076" points="489" reactiontime="+89" swimtime="00:00:28.08" resultid="4162" heatid="7693" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1108" points="334" reactiontime="+92" swimtime="00:02:50.13" resultid="4163" heatid="7726" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:20.24" />
                    <SPLIT distance="150" swimtime="00:02:10.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="467" reactiontime="+88" swimtime="00:00:34.14" resultid="4164" heatid="7771" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1222" points="374" reactiontime="+90" swimtime="00:03:14.96" resultid="4165" heatid="7792" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                    <SPLIT distance="100" swimtime="00:01:30.90" />
                    <SPLIT distance="150" swimtime="00:02:24.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="359" reactiontime="+92" swimtime="00:01:26.25" resultid="4166" heatid="7890" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="WDR" swimtime="00:00:00.00" resultid="4167" entrytime="00:06:45.00" />
                <RESULT eventid="1623" points="262" reactiontime="+72" swimtime="00:03:02.08" resultid="4168" heatid="8015" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:01:24.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="405" reactiontime="+90" swimtime="00:00:37.56" resultid="4169" heatid="8038" lane="3" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-14" firstname="Jakub" gender="M" lastname="Gryczyński" nation="POL" athleteid="4170">
              <RESULTS>
                <RESULT eventid="1286" points="308" reactiontime="+86" swimtime="00:01:21.41" resultid="4171" heatid="7846" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="339" reactiontime="+93" swimtime="00:01:27.93" resultid="4172" heatid="7889" lane="6" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="377" reactiontime="+84" swimtime="00:00:38.49" resultid="4173" heatid="8039" lane="8" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-02" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="4174">
              <RESULTS>
                <RESULT eventid="1076" points="524" reactiontime="+96" swimtime="00:00:27.44" resultid="4175" heatid="7710" lane="8" entrytime="00:00:26.00" />
                <RESULT eventid="1254" points="440" reactiontime="+92" swimtime="00:01:04.43" resultid="4176" heatid="7817" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="365" reactiontime="+95" swimtime="00:00:31.98" resultid="4177" heatid="7917" lane="3" entrytime="00:00:31.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-11-12" firstname="Witold" gender="M" lastname="Pietrowski" nation="POL" athleteid="4178">
              <RESULTS>
                <RESULT eventid="1076" points="414" reactiontime="+86" swimtime="00:00:29.67" resultid="4179" heatid="7704" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1190" points="438" reactiontime="+73" swimtime="00:00:34.88" resultid="4180" heatid="7772" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1254" points="400" reactiontime="+80" swimtime="00:01:06.55" resultid="4181" heatid="7815" lane="7" entrytime="00:01:07.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="413" reactiontime="+77" swimtime="00:00:30.71" resultid="4182" heatid="7917" lane="5" entrytime="00:00:31.19" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="4183" heatid="7995" lane="5" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Rafał" gender="M" lastname="Trudnos" nation="POL" athleteid="4184">
              <RESULTS>
                <RESULT eventid="1076" points="502" reactiontime="+78" swimtime="00:00:27.84" resultid="4185" heatid="7707" lane="8" entrytime="00:00:27.13" />
                <RESULT eventid="1222" points="548" reactiontime="+75" swimtime="00:02:51.69" resultid="4186" heatid="7793" lane="7" entrytime="00:03:00.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:18.87" />
                    <SPLIT distance="150" swimtime="00:02:04.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="506" reactiontime="+76" swimtime="00:01:16.95" resultid="4187" heatid="7893" lane="4" entrytime="00:01:16.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="552" reactiontime="+75" swimtime="00:00:33.90" resultid="4188" heatid="8046" lane="2" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-06-12" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" athleteid="4189">
              <RESULTS>
                <RESULT eventid="1076" points="586" reactiontime="+82" swimtime="00:00:26.44" resultid="4190" heatid="7711" lane="1" entrytime="00:00:25.80" />
                <RESULT eventid="1254" points="550" reactiontime="+79" swimtime="00:00:59.82" resultid="4191" heatid="7822" lane="1" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="458" reactiontime="+80" swimtime="00:00:29.66" resultid="4192" heatid="7923" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1479" points="399" reactiontime="+86" swimtime="00:02:24.58" resultid="4193" heatid="7964" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="100" swimtime="00:01:05.38" />
                    <SPLIT distance="150" swimtime="00:01:44.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="454" reactiontime="+82" swimtime="00:01:08.45" resultid="4194" heatid="8000" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-08-19" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" athleteid="4195">
              <RESULTS>
                <RESULT eventid="1076" points="401" reactiontime="+81" swimtime="00:00:30.01" resultid="4196" heatid="7702" lane="1" entrytime="00:00:28.70" />
                <RESULT eventid="1286" points="324" reactiontime="+86" swimtime="00:01:20.00" resultid="4197" heatid="7845" lane="8" entrytime="00:01:23.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="4198" heatid="8040" lane="1" entrytime="00:00:37.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-04-28" firstname="Kornel" gender="M" lastname="Pintara" nation="POL" athleteid="4199">
              <RESULTS>
                <RESULT eventid="1254" points="495" reactiontime="+82" swimtime="00:01:05.00" resultid="4200" heatid="7819" lane="4" entrytime="00:01:02.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="460" reactiontime="+85" swimtime="00:01:16.47" resultid="4201" heatid="7849" lane="7" entrytime="00:01:14.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="422" reactiontime="+87" swimtime="00:00:34.20" resultid="4202" heatid="7917" lane="6" entrytime="00:00:31.28" />
                <RESULT eventid="1479" points="347" reactiontime="+93" swimtime="00:02:38.59" resultid="4203" heatid="7962" lane="8" entrytime="00:02:27.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="150" swimtime="00:01:55.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="4204" heatid="8017" lane="3" entrytime="00:02:40.00" />
                <RESULT eventid="1655" points="392" reactiontime="+86" swimtime="00:00:39.42" resultid="4205" heatid="8039" lane="4" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="4206">
              <RESULTS>
                <RESULT eventid="1108" points="464" reactiontime="+80" swimtime="00:02:44.43" resultid="4207" heatid="7727" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                    <SPLIT distance="150" swimtime="00:02:05.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="523" swimtime="00:20:53.83" resultid="4208" heatid="8720" lane="1" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:13.62" />
                    <SPLIT distance="200" swimtime="00:02:31.96" />
                    <SPLIT distance="300" swimtime="00:03:55.00" />
                    <SPLIT distance="400" swimtime="00:05:20.01" />
                    <SPLIT distance="500" swimtime="00:06:44.98" />
                    <SPLIT distance="600" swimtime="00:08:10.27" />
                    <SPLIT distance="700" swimtime="00:09:35.10" />
                    <SPLIT distance="800" swimtime="00:11:00.20" />
                    <SPLIT distance="900" swimtime="00:12:24.57" />
                    <SPLIT distance="1000" swimtime="00:13:49.06" />
                    <SPLIT distance="1100" swimtime="00:15:15.17" />
                    <SPLIT distance="1200" swimtime="00:16:40.45" />
                    <SPLIT distance="1300" swimtime="00:18:05.54" />
                    <SPLIT distance="1400" swimtime="00:19:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="623" reactiontime="+77" swimtime="00:00:30.04" resultid="4209" heatid="7913" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="4210" heatid="7998" lane="3" entrytime="00:01:15.00" />
                <RESULT eventid="1703" points="439" reactiontime="+70" swimtime="00:05:18.68" resultid="4211" heatid="9064" lane="6" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:47.25" />
                    <SPLIT distance="200" swimtime="00:02:27.78" />
                    <SPLIT distance="250" swimtime="00:03:09.74" />
                    <SPLIT distance="300" swimtime="00:03:52.13" />
                    <SPLIT distance="350" swimtime="00:04:36.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-04" firstname="Jakub" gender="M" lastname="Sidorowicz" nation="POL" athleteid="4212">
              <RESULTS>
                <RESULT eventid="1108" points="186" reactiontime="+85" swimtime="00:03:26.78" resultid="4213" heatid="7721" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:01:33.50" />
                    <SPLIT distance="150" swimtime="00:02:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="267" reactiontime="+76" swimtime="00:00:41.11" resultid="4214" heatid="7766" lane="8" entrytime="00:00:48.00" />
                <RESULT eventid="1286" points="235" reactiontime="+92" swimtime="00:01:29.08" resultid="4215" heatid="7839" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="254" reactiontime="+101" swimtime="00:01:36.79" resultid="4216" heatid="7882" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="4217" heatid="7935" lane="1" entrytime="00:01:40.00" />
                <RESULT eventid="1655" points="291" reactiontime="+80" swimtime="00:00:41.95" resultid="4218" heatid="8032" lane="8" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-14" firstname="Tomasz" gender="M" lastname="Kotus" nation="POL" athleteid="4226">
              <RESULTS>
                <RESULT eventid="1156" points="521" swimtime="00:20:52.67" resultid="4227" heatid="8719" lane="6" entrytime="00:21:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:12.81" />
                    <SPLIT distance="200" swimtime="00:02:31.16" />
                    <SPLIT distance="400" swimtime="00:05:12.42" />
                    <SPLIT distance="500" swimtime="00:06:36.05" />
                    <SPLIT distance="600" swimtime="00:08:01.70" />
                    <SPLIT distance="700" swimtime="00:09:29.38" />
                    <SPLIT distance="800" swimtime="00:10:54.78" />
                    <SPLIT distance="900" swimtime="00:12:21.14" />
                    <SPLIT distance="1000" swimtime="00:13:48.39" />
                    <SPLIT distance="1100" swimtime="00:15:12.63" />
                    <SPLIT distance="1200" swimtime="00:16:41.79" />
                    <SPLIT distance="1300" swimtime="00:18:06.55" />
                    <SPLIT distance="1400" swimtime="00:19:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="408" reactiontime="+85" swimtime="00:02:47.15" resultid="4228" heatid="7863" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:58.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="513" reactiontime="+84" swimtime="00:00:28.56" resultid="4229" heatid="7922" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1543" points="476" reactiontime="+82" swimtime="00:05:41.82" resultid="4230" heatid="8808" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:13.10" />
                    <SPLIT distance="150" swimtime="00:01:59.69" />
                    <SPLIT distance="200" swimtime="00:02:46.50" />
                    <SPLIT distance="250" swimtime="00:03:37.55" />
                    <SPLIT distance="300" swimtime="00:04:27.62" />
                    <SPLIT distance="350" swimtime="00:05:06.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="463" reactiontime="+89" swimtime="00:01:08.01" resultid="4231" heatid="8000" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="354" reactiontime="+75" swimtime="00:02:44.89" resultid="4232" heatid="8015" lane="7" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:17.14" />
                    <SPLIT distance="150" swimtime="00:02:01.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="WDR" swimtime="00:00:00.00" resultid="4233" heatid="8036" lane="5" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Piatka Konstantynów B" number="1">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+90" swimtime="00:02:07.56" resultid="4245" heatid="7872" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:41.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4161" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="4184" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4206" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="4189" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Piatka Konstantynów Ł. B" number="1">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+78" swimtime="00:01:48.79" resultid="4243" heatid="7973" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                    <SPLIT distance="100" swimtime="00:00:55.28" />
                    <SPLIT distance="150" swimtime="00:01:22.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4184" number="1" />
                    <RELAYPOSITION athleteid="4174" number="2" />
                    <RELAYPOSITION athleteid="4152" number="3" />
                    <RELAYPOSITION athleteid="4189" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Piatka Konstantynów B" number="2">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+71" swimtime="00:02:12.69" resultid="4247" heatid="7871" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:45.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4152" number="1" />
                    <RELAYPOSITION athleteid="4195" number="2" />
                    <RELAYPOSITION athleteid="4199" number="3" />
                    <RELAYPOSITION athleteid="4174" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Piatka Konstantynów Ł. B" number="2">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+81" swimtime="00:01:51.85" resultid="4244" heatid="7973" lane="3" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                    <SPLIT distance="100" swimtime="00:00:56.80" />
                    <SPLIT distance="150" swimtime="00:01:23.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4178" number="1" />
                    <RELAYPOSITION athleteid="4206" number="2" />
                    <RELAYPOSITION athleteid="4226" number="3" />
                    <RELAYPOSITION athleteid="4161" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Piatka Konstantynów Ł. B" number="3">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+81" swimtime="00:02:03.58" resultid="4246" heatid="7973" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="100" swimtime="00:01:00.11" />
                    <SPLIT distance="150" swimtime="00:01:31.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4195" number="1" />
                    <RELAYPOSITION athleteid="4199" number="2" />
                    <RELAYPOSITION athleteid="4170" number="3" />
                    <RELAYPOSITION athleteid="4212" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Piątka Konstantynów B" number="3">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+73" swimtime="00:02:18.42" resultid="4248" heatid="7871" lane="1" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                    <SPLIT distance="100" swimtime="00:01:19.19" />
                    <SPLIT distance="150" swimtime="00:01:50.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4212" number="1" />
                    <RELAYPOSITION athleteid="4170" number="2" />
                    <RELAYPOSITION athleteid="4178" number="3" />
                    <RELAYPOSITION athleteid="4226" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00706" nation="POL" region="06" clubid="1861" name="UKS SP 8 Chrzanów" shortname="UKS SP 8 Chrzanów             ">
          <CONTACT city="Chrzanów" email="abalp@poczta.onet.pl" name="Zabrzański Alfred" phone="692076808" state="MAŁOP" street="Niepodległości 7/46" zip="32-500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="1862">
              <RESULTS>
                <RESULT eventid="1076" points="645" reactiontime="+84" swimtime="00:00:30.17" resultid="1863" heatid="7697" lane="1" entrytime="00:00:30.20" entrycourse="SCM" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="1864" heatid="8721" lane="2" entrytime="00:24:15.00" entrycourse="SCM" />
                <RESULT eventid="1254" points="618" reactiontime="+81" swimtime="00:01:08.12" resultid="1865" heatid="7814" lane="6" entrytime="00:01:09.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="570" reactiontime="+84" swimtime="00:01:23.41" resultid="1866" heatid="7844" lane="4" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="1867" heatid="7959" lane="6" entrytime="00:02:39.00" entrycourse="SCM" />
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="1868" heatid="9066" lane="1" entrytime="00:05:52.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TROBO" nation="POL" region="15" clubid="2402" name="UKS Trójka Oborniki" shortname="Trójka Oborniki">
          <CONTACT city="Oborniki" email="janwol@poczta.onet.pl" name="Wolniewicz" phone="791064667" state="WIE" street="Piłsudskiego 49/42" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="2403">
              <RESULTS>
                <RESULT eventid="1076" points="487" reactiontime="+108" swimtime="00:00:35.80" resultid="2404" heatid="7689" lane="2" entrytime="00:00:35.08" />
                <RESULT eventid="1156" points="430" swimtime="00:29:08.91" resultid="2405" heatid="8723" lane="6" entrytime="00:27:27.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.78" />
                    <SPLIT distance="100" swimtime="00:01:40.57" />
                    <SPLIT distance="200" swimtime="00:03:31.71" />
                    <SPLIT distance="300" swimtime="00:05:25.20" />
                    <SPLIT distance="400" swimtime="00:07:20.66" />
                    <SPLIT distance="500" swimtime="00:09:16.83" />
                    <SPLIT distance="600" swimtime="00:11:12.93" />
                    <SPLIT distance="700" swimtime="00:13:10.47" />
                    <SPLIT distance="800" swimtime="00:15:09.37" />
                    <SPLIT distance="900" swimtime="00:17:08.81" />
                    <SPLIT distance="1000" swimtime="00:19:08.71" />
                    <SPLIT distance="1100" swimtime="00:21:08.33" />
                    <SPLIT distance="1200" swimtime="00:23:09.78" />
                    <SPLIT distance="1300" swimtime="00:25:11.20" />
                    <SPLIT distance="1400" swimtime="00:27:12.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="476" reactiontime="+107" swimtime="00:01:21.17" resultid="2406" heatid="7808" lane="4" entrytime="00:01:21.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="407" reactiontime="+116" swimtime="00:03:16.86" resultid="2407" heatid="7954" lane="7" entrytime="00:03:18.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                    <SPLIT distance="100" swimtime="00:01:32.79" />
                    <SPLIT distance="150" swimtime="00:02:25.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="334" reactiontime="+110" swimtime="00:07:22.63" resultid="2408" heatid="9069" lane="1" entrytime="00:07:20.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.81" />
                    <SPLIT distance="100" swimtime="00:01:41.07" />
                    <SPLIT distance="150" swimtime="00:02:37.05" />
                    <SPLIT distance="200" swimtime="00:03:33.12" />
                    <SPLIT distance="250" swimtime="00:04:30.16" />
                    <SPLIT distance="300" swimtime="00:05:28.37" />
                    <SPLIT distance="350" swimtime="00:06:25.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02914" nation="POL" region="14" clubid="3004" name="UKS Victoria Józefów" shortname="Victoria Józefów">
          <CONTACT email="ali90@o2.pl" name="KOWALCZYK ALICJA" />
          <ATHLETES>
            <ATHLETE birthdate="1966-03-01" firstname="Jan" gender="M" lastname="Kośmider" nation="POL" athleteid="3013">
              <RESULTS>
                <RESULT eventid="1076" points="609" reactiontime="+83" swimtime="00:00:28.52" resultid="3014" heatid="7700" lane="8" entrytime="00:00:29.51" />
                <RESULT eventid="1156" points="449" swimtime="00:21:31.05" resultid="3015" heatid="8718" lane="3" entrytime="00:20:50.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="200" swimtime="00:02:41.41" />
                    <SPLIT distance="300" swimtime="00:04:04.70" />
                    <SPLIT distance="400" swimtime="00:05:29.55" />
                    <SPLIT distance="500" swimtime="00:06:55.31" />
                    <SPLIT distance="600" swimtime="00:08:22.07" />
                    <SPLIT distance="700" swimtime="00:09:49.59" />
                    <SPLIT distance="800" swimtime="00:11:17.38" />
                    <SPLIT distance="900" swimtime="00:12:45.93" />
                    <SPLIT distance="1000" swimtime="00:14:13.70" />
                    <SPLIT distance="1100" swimtime="00:15:40.38" />
                    <SPLIT distance="1200" swimtime="00:17:08.31" />
                    <SPLIT distance="1300" swimtime="00:18:36.35" />
                    <SPLIT distance="1400" swimtime="00:20:04.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="601" reactiontime="+82" swimtime="00:02:56.80" resultid="3016" heatid="7793" lane="1" entrytime="00:03:02.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:25.31" />
                    <SPLIT distance="150" swimtime="00:02:11.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="637" reactiontime="+96" swimtime="00:01:18.12" resultid="3017" heatid="7890" lane="3" entrytime="00:01:24.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="647" reactiontime="+91" swimtime="00:05:51.57" resultid="3018" heatid="8807" lane="7" entrytime="00:05:50.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:28.88" />
                    <SPLIT distance="150" swimtime="00:02:15.36" />
                    <SPLIT distance="200" swimtime="00:03:00.22" />
                    <SPLIT distance="250" swimtime="00:03:47.89" />
                    <SPLIT distance="300" swimtime="00:04:35.24" />
                    <SPLIT distance="350" swimtime="00:05:15.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="687" reactiontime="+79" swimtime="00:00:34.76" resultid="3019" heatid="8042" lane="7" entrytime="00:00:36.50" />
                <RESULT eventid="1703" points="495" reactiontime="+83" swimtime="00:05:10.74" resultid="3020" heatid="9061" lane="4" entrytime="00:04:55.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:13.44" />
                    <SPLIT distance="150" swimtime="00:01:52.97" />
                    <SPLIT distance="200" swimtime="00:02:33.36" />
                    <SPLIT distance="250" swimtime="00:03:13.50" />
                    <SPLIT distance="300" swimtime="00:03:53.17" />
                    <SPLIT distance="350" swimtime="00:04:32.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03311" nation="POL" region="11" clubid="5830" name="UKS Wodnik 29 Katowice" shortname="Wodnik 29 Katowice">
          <CONTACT email="skoczyt@gmail.com" name="Skoczylas Tomasz" phone="662297707" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-10" firstname="Sandra" gender="F" lastname="Pietrzak" nation="POL" athleteid="5838">
              <RESULTS>
                <RESULT eventid="1173" status="DNS" swimtime="00:00:00.00" resultid="5839" heatid="7760" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1238" points="659" reactiontime="+77" swimtime="00:01:06.49" resultid="5840" heatid="7805" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="556" reactiontime="+82" swimtime="00:00:34.80" resultid="5841" heatid="7903" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1431" points="555" reactiontime="+80" swimtime="00:01:19.33" resultid="5842" heatid="7931" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" status="WDR" swimtime="00:00:00.00" resultid="5843" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-19" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="5864">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5865" heatid="7694" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="1254" points="550" reactiontime="+94" swimtime="00:01:13.03" resultid="5866" heatid="7811" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="411" reactiontime="+95" swimtime="00:03:34.77" resultid="5867" heatid="7862" lane="8" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:39.02" />
                    <SPLIT distance="150" swimtime="00:02:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="668" reactiontime="+94" swimtime="00:00:34.25" resultid="5868" heatid="7914" lane="3" entrytime="00:00:33.99" />
                <RESULT eventid="1479" points="451" reactiontime="+99" swimtime="00:02:59.77" resultid="5869" heatid="7956" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:23.11" />
                    <SPLIT distance="150" swimtime="00:02:13.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="5870" heatid="7994" lane="8" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="5871">
              <RESULTS>
                <RESULT eventid="1059" points="672" reactiontime="+81" swimtime="00:00:29.84" resultid="5872" heatid="7682" lane="3" entrytime="00:00:29.90" />
                <RESULT eventid="1140" points="549" reactiontime="+95" swimtime="00:11:45.91" resultid="5873" heatid="8712" lane="7" entrytime="00:10:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:18.35" />
                    <SPLIT distance="150" swimtime="00:02:01.67" />
                    <SPLIT distance="200" swimtime="00:02:45.92" />
                    <SPLIT distance="250" swimtime="00:03:31.04" />
                    <SPLIT distance="300" swimtime="00:04:16.53" />
                    <SPLIT distance="350" swimtime="00:05:01.52" />
                    <SPLIT distance="400" swimtime="00:05:46.83" />
                    <SPLIT distance="450" swimtime="00:06:32.40" />
                    <SPLIT distance="500" swimtime="00:07:18.01" />
                    <SPLIT distance="550" swimtime="00:08:03.46" />
                    <SPLIT distance="600" swimtime="00:08:48.65" />
                    <SPLIT distance="650" swimtime="00:09:33.77" />
                    <SPLIT distance="700" swimtime="00:10:18.35" />
                    <SPLIT distance="750" swimtime="00:10:59.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="644" reactiontime="+84" swimtime="00:01:06.53" resultid="5874" heatid="7804" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="734" reactiontime="+87" swimtime="00:00:32.21" resultid="5875" heatid="7905" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1463" points="575" reactiontime="+90" swimtime="00:02:31.41" resultid="5876" heatid="7950" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:11.46" />
                    <SPLIT distance="150" swimtime="00:01:51.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="573" reactiontime="+88" swimtime="00:01:16.78" resultid="5877" heatid="7991" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" status="WDR" swimtime="00:00:00.00" resultid="5878" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-08-07" firstname="Marzena" gender="F" lastname="Fligier" nation="POL" athleteid="5879">
              <RESULTS>
                <RESULT eventid="1206" points="334" reactiontime="+123" swimtime="00:03:59.38" resultid="5880" heatid="7780" lane="3" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.57" />
                    <SPLIT distance="100" swimtime="00:01:52.87" />
                    <SPLIT distance="150" swimtime="00:02:56.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="311" reactiontime="+141" swimtime="00:01:51.69" resultid="5881" heatid="7876" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="5882">
              <RESULTS>
                <RESULT eventid="1076" points="670" reactiontime="+85" swimtime="00:00:27.62" resultid="5883" heatid="7701" lane="4" entrytime="00:00:28.91" />
                <RESULT eventid="1156" points="560" swimtime="00:19:59.15" resultid="5884" heatid="8719" lane="8" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="200" swimtime="00:02:33.02" />
                    <SPLIT distance="300" swimtime="00:03:52.46" />
                    <SPLIT distance="400" swimtime="00:05:11.78" />
                    <SPLIT distance="500" swimtime="00:06:32.35" />
                    <SPLIT distance="600" swimtime="00:07:52.81" />
                    <SPLIT distance="700" swimtime="00:09:12.78" />
                    <SPLIT distance="800" swimtime="00:10:32.66" />
                    <SPLIT distance="900" swimtime="00:11:53.17" />
                    <SPLIT distance="1000" swimtime="00:13:14.99" />
                    <SPLIT distance="1100" swimtime="00:14:36.20" />
                    <SPLIT distance="1200" swimtime="00:15:58.04" />
                    <SPLIT distance="1300" swimtime="00:17:19.73" />
                    <SPLIT distance="1400" swimtime="00:18:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="606" reactiontime="+97" swimtime="00:00:33.85" resultid="5885" heatid="7771" lane="3" entrytime="00:00:35.50" />
                <RESULT eventid="1254" points="667" reactiontime="+82" swimtime="00:01:00.56" resultid="5886" heatid="7820" lane="3" entrytime="00:01:01.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="603" reactiontime="+86" swimtime="00:01:13.54" resultid="5887" heatid="7939" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="564" reactiontime="+101" swimtime="00:02:18.83" resultid="5888" heatid="7963" lane="8" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="613" reactiontime="+89" swimtime="00:02:40.40" resultid="5889" heatid="8017" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:18.63" />
                    <SPLIT distance="150" swimtime="00:01:59.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="573" reactiontime="+99" swimtime="00:04:55.96" resultid="5890" heatid="9062" lane="3" entrytime="00:05:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:10.22" />
                    <SPLIT distance="150" swimtime="00:01:48.00" />
                    <SPLIT distance="200" swimtime="00:02:26.89" />
                    <SPLIT distance="250" swimtime="00:03:05.32" />
                    <SPLIT distance="300" swimtime="00:03:43.56" />
                    <SPLIT distance="350" swimtime="00:04:20.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="5891">
              <RESULTS>
                <RESULT eventid="1222" points="573" reactiontime="+75" swimtime="00:03:06.27" resultid="5892" heatid="7792" lane="6" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                    <SPLIT distance="100" swimtime="00:01:28.11" />
                    <SPLIT distance="150" swimtime="00:02:16.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="651" reactiontime="+80" swimtime="00:01:15.53" resultid="5893" heatid="7847" lane="7" entrytime="00:01:17.00" />
                <RESULT eventid="1383" points="602" reactiontime="+81" swimtime="00:01:22.33" resultid="5894" heatid="7891" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="5895" heatid="7957" lane="5" entrytime="00:02:45.00" />
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)  (Czas: 11:37)" eventid="1655" reactiontime="+61" status="DSQ" swimtime="00:00:35.43" resultid="5896" heatid="8043" lane="1" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-16" firstname="Elżbieta" gender="F" lastname="Fira" nation="POL" athleteid="5897">
              <RESULTS>
                <RESULT eventid="1059" points="410" reactiontime="+82" swimtime="00:00:36.56" resultid="5898" heatid="7675" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1238" points="359" reactiontime="+84" swimtime="00:01:21.31" resultid="5899" heatid="7800" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="376" reactiontime="+84" swimtime="00:01:34.02" resultid="5900" heatid="7829" lane="5" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="410" reactiontime="+85" swimtime="00:00:39.72" resultid="5901" heatid="7899" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1463" points="303" reactiontime="+84" swimtime="00:03:10.57" resultid="5902" heatid="7946" lane="3" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                    <SPLIT distance="100" swimtime="00:01:32.73" />
                    <SPLIT distance="150" swimtime="00:02:22.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="352" reactiontime="+96" swimtime="00:00:47.98" resultid="5903" heatid="8023" lane="6" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-05-18" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="5904">
              <RESULTS>
                <RESULT eventid="1059" points="369" reactiontime="+131" swimtime="00:01:07.75" resultid="5905" heatid="7671" lane="5" entrytime="00:01:05.00" />
                <RESULT eventid="1140" points="421" swimtime="00:24:45.59" resultid="5906" heatid="8716" lane="6" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.20" />
                    <SPLIT distance="100" swimtime="00:02:40.14" />
                    <SPLIT distance="200" swimtime="00:05:41.80" />
                    <SPLIT distance="300" swimtime="00:08:47.92" />
                    <SPLIT distance="400" swimtime="00:11:59.47" />
                    <SPLIT distance="500" swimtime="00:15:09.94" />
                    <SPLIT distance="600" swimtime="00:18:29.90" />
                    <SPLIT distance="700" swimtime="00:21:39.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="394" reactiontime="+88" swimtime="00:01:13.02" resultid="5907" heatid="7754" lane="7" entrytime="00:01:10.00" />
                <RESULT eventid="1238" points="353" reactiontime="+127" swimtime="00:02:42.93" resultid="5908" heatid="7796" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" status="DNS" swimtime="00:00:00.00" resultid="5909" heatid="7926" lane="2" entrytime="00:02:38.00" />
                <RESULT eventid="1687" points="320" reactiontime="+112" swimtime="00:11:57.07" resultid="5910" heatid="9053" lane="5" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.71" />
                    <SPLIT distance="100" swimtime="00:02:46.27" />
                    <SPLIT distance="150" swimtime="00:04:19.80" />
                    <SPLIT distance="200" swimtime="00:05:52.89" />
                    <SPLIT distance="250" swimtime="00:07:26.78" />
                    <SPLIT distance="300" swimtime="00:08:59.91" />
                    <SPLIT distance="350" swimtime="00:10:32.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-15" firstname="Andrzej" gender="M" lastname="Porszke" nation="POL" athleteid="5911">
              <RESULTS>
                <RESULT eventid="1222" points="306" reactiontime="+112" swimtime="00:03:31.28" resultid="5912" heatid="7789" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.06" />
                    <SPLIT distance="100" swimtime="00:01:38.96" />
                    <SPLIT distance="150" swimtime="00:02:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="333" reactiontime="+95" swimtime="00:01:32.32" resultid="5913" heatid="7887" lane="2" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="354" reactiontime="+96" swimtime="00:00:40.80" resultid="5914" heatid="8037" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-08" firstname="Paweł" gender="M" lastname="Dygdoń" nation="POL" athleteid="5915">
              <RESULTS>
                <RESULT eventid="1108" points="481" reactiontime="+80" swimtime="00:02:42.40" resultid="5916" heatid="7728" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="150" swimtime="00:02:02.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="473" swimtime="00:21:36.55" resultid="5917" heatid="8718" lane="6" entrytime="00:20:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:13.40" />
                    <SPLIT distance="200" swimtime="00:02:35.09" />
                    <SPLIT distance="300" swimtime="00:04:00.81" />
                    <SPLIT distance="400" swimtime="00:05:27.48" />
                    <SPLIT distance="500" swimtime="00:06:54.72" />
                    <SPLIT distance="600" swimtime="00:08:22.75" />
                    <SPLIT distance="700" swimtime="00:09:51.06" />
                    <SPLIT distance="800" swimtime="00:11:19.24" />
                    <SPLIT distance="900" swimtime="00:12:47.31" />
                    <SPLIT distance="1000" swimtime="00:14:15.70" />
                    <SPLIT distance="1100" swimtime="00:15:44.24" />
                    <SPLIT distance="1200" swimtime="00:17:12.93" />
                    <SPLIT distance="1300" swimtime="00:18:41.43" />
                    <SPLIT distance="1400" swimtime="00:20:10.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="506" reactiontime="+74" swimtime="00:01:14.10" resultid="5918" heatid="7848" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="5919" heatid="7864" lane="7" entrytime="00:02:50.00" />
                <RESULT eventid="1447" points="474" reactiontime="+82" swimtime="00:01:15.80" resultid="5920" heatid="7937" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="465" reactiontime="+86" swimtime="00:05:52.13" resultid="5921" heatid="8809" lane="4" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="150" swimtime="00:01:59.11" />
                    <SPLIT distance="200" swimtime="00:02:44.70" />
                    <SPLIT distance="250" swimtime="00:03:35.55" />
                    <SPLIT distance="300" swimtime="00:04:27.06" />
                    <SPLIT distance="350" swimtime="00:05:10.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="492" reactiontime="+83" swimtime="00:01:12.02" resultid="5922" heatid="7997" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="471" reactiontime="+92" swimtime="00:02:46.98" resultid="5923" heatid="8017" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                    <SPLIT distance="150" swimtime="00:02:03.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-26" firstname="Piotr" gender="M" lastname="Klepacki" nation="POL" athleteid="5924">
              <RESULTS>
                <RESULT eventid="1222" points="165" reactiontime="+85" swimtime="00:04:19.40" resultid="5925" heatid="7786" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.27" />
                    <SPLIT distance="100" swimtime="00:01:57.25" />
                    <SPLIT distance="150" swimtime="00:03:07.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="200" reactiontime="+69" swimtime="00:01:49.44" resultid="5926" heatid="7883" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-12-22" firstname="Sylwia" gender="F" lastname="Kornaś" nation="POL" athleteid="5927">
              <RESULTS>
                <RESULT eventid="1059" points="388" swimtime="00:00:35.83" resultid="5928" heatid="7677" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1173" points="311" reactiontime="+79" swimtime="00:00:44.79" resultid="5929" heatid="7757" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1270" points="300" reactiontime="+87" swimtime="00:01:37.16" resultid="5930" heatid="7829" lane="4" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="343" reactiontime="+91" swimtime="00:01:43.81" resultid="5931" heatid="7877" lane="7" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="311" reactiontime="+77" swimtime="00:01:38.12" resultid="5932" heatid="7927" lane="6" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="312" reactiontime="+78" swimtime="00:03:28.79" resultid="5933" heatid="8006" lane="8" entrytime="00:03:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.22" />
                    <SPLIT distance="100" swimtime="00:01:41.85" />
                    <SPLIT distance="150" swimtime="00:02:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="284" reactiontime="+86" swimtime="00:00:48.26" resultid="5934" heatid="8024" lane="5" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-03-15" firstname="Jolanta" gender="F" lastname="Stefanek" nation="POL" athleteid="5935">
              <RESULTS>
                <RESULT eventid="1206" points="544" reactiontime="+70" swimtime="00:03:37.37" resultid="5936" heatid="7782" lane="1" entrytime="00:03:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.50" />
                    <SPLIT distance="100" swimtime="00:01:41.27" />
                    <SPLIT distance="150" swimtime="00:02:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="356" reactiontime="+86" swimtime="00:01:42.37" resultid="5937" heatid="7830" lane="1" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="516" reactiontime="+76" swimtime="00:01:39.99" resultid="5938" heatid="7878" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="235" reactiontime="+81" swimtime="00:00:50.43" resultid="5939" heatid="7900" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1639" points="527" reactiontime="+88" swimtime="00:00:45.37" resultid="5940" heatid="8026" lane="2" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-06-09" firstname="Edyta" gender="F" lastname="Mróz" nation="POL" athleteid="5941">
              <RESULTS>
                <RESULT eventid="1431" points="582" reactiontime="+92" swimtime="00:01:19.67" resultid="5942" heatid="7930" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="489" reactiontime="+89" swimtime="00:02:39.83" resultid="5943" heatid="7949" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                    <SPLIT distance="150" swimtime="00:01:58.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="546" reactiontime="+89" swimtime="00:02:53.16" resultid="5944" heatid="8008" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:23.93" />
                    <SPLIT distance="150" swimtime="00:02:09.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="510" reactiontime="+91" swimtime="00:05:42.28" resultid="5945" heatid="9049" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="100" swimtime="00:01:19.70" />
                    <SPLIT distance="150" swimtime="00:02:03.56" />
                    <SPLIT distance="200" swimtime="00:02:48.16" />
                    <SPLIT distance="250" swimtime="00:03:32.13" />
                    <SPLIT distance="300" swimtime="00:04:16.23" />
                    <SPLIT distance="350" swimtime="00:05:00.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="5946">
              <RESULTS>
                <RESULT eventid="1076" points="734" reactiontime="+93" swimtime="00:00:28.90" resultid="5947" heatid="7701" lane="5" entrytime="00:00:28.94" />
                <RESULT eventid="1254" points="637" reactiontime="+91" swimtime="00:01:07.42" resultid="5948" heatid="7815" lane="2" entrytime="00:01:07.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="726" reactiontime="+94" swimtime="00:00:31.73" resultid="5949" heatid="7917" lane="8" entrytime="00:00:31.40" />
                <RESULT eventid="1591" points="708" reactiontime="+98" swimtime="00:01:12.67" resultid="5950" heatid="7998" lane="8" entrytime="00:01:16.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-05" firstname="Marcin" gender="M" lastname="Szczypiński" nation="POL" athleteid="5951">
              <RESULTS>
                <RESULT eventid="1076" points="863" reactiontime="+73" swimtime="00:00:23.99" resultid="5952" heatid="7712" lane="1" entrytime="00:00:25.00" />
                <RESULT eventid="1156" points="791" reactiontime="+87" swimtime="00:17:27.30" resultid="5953" heatid="8717" lane="4" entrytime="00:17:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:05.56" />
                    <SPLIT distance="150" swimtime="00:01:40.36" />
                    <SPLIT distance="200" swimtime="00:02:15.69" />
                    <SPLIT distance="250" swimtime="00:02:50.69" />
                    <SPLIT distance="300" swimtime="00:03:26.11" />
                    <SPLIT distance="350" swimtime="00:04:01.56" />
                    <SPLIT distance="400" swimtime="00:04:36.88" />
                    <SPLIT distance="450" swimtime="00:05:12.12" />
                    <SPLIT distance="500" swimtime="00:05:47.35" />
                    <SPLIT distance="550" swimtime="00:06:22.62" />
                    <SPLIT distance="600" swimtime="00:06:58.10" />
                    <SPLIT distance="650" swimtime="00:07:32.92" />
                    <SPLIT distance="700" swimtime="00:08:07.85" />
                    <SPLIT distance="750" swimtime="00:08:42.45" />
                    <SPLIT distance="800" swimtime="00:09:17.38" />
                    <SPLIT distance="850" swimtime="00:09:52.37" />
                    <SPLIT distance="900" swimtime="00:10:27.30" />
                    <SPLIT distance="950" swimtime="00:11:02.57" />
                    <SPLIT distance="1000" swimtime="00:11:37.76" />
                    <SPLIT distance="1050" swimtime="00:12:13.28" />
                    <SPLIT distance="1100" swimtime="00:12:48.64" />
                    <SPLIT distance="1150" swimtime="00:13:23.70" />
                    <SPLIT distance="1200" swimtime="00:13:59.08" />
                    <SPLIT distance="1250" swimtime="00:14:34.28" />
                    <SPLIT distance="1300" swimtime="00:15:09.72" />
                    <SPLIT distance="1350" swimtime="00:15:44.80" />
                    <SPLIT distance="1400" swimtime="00:16:20.10" />
                    <SPLIT distance="1450" swimtime="00:16:54.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="695" reactiontime="+67" swimtime="00:00:28.28" resultid="5954" heatid="7777" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="1254" points="797" reactiontime="+76" swimtime="00:00:52.38" resultid="5955" heatid="7825" lane="6" entrytime="00:00:54.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="762" reactiontime="+75" swimtime="00:00:25.94" resultid="5956" heatid="7925" lane="1" entrytime="00:00:26.80" />
                <RESULT eventid="1479" points="812" reactiontime="+77" swimtime="00:02:00.62" resultid="5957" heatid="7967" lane="3" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                    <SPLIT distance="100" swimtime="00:00:57.47" />
                    <SPLIT distance="150" swimtime="00:01:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="822" reactiontime="+78" swimtime="00:00:57.57" resultid="5958" heatid="8003" lane="7" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="819" reactiontime="+82" swimtime="00:04:21.22" resultid="5959" heatid="9059" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:04.10" />
                    <SPLIT distance="150" swimtime="00:01:37.51" />
                    <SPLIT distance="200" swimtime="00:02:11.23" />
                    <SPLIT distance="250" swimtime="00:02:44.71" />
                    <SPLIT distance="300" swimtime="00:03:18.36" />
                    <SPLIT distance="350" swimtime="00:03:50.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-16" firstname="Michał" gender="M" lastname="Spławiński" nation="POL" athleteid="5960">
              <RESULTS>
                <RESULT eventid="1076" points="693" reactiontime="+69" swimtime="00:00:25.00" resultid="5961" heatid="7712" lane="2" entrytime="00:00:24.99" />
                <RESULT eventid="1108" points="524" reactiontime="+82" swimtime="00:02:26.52" resultid="5962" heatid="7729" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="150" swimtime="00:01:52.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="679" reactiontime="+67" swimtime="00:00:30.15" resultid="5963" heatid="7775" lane="6" entrytime="00:00:30.90" />
                <RESULT eventid="1286" points="682" reactiontime="+76" swimtime="00:01:02.46" resultid="5964" heatid="7856" lane="7" entrytime="00:01:02.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="751" reactiontime="+82" swimtime="00:01:07.48" resultid="5965" heatid="7895" lane="7" entrytime="00:01:11.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="648" reactiontime="+77" swimtime="00:00:26.42" resultid="5966" heatid="7925" lane="8" entrytime="00:00:26.88" />
                <RESULT eventid="1655" points="747" reactiontime="+75" swimtime="00:00:30.65" resultid="5967" heatid="8048" lane="1" entrytime="00:00:30.78" />
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="5968" entrytime="00:05:00.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-11-14" firstname="Aleksander" gender="M" lastname="Aleksandrowicz" nation="POL" athleteid="5969">
              <RESULTS>
                <RESULT eventid="1190" points="368" reactiontime="+77" swimtime="00:00:55.66" resultid="5970" heatid="7764" lane="3" entrytime="00:00:54.70" />
                <RESULT eventid="1222" points="304" reactiontime="+109" swimtime="00:04:50.62" resultid="5971" heatid="7785" lane="5" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.16" />
                    <SPLIT distance="100" swimtime="00:02:18.69" />
                    <SPLIT distance="150" swimtime="00:03:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="271" reactiontime="+112" swimtime="00:02:13.92" resultid="5972" heatid="7881" lane="4" entrytime="00:02:13.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="293" reactiontime="+98" swimtime="00:00:59.02" resultid="5973" heatid="8030" lane="6" entrytime="00:00:59.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-08-30" firstname="Aleksandra" gender="F" lastname="Kącki" nation="POL" athleteid="5977">
              <RESULTS>
                <RESULT eventid="1059" points="288" reactiontime="+129" swimtime="00:00:41.12" resultid="5978" heatid="7674" lane="5" entrytime="00:00:41.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-07-07" firstname="Tomasz" gender="M" lastname="Szabelka" nation="POL" athleteid="5979">
              <RESULTS>
                <RESULT eventid="1076" points="380" reactiontime="+110" swimtime="00:00:32.72" resultid="5980" heatid="7691" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1254" points="311" reactiontime="+108" swimtime="00:01:15.91" resultid="5981" heatid="7810" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="295" reactiontime="+113" swimtime="00:02:47.40" resultid="5982" heatid="7956" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="325" reactiontime="+101" swimtime="00:05:52.41" resultid="5983" heatid="9066" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:02:05.45" />
                    <SPLIT distance="200" swimtime="00:02:50.24" />
                    <SPLIT distance="250" swimtime="00:03:35.63" />
                    <SPLIT distance="300" swimtime="00:04:21.23" />
                    <SPLIT distance="350" swimtime="00:05:07.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Wodnik 29 Katowice C" number="2">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+83" swimtime="00:01:45.54" resultid="5985" heatid="7974" lane="7" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                    <SPLIT distance="100" swimtime="00:00:56.17" />
                    <SPLIT distance="150" swimtime="00:01:21.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5882" number="1" />
                    <RELAYPOSITION athleteid="5946" number="2" />
                    <RELAYPOSITION athleteid="5960" number="3" />
                    <RELAYPOSITION athleteid="5951" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Wodnik 29 Katowice D" number="4">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+78" swimtime="00:02:15.21" resultid="5988" heatid="7870" lane="6" entrytime="00:02:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                    <SPLIT distance="150" swimtime="00:01:43.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5882" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="5891" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="5864" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="5946" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Wodnik 29 Katowice B" number="3">
              <RESULTS>
                <RESULT eventid="1495" reactiontime="+90" swimtime="00:02:23.30" resultid="5986" heatid="7968" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                    <SPLIT distance="150" swimtime="00:01:52.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5941" number="1" />
                    <RELAYPOSITION athleteid="5897" number="2" />
                    <RELAYPOSITION athleteid="5935" number="3" />
                    <RELAYPOSITION athleteid="5871" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" reactiontime="+76" swimtime="00:02:42.37" resultid="5987" heatid="7867" lane="8" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                    <SPLIT distance="100" swimtime="00:01:31.93" />
                    <SPLIT distance="150" swimtime="00:02:05.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5927" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="5935" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="5871" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="5897" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Wodnik 29 Katowice B" number="1">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+84" swimtime="00:02:03.63" resultid="5984" heatid="8052" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                    <SPLIT distance="150" swimtime="00:01:33.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5941" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="5960" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="5951" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="5871" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01711" nation="POL" region="11" clubid="2600" name="UKS Wodnik Siemianowice Śl." shortname="Wodnik Siemianowice Śl.">
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="2601">
              <RESULTS>
                <RESULT eventid="1156" points="528" swimtime="00:22:01.12" resultid="2602" heatid="8719" lane="4" entrytime="00:21:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:20.83" />
                    <SPLIT distance="200" swimtime="00:02:50.73" />
                    <SPLIT distance="300" swimtime="00:04:20.38" />
                    <SPLIT distance="400" swimtime="00:05:49.99" />
                    <SPLIT distance="500" swimtime="00:07:20.23" />
                    <SPLIT distance="600" swimtime="00:08:49.00" />
                    <SPLIT distance="700" swimtime="00:10:18.00" />
                    <SPLIT distance="800" swimtime="00:11:47.63" />
                    <SPLIT distance="900" swimtime="00:13:17.40" />
                    <SPLIT distance="1000" swimtime="00:14:46.64" />
                    <SPLIT distance="1100" swimtime="00:16:14.19" />
                    <SPLIT distance="1200" swimtime="00:17:43.15" />
                    <SPLIT distance="1300" swimtime="00:19:11.29" />
                    <SPLIT distance="1400" swimtime="00:20:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="473" reactiontime="+87" swimtime="00:00:35.35" resultid="2603" heatid="7913" lane="8" entrytime="00:00:35.14" />
                <RESULT eventid="1543" points="513" reactiontime="+101" swimtime="00:06:25.01" resultid="2604" heatid="8809" lane="5" entrytime="00:06:22.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:32.81" />
                    <SPLIT distance="150" swimtime="00:02:23.16" />
                    <SPLIT distance="200" swimtime="00:03:12.52" />
                    <SPLIT distance="250" swimtime="00:04:07.74" />
                    <SPLIT distance="300" swimtime="00:05:02.97" />
                    <SPLIT distance="350" swimtime="00:05:44.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" nation="POL" region="14" clubid="4389" name="Ursynów Masters">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1985-05-26" firstname="Urszula" gender="F" lastname="Grycz" nation="POL" athleteid="4408">
              <RESULTS>
                <RESULT eventid="1140" points="431" swimtime="00:12:16.41" resultid="4409" heatid="8713" lane="3" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                    <SPLIT distance="100" swimtime="00:01:25.04" />
                    <SPLIT distance="200" swimtime="00:02:56.19" />
                    <SPLIT distance="300" swimtime="00:04:29.12" />
                    <SPLIT distance="400" swimtime="00:06:02.45" />
                    <SPLIT distance="500" swimtime="00:07:36.76" />
                    <SPLIT distance="600" swimtime="00:09:11.26" />
                    <SPLIT distance="700" swimtime="00:10:45.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="522" reactiontime="+91" swimtime="00:01:12.49" resultid="4410" heatid="7803" lane="1" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="404" reactiontime="+95" swimtime="00:01:35.53" resultid="4411" heatid="7878" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="481" reactiontime="+97" swimtime="00:02:40.82" resultid="4412" heatid="7949" lane="7" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:01:59.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="455" reactiontime="+87" swimtime="00:05:48.26" resultid="4413" heatid="9050" lane="4" entrytime="00:05:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:21.30" />
                    <SPLIT distance="150" swimtime="00:02:05.31" />
                    <SPLIT distance="200" swimtime="00:02:49.96" />
                    <SPLIT distance="250" swimtime="00:03:35.11" />
                    <SPLIT distance="300" swimtime="00:04:20.68" />
                    <SPLIT distance="350" swimtime="00:05:05.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-03" firstname="Alicja" gender="F" lastname="Cicha-Mikołajczyk" nation="POL" athleteid="4414">
              <RESULTS>
                <RESULT eventid="1431" status="DNS" swimtime="00:00:00.00" resultid="4415" heatid="7926" lane="3" entrytime="00:02:25.00" />
                <RESULT eventid="1463" points="142" reactiontime="+134" swimtime="00:04:15.97" resultid="4416" heatid="7944" lane="3" entrytime="00:04:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.37" />
                    <SPLIT distance="100" swimtime="00:02:06.19" />
                    <SPLIT distance="150" swimtime="00:03:14.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="125" reactiontime="+89" swimtime="00:05:06.74" resultid="4417" heatid="8004" lane="4" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.49" />
                    <SPLIT distance="100" swimtime="00:02:31.68" />
                    <SPLIT distance="150" swimtime="00:03:50.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="147" reactiontime="+124" swimtime="00:08:57.57" resultid="4418" heatid="9052" lane="1" entrytime="00:08:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.48" />
                    <SPLIT distance="100" swimtime="00:02:05.96" />
                    <SPLIT distance="150" swimtime="00:03:14.82" />
                    <SPLIT distance="200" swimtime="00:04:24.50" />
                    <SPLIT distance="250" swimtime="00:05:34.06" />
                    <SPLIT distance="300" swimtime="00:06:44.40" />
                    <SPLIT distance="350" swimtime="00:07:54.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="Nowak" nation="POL" athleteid="4419">
              <RESULTS>
                <RESULT eventid="1108" points="763" reactiontime="+88" swimtime="00:02:59.73" resultid="4420" heatid="7725" lane="3" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:01:27.05" />
                    <SPLIT distance="150" swimtime="00:02:17.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="828" reactiontime="+90" swimtime="00:03:06.31" resultid="4421" heatid="7792" lane="5" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:27.50" />
                    <SPLIT distance="150" swimtime="00:02:15.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="806" reactiontime="+74" swimtime="00:01:17.83" resultid="4422" heatid="7846" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="891" reactiontime="+79" swimtime="00:01:21.19" resultid="4423" heatid="7891" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="592" reactiontime="+83" swimtime="00:06:55.26" resultid="4424" heatid="8810" lane="4" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:01:38.03" />
                    <SPLIT distance="150" swimtime="00:03:22.60" />
                    <SPLIT distance="200" swimtime="00:04:17.81" />
                    <SPLIT distance="250" swimtime="00:05:13.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="395" reactiontime="+90" swimtime="00:01:33.08" resultid="4425" heatid="7996" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="815" reactiontime="+74" swimtime="00:00:36.19" resultid="4426" heatid="8041" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="Rybarczyk" nation="POL" athleteid="4427">
              <RESULTS>
                <RESULT eventid="1076" points="513" reactiontime="+90" swimtime="00:00:29.68" resultid="4428" heatid="7699" lane="4" entrytime="00:00:29.57" />
                <RESULT eventid="1190" points="240" reactiontime="+79" swimtime="00:00:43.63" resultid="4429" heatid="7767" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="1254" points="506" reactiontime="+93" swimtime="00:01:05.34" resultid="4430" heatid="7817" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="468" reactiontime="+90" swimtime="00:00:32.35" resultid="4431" heatid="7914" lane="5" entrytime="00:00:33.64" />
                <RESULT eventid="1479" points="415" reactiontime="+89" swimtime="00:02:31.48" resultid="4432" heatid="7960" lane="3" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:10.58" />
                    <SPLIT distance="150" swimtime="00:01:51.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="357" reactiontime="+91" swimtime="00:01:19.76" resultid="4433" heatid="7997" lane="8" entrytime="00:01:21.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="389" reactiontime="+98" swimtime="00:05:29.53" resultid="4434" heatid="9067" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:15.09" />
                    <SPLIT distance="150" swimtime="00:01:56.98" />
                    <SPLIT distance="200" swimtime="00:02:40.17" />
                    <SPLIT distance="250" swimtime="00:03:23.36" />
                    <SPLIT distance="300" swimtime="00:04:07.12" />
                    <SPLIT distance="350" swimtime="00:04:50.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-03-23" firstname="Ryszard" gender="M" lastname="Rybarczyk" nation="POL" athleteid="4435">
              <RESULTS>
                <RESULT eventid="1076" points="356" reactiontime="+101" swimtime="00:00:40.89" resultid="4436" heatid="7686" lane="8" entrytime="00:00:41.75" />
                <RESULT eventid="1190" points="271" reactiontime="+94" swimtime="00:00:53.57" resultid="4437" heatid="7764" lane="4" entrytime="00:00:53.85" />
                <RESULT eventid="1222" points="477" reactiontime="+99" swimtime="00:03:57.05" resultid="4438" heatid="7786" lane="2" entrytime="00:04:09.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.64" />
                    <SPLIT distance="100" swimtime="00:01:55.73" />
                    <SPLIT distance="150" swimtime="00:03:00.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="4439" heatid="7883" lane="2" entrytime="00:01:47.47" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="4440" heatid="7952" lane="6" entrytime="00:05:42.58" />
                <RESULT eventid="1655" points="504" reactiontime="+102" swimtime="00:00:47.03" resultid="4441" heatid="8032" lane="3" entrytime="00:00:45.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-11" firstname="Maciej" gender="M" lastname="Rybicki" nation="POL" athleteid="4442">
              <RESULTS>
                <RESULT eventid="1076" status="WDR" swimtime="00:00:00.00" resultid="4443" heatid="7696" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="1190" status="WDR" swimtime="00:00:00.00" resultid="4444" heatid="7769" lane="1" entrytime="00:00:40.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VIELB" nation="POL" region="13" clubid="3123" name="Victory Masters Elbląg">
          <CONTACT name="Latecki Grzegorz" street="Łokietka 45" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="3124">
              <RESULTS>
                <RESULT eventid="1059" points="242" reactiontime="+97" swimtime="00:00:42.54" resultid="3125" heatid="7674" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1140" points="256" reactiontime="+102" swimtime="00:14:35.52" resultid="3126" heatid="8712" lane="8" entrytime="00:12:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.62" />
                    <SPLIT distance="100" swimtime="00:01:41.71" />
                    <SPLIT distance="150" swimtime="00:04:27.41" />
                    <SPLIT distance="200" swimtime="00:05:22.99" />
                    <SPLIT distance="250" swimtime="00:06:18.62" />
                    <SPLIT distance="300" swimtime="00:09:07.57" />
                    <SPLIT distance="350" swimtime="00:11:54.15" />
                    <SPLIT distance="400" swimtime="00:12:49.74" />
                    <SPLIT distance="450" swimtime="00:13:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="231" reactiontime="+91" swimtime="00:01:35.15" resultid="3127" heatid="7798" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="245" reactiontime="+107" swimtime="00:03:21.22" resultid="3128" heatid="7946" lane="5" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                    <SPLIT distance="100" swimtime="00:01:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="243" reactiontime="+103" swimtime="00:07:09.18" resultid="3129" heatid="9052" lane="5" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                    <SPLIT distance="150" swimtime="00:03:35.61" />
                    <SPLIT distance="200" swimtime="00:04:31.36" />
                    <SPLIT distance="250" swimtime="00:05:25.60" />
                    <SPLIT distance="300" swimtime="00:06:19.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karaś" nation="POL" athleteid="3130">
              <RESULTS>
                <RESULT eventid="1092" points="270" reactiontime="+109" swimtime="00:04:00.28" resultid="3131" heatid="7714" lane="5" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.65" />
                    <SPLIT distance="100" swimtime="00:01:56.52" />
                    <SPLIT distance="150" swimtime="00:03:09.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="303" swimtime="00:14:30.36" resultid="3132" heatid="8715" lane="4" entrytime="00:14:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.26" />
                    <SPLIT distance="100" swimtime="00:01:49.15" />
                    <SPLIT distance="200" swimtime="00:03:39.33" />
                    <SPLIT distance="300" swimtime="00:05:29.38" />
                    <SPLIT distance="400" swimtime="00:07:19.04" />
                    <SPLIT distance="500" swimtime="00:09:08.02" />
                    <SPLIT distance="600" swimtime="00:10:56.74" />
                    <SPLIT distance="700" swimtime="00:12:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="278" reactiontime="+115" swimtime="00:01:34.85" resultid="3133" heatid="7798" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="321" reactiontime="+114" swimtime="00:04:08.59" resultid="3134" heatid="7857" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                    <SPLIT distance="100" swimtime="00:01:57.97" />
                    <SPLIT distance="150" swimtime="00:03:03.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="276" reactiontime="+115" swimtime="00:03:27.00" resultid="3135" heatid="7946" lane="8" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                    <SPLIT distance="100" swimtime="00:01:40.77" />
                    <SPLIT distance="150" swimtime="00:02:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="291" reactiontime="+116" swimtime="00:08:26.88" resultid="3136" heatid="8803" lane="8" entrytime="00:08:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.41" />
                    <SPLIT distance="100" swimtime="00:01:58.11" />
                    <SPLIT distance="150" swimtime="00:03:05.76" />
                    <SPLIT distance="200" swimtime="00:04:09.95" />
                    <SPLIT distance="250" swimtime="00:05:24.58" />
                    <SPLIT distance="300" swimtime="00:06:41.02" />
                    <SPLIT distance="350" swimtime="00:07:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="231" reactiontime="+100" swimtime="00:01:55.23" resultid="3137" heatid="7989" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="301" reactiontime="+101" swimtime="00:07:06.82" resultid="3138" heatid="9052" lane="6" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.51" />
                    <SPLIT distance="100" swimtime="00:01:40.56" />
                    <SPLIT distance="150" swimtime="00:02:35.50" />
                    <SPLIT distance="200" swimtime="00:03:29.64" />
                    <SPLIT distance="250" swimtime="00:04:24.60" />
                    <SPLIT distance="300" swimtime="00:05:19.80" />
                    <SPLIT distance="350" swimtime="00:06:14.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner Mateusiak" nation="POL" athleteid="3139">
              <RESULTS>
                <RESULT eventid="1059" points="225" reactiontime="+136" swimtime="00:00:49.73" resultid="3140" heatid="7672" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1173" points="197" reactiontime="+97" swimtime="00:01:02.53" resultid="3141" heatid="7754" lane="2" entrytime="00:01:10.00" />
                <RESULT eventid="1238" points="175" swimtime="00:02:02.40" resultid="3142" heatid="7797" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.83" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K15 - Brak dotknięcia ściany obydwoma rozłączonymi dłońmi przy nawrocie lub na zakończenie wyścigu" eventid="1366" reactiontime="+110" status="DSQ" swimtime="00:02:36.47" resultid="3143" heatid="7874" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" status="DNS" swimtime="00:00:00.00" resultid="3144" heatid="7926" lane="6" entrytime="00:02:33.00" />
                <RESULT eventid="1639" points="149" reactiontime="+112" swimtime="00:01:10.72" resultid="3145" heatid="8021" lane="7" entrytime="00:01:07.00" />
                <RESULT eventid="1140" status="DNF" swimtime="00:00:00.00" resultid="6141" heatid="8715" lane="1" entrytime="00:18:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOPKK" nation="POL" region="07" clubid="2192" name="WOPR Kędzierzyn Koźle">
          <ATHLETES>
            <ATHLETE birthdate="1959-07-07" firstname="Ryszard" gender="M" lastname="Tatarczuk" nation="POL" athleteid="2193">
              <RESULTS>
                <RESULT eventid="1076" points="424" reactiontime="+89" swimtime="00:00:33.81" resultid="2194" heatid="7691" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1156" points="326" swimtime="00:25:50.89" resultid="2195" heatid="8723" lane="5" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:01:31.41" />
                    <SPLIT distance="200" swimtime="00:03:12.41" />
                    <SPLIT distance="300" swimtime="00:04:52.82" />
                    <SPLIT distance="400" swimtime="00:06:36.06" />
                    <SPLIT distance="500" swimtime="00:08:20.88" />
                    <SPLIT distance="600" swimtime="00:10:05.18" />
                    <SPLIT distance="700" swimtime="00:11:50.03" />
                    <SPLIT distance="800" swimtime="00:13:36.41" />
                    <SPLIT distance="900" swimtime="00:15:21.42" />
                    <SPLIT distance="1000" swimtime="00:17:07.21" />
                    <SPLIT distance="1100" swimtime="00:18:52.28" />
                    <SPLIT distance="1200" swimtime="00:20:37.80" />
                    <SPLIT distance="1300" swimtime="00:22:23.57" />
                    <SPLIT distance="1400" swimtime="00:24:10.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-11-01" firstname="Stanisław" gender="M" lastname="Zajfert" nation="POL" athleteid="2196">
              <RESULTS>
                <RESULT eventid="1076" points="477" reactiontime="+93" swimtime="00:00:36.05" resultid="2197" heatid="7688" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1156" points="534" swimtime="00:27:07.94" resultid="2198" heatid="8723" lane="3" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                    <SPLIT distance="100" swimtime="00:01:36.54" />
                    <SPLIT distance="200" swimtime="00:03:24.26" />
                    <SPLIT distance="300" swimtime="00:05:12.31" />
                    <SPLIT distance="400" swimtime="00:07:01.45" />
                    <SPLIT distance="500" swimtime="00:08:51.39" />
                    <SPLIT distance="600" swimtime="00:10:41.71" />
                    <SPLIT distance="700" swimtime="00:12:32.90" />
                    <SPLIT distance="800" swimtime="00:14:24.39" />
                    <SPLIT distance="900" swimtime="00:16:13.71" />
                    <SPLIT distance="1000" swimtime="00:18:03.02" />
                    <SPLIT distance="1100" swimtime="00:19:51.43" />
                    <SPLIT distance="1200" swimtime="00:21:42.17" />
                    <SPLIT distance="1300" swimtime="00:23:32.99" />
                    <SPLIT distance="1400" swimtime="00:02:52.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="5225" name="Warsaw Masters Team">
          <CONTACT city="Warszawa" email="wojciech.kaluzynski@gmail.com" internet="www.masters.waw.pl" name="Kałużyński Wojciech" phone="607 45 44 44" state="MAZ" />
          <ATHLETES>
            <ATHLETE birthdate="1986-04-21" firstname="Marianna" gender="F" lastname="Gajdus" nation="POL" athleteid="5233">
              <RESULTS>
                <RESULT eventid="1206" points="441" reactiontime="+78" swimtime="00:03:21.80" resultid="5234" heatid="7782" lane="5" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.75" />
                    <SPLIT distance="100" swimtime="00:01:36.98" />
                    <SPLIT distance="150" swimtime="00:02:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="528" reactiontime="+81" swimtime="00:01:20.91" resultid="5235" heatid="7835" lane="3" entrytime="00:01:19.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="569" reactiontime="+73" swimtime="00:00:35.07" resultid="5236" heatid="7902" lane="4" entrytime="00:00:35.21" entrycourse="SCM" />
                <RESULT eventid="1463" points="477" reactiontime="+84" swimtime="00:02:41.28" resultid="5237" heatid="7949" lane="3" entrytime="00:02:40.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="100" swimtime="00:01:18.30" />
                    <SPLIT distance="150" swimtime="00:02:00.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="503" reactiontime="+77" swimtime="00:01:20.43" resultid="5238" heatid="7990" lane="6" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="467" reactiontime="+79" swimtime="00:05:45.14" resultid="5239" heatid="9048" lane="4" entrytime="00:05:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                    <SPLIT distance="100" swimtime="00:01:21.12" />
                    <SPLIT distance="150" swimtime="00:02:05.44" />
                    <SPLIT distance="200" swimtime="00:02:50.48" />
                    <SPLIT distance="250" swimtime="00:03:35.32" />
                    <SPLIT distance="300" swimtime="00:04:20.30" />
                    <SPLIT distance="350" swimtime="00:05:04.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-14" firstname="Wojciech" gender="M" lastname="Kałużyński" nation="POL" athleteid="5240">
              <RESULTS>
                <RESULT eventid="1108" points="281" reactiontime="+83" swimtime="00:03:00.32" resultid="5241" heatid="7725" lane="4" entrytime="00:03:01.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:01:24.62" />
                    <SPLIT distance="150" swimtime="00:02:18.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="384" reactiontime="+82" swimtime="00:01:07.43" resultid="5242" heatid="7815" lane="5" entrytime="00:01:06.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="323" reactiontime="+91" swimtime="00:01:20.09" resultid="5243" heatid="7846" lane="3" entrytime="00:01:18.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="226" reactiontime="+92" swimtime="00:00:37.50" resultid="5244" heatid="7906" lane="7" />
                <RESULT eventid="1479" points="297" reactiontime="+88" swimtime="00:02:39.51" resultid="5245" heatid="7961" lane="8" entrytime="00:02:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:01:13.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="5246" heatid="8032" lane="5" entrytime="00:00:45.37" entrycourse="SCM" />
                <RESULT eventid="1703" points="362" reactiontime="+87" swimtime="00:05:36.90" resultid="5247" heatid="9064" lane="5" entrytime="00:05:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:18.69" />
                    <SPLIT distance="150" swimtime="00:02:01.26" />
                    <SPLIT distance="200" swimtime="00:02:44.48" />
                    <SPLIT distance="250" swimtime="00:03:27.70" />
                    <SPLIT distance="300" swimtime="00:04:11.18" />
                    <SPLIT distance="350" swimtime="00:04:55.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="5248">
              <RESULTS>
                <RESULT eventid="1108" points="294" reactiontime="+113" swimtime="00:04:45.78" resultid="5249" heatid="7720" lane="7" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.73" />
                    <SPLIT distance="100" swimtime="00:02:26.93" />
                    <SPLIT distance="150" swimtime="00:03:40.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="351" reactiontime="+119" swimtime="00:04:37.18" resultid="5250" heatid="7785" lane="6" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.39" />
                    <SPLIT distance="100" swimtime="00:02:17.89" />
                    <SPLIT distance="150" swimtime="00:03:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="176" reactiontime="+114" swimtime="00:06:08.64" resultid="5251" heatid="7859" lane="7" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.59" />
                    <SPLIT distance="100" swimtime="00:02:58.09" />
                    <SPLIT distance="150" swimtime="00:04:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="251" reactiontime="+115" swimtime="00:00:58.87" resultid="5252" heatid="7906" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1543" points="309" reactiontime="+126" swimtime="00:10:09.81" resultid="5253" heatid="8812" lane="3" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.89" />
                    <SPLIT distance="100" swimtime="00:02:44.35" />
                    <SPLIT distance="150" swimtime="00:04:03.69" />
                    <SPLIT distance="200" swimtime="00:05:22.34" />
                    <SPLIT distance="250" swimtime="00:06:38.58" />
                    <SPLIT distance="300" swimtime="00:07:55.86" />
                    <SPLIT distance="350" swimtime="00:09:03.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="194" reactiontime="+116" swimtime="00:02:39.00" resultid="5254" heatid="7992" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G8 - Ukończenie wyścigu nie w położeniu na plecach" eventid="1623" reactiontime="+85" status="DSQ" swimtime="00:04:45.97" resultid="5255" heatid="8010" lane="6" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.44" />
                    <SPLIT distance="100" swimtime="00:02:20.40" />
                    <SPLIT distance="150" swimtime="00:03:33.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-09" firstname="Alina" gender="F" lastname="Wieczorkiewicz" nation="POL" athleteid="5256">
              <RESULTS>
                <RESULT eventid="1092" points="111" reactiontime="+108" swimtime="00:06:39.65" resultid="5257" heatid="7713" lane="5" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:41.05" />
                    <SPLIT distance="100" swimtime="00:03:12.78" />
                    <SPLIT distance="150" swimtime="00:05:01.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="153" reactiontime="+96" swimtime="00:01:18.14" resultid="5258" heatid="7753" lane="4" entrytime="00:01:25.00" />
                <RESULT eventid="1270" points="105" reactiontime="+106" swimtime="00:03:05.20" resultid="5259" heatid="7826" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="108" reactiontime="+108" swimtime="00:03:23.49" resultid="5260" heatid="7874" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G3 - Nieutrzymanie pozycji na plecach (z wyjątkiem wykonania cyklu nawrotu)" eventid="1431" status="DSQ" swimtime="00:00:00.00" resultid="5261" heatid="7926" lane="7" entrytime="00:02:50.00" />
                <RESULT eventid="1607" points="139" reactiontime="+93" swimtime="00:06:21.15" resultid="5262" heatid="8004" lane="5" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.25" />
                    <SPLIT distance="100" swimtime="00:03:06.06" />
                    <SPLIT distance="150" swimtime="00:04:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="108" reactiontime="+114" swimtime="00:01:30.51" resultid="5263" heatid="8021" lane="8" entrytime="00:01:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="5264">
              <RESULTS>
                <RESULT eventid="1076" points="300" reactiontime="+105" swimtime="00:00:37.94" resultid="5265" heatid="7688" lane="8" entrytime="00:00:36.41" />
                <RESULT eventid="1190" points="165" reactiontime="+107" swimtime="00:00:53.46" resultid="5266" heatid="7765" lane="8" entrytime="00:00:52.35" />
                <RESULT eventid="1286" points="238" reactiontime="+98" swimtime="00:01:45.66" resultid="5267" heatid="7838" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="196" reactiontime="+107" swimtime="00:00:47.39" resultid="5268" heatid="7908" lane="7" entrytime="00:00:44.64" />
                <RESULT eventid="1479" points="287" reactiontime="+107" swimtime="00:03:10.57" resultid="5269" heatid="7955" lane="8" entrytime="00:03:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:29.27" />
                    <SPLIT distance="150" swimtime="00:02:20.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="265" reactiontime="+102" swimtime="00:06:54.50" resultid="5270" heatid="9061" lane="8" entrytime="00:05:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:01:32.58" />
                    <SPLIT distance="150" swimtime="00:02:26.37" />
                    <SPLIT distance="250" swimtime="00:04:17.14" />
                    <SPLIT distance="300" swimtime="00:05:13.38" />
                    <SPLIT distance="350" swimtime="00:06:07.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="5271">
              <RESULTS>
                <RESULT eventid="1076" points="283" reactiontime="+102" swimtime="00:00:36.82" resultid="5272" heatid="7688" lane="7" entrytime="00:00:36.01" />
                <RESULT eventid="1222" points="376" reactiontime="+101" swimtime="00:03:26.71" resultid="5273" heatid="7790" lane="2" entrytime="00:03:22.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:37.82" />
                    <SPLIT distance="150" swimtime="00:02:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="353" reactiontime="+106" swimtime="00:01:35.06" resultid="5274" heatid="7881" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="242" reactiontime="+100" swimtime="00:00:42.41" resultid="5275" heatid="7908" lane="3" entrytime="00:00:43.08" />
                <RESULT eventid="1591" points="162" reactiontime="+94" swimtime="00:01:47.72" resultid="5276" heatid="7993" lane="2" entrytime="00:01:53.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="344" reactiontime="+91" swimtime="00:00:43.75" resultid="5277" heatid="8034" lane="4" entrytime="00:00:42.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-28" firstname="Katarzyna" gender="F" lastname="Dobczyńska" nation="POL" athleteid="5278">
              <RESULTS>
                <RESULT eventid="1059" points="368" reactiontime="+110" swimtime="00:00:37.89" resultid="5279" heatid="7675" lane="7" entrytime="00:00:39.91" />
                <RESULT eventid="1173" points="411" reactiontime="+101" swimtime="00:00:42.89" resultid="5280" heatid="7755" lane="4" entrytime="00:00:46.90" />
                <RESULT eventid="1238" points="325" reactiontime="+109" swimtime="00:01:24.00" resultid="5281" heatid="7800" lane="3" entrytime="00:01:22.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="383" reactiontime="+91" swimtime="00:01:30.71" resultid="5282" heatid="7928" lane="2" entrytime="00:01:33.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="351" reactiontime="+112" swimtime="00:03:01.46" resultid="5283" heatid="7947" lane="7" entrytime="00:03:06.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                    <SPLIT distance="100" swimtime="00:01:28.40" />
                    <SPLIT distance="150" swimtime="00:02:15.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="383" reactiontime="+104" swimtime="00:03:16.51" resultid="5284" heatid="8006" lane="7" entrytime="00:03:20.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:36.96" />
                    <SPLIT distance="150" swimtime="00:02:28.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-18" firstname="Robert" gender="M" lastname="Nowicki" nation="POL" athleteid="5285">
              <RESULTS>
                <RESULT eventid="1076" points="259" reactiontime="+105" swimtime="00:00:39.84" resultid="5286" heatid="7686" lane="3" entrytime="00:00:40.90" />
                <RESULT eventid="1156" status="WDR" swimtime="00:00:00.00" resultid="5287" entrytime="00:29:23.49" />
                <RESULT eventid="1254" points="247" reactiontime="+112" swimtime="00:01:29.93" resultid="5288" heatid="7807" lane="4" entrytime="00:01:31.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="247" reactiontime="+111" swimtime="00:03:20.33" resultid="5289" heatid="7953" lane="5" entrytime="00:03:22.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:34.68" />
                    <SPLIT distance="150" swimtime="00:02:27.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="5290">
              <RESULTS>
                <RESULT eventid="1076" points="869" reactiontime="+73" swimtime="00:00:26.62" resultid="5291" heatid="7708" lane="2" entrytime="00:00:26.78" />
                <RESULT eventid="1254" points="954" reactiontime="+77" swimtime="00:00:57.32" resultid="5292" heatid="7806" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="950" reactiontime="+77" swimtime="00:01:06.61" resultid="5293" heatid="7854" lane="8" entrytime="00:01:07.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="5294" heatid="7966" lane="8" entrytime="00:02:11.12" />
                <RESULT eventid="1655" points="765" reactiontime="+78" swimtime="00:00:34.30" resultid="5295" heatid="8043" lane="2" entrytime="00:00:35.78" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-07" firstname="Michał" gender="M" lastname="Wasielak" nation="POL" athleteid="5296">
              <RESULTS>
                <RESULT eventid="1076" points="306" reactiontime="+93" swimtime="00:00:32.81" resultid="5297" heatid="7692" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1254" points="280" reactiontime="+89" swimtime="00:01:14.88" resultid="5298" heatid="7811" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="274" reactiontime="+112" swimtime="00:02:43.94" resultid="5299" heatid="7957" lane="7" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:18.40" />
                    <SPLIT distance="150" swimtime="00:02:02.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="310" reactiontime="+88" swimtime="00:05:54.96" resultid="5300" heatid="9067" lane="3" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:01:19.71" />
                    <SPLIT distance="150" swimtime="00:02:03.65" />
                    <SPLIT distance="200" swimtime="00:02:48.77" />
                    <SPLIT distance="250" swimtime="00:03:35.66" />
                    <SPLIT distance="300" swimtime="00:04:22.76" />
                    <SPLIT distance="350" swimtime="00:05:09.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-12-16" firstname="Przemysław" gender="M" lastname="Wołosz" nation="POL" athleteid="5301">
              <RESULTS>
                <RESULT eventid="1286" points="383" reactiontime="+83" swimtime="00:01:21.31" resultid="5302" heatid="7843" lane="1" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="381" reactiontime="+92" swimtime="00:01:28.25" resultid="5303" heatid="7888" lane="6" entrytime="00:01:29.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="403" reactiontime="+83" swimtime="00:00:34.72" resultid="5304" heatid="7912" lane="3" entrytime="00:00:35.62" />
                <RESULT eventid="1447" points="315" reactiontime="+89" swimtime="00:01:26.81" resultid="5305" heatid="7937" lane="1" entrytime="00:01:25.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-20" firstname="Anna" gender="F" lastname="Stanisławska" nation="POL" athleteid="5306">
              <RESULTS>
                <RESULT eventid="1059" points="386" reactiontime="+100" swimtime="00:00:36.40" resultid="5307" heatid="7676" lane="5" entrytime="00:00:36.74" />
                <RESULT eventid="1140" points="354" swimtime="00:13:06.12" resultid="5308" heatid="8714" lane="3" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="100" swimtime="00:01:29.96" />
                    <SPLIT distance="200" swimtime="00:03:07.65" />
                    <SPLIT distance="300" swimtime="00:04:47.50" />
                    <SPLIT distance="400" swimtime="00:06:28.38" />
                    <SPLIT distance="500" swimtime="00:08:09.51" />
                    <SPLIT distance="600" swimtime="00:09:49.41" />
                    <SPLIT distance="700" swimtime="00:11:29.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="384" reactiontime="+105" swimtime="00:01:20.28" resultid="5309" heatid="7799" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="287" reactiontime="+123" swimtime="00:03:33.29" resultid="5310" heatid="7858" lane="2" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.23" />
                    <SPLIT distance="100" swimtime="00:01:39.01" />
                    <SPLIT distance="150" swimtime="00:02:35.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="356" reactiontime="+111" swimtime="00:00:41.01" resultid="5311" heatid="7899" lane="6" entrytime="00:00:41.38" />
                <RESULT eventid="1527" points="332" reactiontime="+111" swimtime="00:07:19.43" resultid="5312" heatid="8803" lane="2" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                    <SPLIT distance="100" swimtime="00:01:38.02" />
                    <SPLIT distance="150" swimtime="00:02:40.19" />
                    <SPLIT distance="200" swimtime="00:03:38.66" />
                    <SPLIT distance="250" swimtime="00:04:38.82" />
                    <SPLIT distance="300" swimtime="00:05:41.91" />
                    <SPLIT distance="350" swimtime="00:06:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="272" reactiontime="+121" swimtime="00:01:38.72" resultid="5313" heatid="7988" lane="7" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="318" reactiontime="+125" swimtime="00:06:32.14" resultid="5314" heatid="9051" lane="3" entrytime="00:06:27.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.57" />
                    <SPLIT distance="100" swimtime="00:01:32.12" />
                    <SPLIT distance="150" swimtime="00:02:23.25" />
                    <SPLIT distance="200" swimtime="00:03:13.43" />
                    <SPLIT distance="250" swimtime="00:04:03.61" />
                    <SPLIT distance="300" swimtime="00:04:54.46" />
                    <SPLIT distance="350" swimtime="00:05:43.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-10-02" firstname="Andrzej" gender="M" lastname="Wiszniewski" nation="POL" athleteid="5315">
              <RESULTS>
                <RESULT eventid="1076" points="243" reactiontime="+105" swimtime="00:00:40.67" resultid="5316" heatid="7686" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1108" points="251" reactiontime="+107" swimtime="00:03:46.49" resultid="5317" heatid="7721" lane="3" entrytime="00:03:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.78" />
                    <SPLIT distance="100" swimtime="00:01:59.81" />
                    <SPLIT distance="150" swimtime="00:02:59.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="317" reactiontime="+108" swimtime="00:03:46.79" resultid="5318" heatid="7788" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.36" />
                    <SPLIT distance="100" swimtime="00:01:49.97" />
                    <SPLIT distance="150" swimtime="00:02:49.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="231" reactiontime="+104" swimtime="00:03:53.29" resultid="5319" heatid="7861" lane="1" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.41" />
                    <SPLIT distance="100" swimtime="00:01:54.13" />
                    <SPLIT distance="150" swimtime="00:02:55.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="156" reactiontime="+83" swimtime="00:02:00.44" resultid="5320" heatid="7933" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="WDR" swimtime="00:00:00.00" resultid="5321" entrytime="00:08:30.00" />
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="5322" heatid="8011" lane="1" entrytime="00:04:20.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="5323" heatid="8031" lane="4" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-11-09" firstname="Tadeusz" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="5324">
              <RESULTS>
                <RESULT eventid="1076" points="537" reactiontime="+130" swimtime="00:00:39.35" resultid="5325" heatid="7686" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-22" firstname="Karol" gender="M" lastname="Dzięcioł" nation="POL" athleteid="5326">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)  (Czas: 17:00)" eventid="1076" reactiontime="+51" status="DSQ" swimtime="00:00:25.38" resultid="5327" heatid="7711" lane="5" entrytime="00:00:25.48" />
                <RESULT eventid="1254" points="675" reactiontime="+74" swimtime="00:00:55.89" resultid="5328" heatid="7825" lane="8" entrytime="00:00:55.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="5329">
              <RESULTS>
                <RESULT eventid="1092" points="359" reactiontime="+84" swimtime="00:03:21.13" resultid="6462" heatid="7715" lane="2" entrytime="00:03:18.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:01:34.41" />
                    <SPLIT distance="150" swimtime="00:02:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="371" reactiontime="+91" swimtime="00:01:30.58" resultid="6463" heatid="7831" lane="1" entrytime="00:01:30.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="367" reactiontime="+89" swimtime="00:00:40.57" resultid="6464" heatid="7900" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1687" points="389" reactiontime="+90" swimtime="00:06:14.65" resultid="6465" heatid="9050" lane="1" entrytime="00:06:20.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:01:27.70" />
                    <SPLIT distance="150" swimtime="00:02:14.67" />
                    <SPLIT distance="200" swimtime="00:03:02.23" />
                    <SPLIT distance="250" swimtime="00:03:50.20" />
                    <SPLIT distance="300" swimtime="00:04:38.44" />
                    <SPLIT distance="350" swimtime="00:05:27.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-13" firstname="Ewa" gender="F" lastname="Krzyżanowska" nation="POL" athleteid="5334">
              <RESULTS>
                <RESULT eventid="1059" points="552" reactiontime="+103" swimtime="00:00:33.13" resultid="6457" heatid="7680" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1173" points="537" reactiontime="+75" swimtime="00:00:38.91" resultid="6458" heatid="7758" lane="5" entrytime="00:00:39.49" />
                <RESULT eventid="1238" points="488" reactiontime="+110" swimtime="00:01:15.48" resultid="6459" heatid="7802" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="468" reactiontime="+78" swimtime="00:01:27.53" resultid="6460" heatid="7928" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="418" reactiontime="+106" swimtime="00:06:10.25" resultid="6461" heatid="9050" lane="7" entrytime="00:06:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:01:23.42" />
                    <SPLIT distance="150" swimtime="00:02:10.07" />
                    <SPLIT distance="200" swimtime="00:02:58.26" />
                    <SPLIT distance="250" swimtime="00:03:46.86" />
                    <SPLIT distance="300" swimtime="00:05:24.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-02-15" firstname="Anna" gender="F" lastname="MIchalska" nation="POL" athleteid="5340">
              <RESULTS>
                <RESULT eventid="1206" points="503" reactiontime="+81" swimtime="00:03:34.25" resultid="6466" heatid="7781" lane="2" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                    <SPLIT distance="100" swimtime="00:01:44.93" />
                    <SPLIT distance="150" swimtime="00:02:39.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="488" reactiontime="+86" swimtime="00:01:40.18" resultid="6467" heatid="7878" lane="1" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="463" reactiontime="+79" swimtime="00:00:45.78" resultid="6468" heatid="8025" lane="3" entrytime="00:00:45.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="5344">
              <RESULTS>
                <RESULT eventid="1190" points="793" reactiontime="+75" swimtime="00:00:30.96" resultid="5345" heatid="7775" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1286" points="698" reactiontime="+85" swimtime="00:01:08.17" resultid="5346" heatid="7853" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="798" reactiontime="+75" swimtime="00:01:06.99" resultid="5347" heatid="7942" lane="8" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="711" reactiontime="+78" swimtime="00:02:32.69" resultid="5348" heatid="8018" lane="5" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:12.88" />
                    <SPLIT distance="150" swimtime="00:01:53.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-09" firstname="Tomasz" gender="M" lastname="Makomaski" nation="POL" athleteid="5349">
              <RESULTS>
                <RESULT eventid="1076" points="572" reactiontime="+90" swimtime="00:00:27.50" resultid="5350" heatid="7707" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1222" points="451" reactiontime="+90" swimtime="00:03:00.38" resultid="5351" heatid="7794" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:25.93" />
                    <SPLIT distance="150" swimtime="00:02:14.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="472" reactiontime="+91" swimtime="00:01:02.39" resultid="5352" heatid="7819" lane="3" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="518" reactiontime="+91" swimtime="00:01:17.23" resultid="5353" heatid="7893" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="423" reactiontime="+94" swimtime="00:00:31.55" resultid="5354" heatid="7922" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1655" points="551" reactiontime="+87" swimtime="00:00:34.46" resultid="5355" heatid="8046" lane="6" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-30" firstname="Piotr" gender="M" lastname="Safrończyk" nation="POL" athleteid="5356">
              <RESULTS>
                <RESULT eventid="1286" points="831" reactiontime="+67" swimtime="00:00:58.70" resultid="5357" heatid="7856" lane="4" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="910" reactiontime="+70" swimtime="00:01:03.99" resultid="5358" heatid="7896" lane="4" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="944" reactiontime="+65" swimtime="00:00:28.80" resultid="5359" heatid="8048" lane="4" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-06" firstname="Barbara" gender="F" lastname="Tkacz" nation="POL" athleteid="5360">
              <RESULTS>
                <RESULT eventid="1238" points="297" reactiontime="+105" swimtime="00:01:27.50" resultid="5361" heatid="7799" lane="2" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="225" reactiontime="+102" swimtime="00:00:47.75" resultid="5362" heatid="7898" lane="4" entrytime="00:00:46.00" />
                <RESULT eventid="1463" points="241" reactiontime="+106" swimtime="00:03:22.37" resultid="5363" heatid="7946" lane="4" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:01:32.30" />
                    <SPLIT distance="150" swimtime="00:02:26.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" status="DNS" swimtime="00:00:00.00" resultid="5364" heatid="9052" lane="3" entrytime="00:07:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-11-07" firstname="Barbara" gender="F" lastname="Mancewicz" nation="POL" athleteid="5365">
              <RESULTS>
                <RESULT eventid="1270" points="235" reactiontime="+100" swimtime="00:01:45.99" resultid="5366" heatid="7829" lane="1" entrytime="00:01:41.00" />
                <RESULT comment="M8 - Przenoszenie ramion do przodu pod powierzchnią wody podczas ostatniego cyklu pracy ramion przed nawrotem lub na zakończenie wyścigu" eventid="1399" reactiontime="+125" status="DSQ" swimtime="00:00:45.53" resultid="5367" heatid="7898" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="1639" status="DNS" swimtime="00:00:00.00" resultid="5368" heatid="8024" lane="6" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="5369">
              <RESULTS>
                <RESULT eventid="1059" points="497" reactiontime="+87" swimtime="00:00:35.05" resultid="5370" heatid="7679" lane="8" entrytime="00:00:34.10" />
                <RESULT eventid="1206" points="695" reactiontime="+84" swimtime="00:03:12.36" resultid="5371" heatid="7783" lane="7" entrytime="00:03:06.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                    <SPLIT distance="100" swimtime="00:01:34.01" />
                    <SPLIT distance="150" swimtime="00:02:23.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="699" reactiontime="+86" swimtime="00:01:28.88" resultid="5372" heatid="7880" lane="1" entrytime="00:01:26.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" status="DNS" swimtime="00:00:00.00" resultid="5373" heatid="7949" lane="6" entrytime="00:02:41.22" />
                <RESULT eventid="1639" points="698" reactiontime="+82" swimtime="00:00:39.93" resultid="5374" heatid="8028" lane="8" entrytime="00:00:39.43" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-07" firstname="Andrzej" gender="M" lastname="Lewandowski" nation="POL" athleteid="5375">
              <RESULTS>
                <RESULT eventid="1076" points="423" reactiontime="+188" swimtime="00:00:32.21" resultid="5376" heatid="7696" lane="6" entrytime="00:00:30.65" />
                <RESULT eventid="1222" points="488" reactiontime="+96" swimtime="00:03:09.57" resultid="5377" heatid="7791" lane="6" entrytime="00:03:12.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                    <SPLIT distance="100" swimtime="00:01:30.15" />
                    <SPLIT distance="150" swimtime="00:02:20.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="526" reactiontime="+85" swimtime="00:01:23.23" resultid="5378" heatid="7891" lane="7" entrytime="00:01:23.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="626" reactiontime="+76" swimtime="00:00:35.85" resultid="5379" heatid="8043" lane="7" entrytime="00:00:35.95" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="Kozak" nation="POL" athleteid="5380">
              <RESULTS>
                <RESULT eventid="1222" points="706" reactiontime="+88" swimtime="00:02:35.43" resultid="5381" heatid="7795" lane="2" entrytime="00:02:39.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                    <SPLIT distance="150" swimtime="00:01:54.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K16 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu" eventid="1383" reactiontime="+101" status="DSQ" swimtime="00:01:10.05" resultid="5382" heatid="7896" lane="8" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="486" reactiontime="+88" swimtime="00:00:30.13" resultid="5383" heatid="7920" lane="1" entrytime="00:00:29.99" />
                <RESULT eventid="1655" points="729" reactiontime="+90" swimtime="00:00:31.39" resultid="5384" heatid="8048" lane="8" entrytime="00:00:30.91" />
                <RESULT eventid="1703" points="526" reactiontime="+91" swimtime="00:05:02.77" resultid="5385" heatid="9061" lane="6" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:52.62" />
                    <SPLIT distance="200" swimtime="00:02:32.06" />
                    <SPLIT distance="250" swimtime="00:03:11.72" />
                    <SPLIT distance="300" swimtime="00:03:51.47" />
                    <SPLIT distance="350" swimtime="00:04:28.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="5386">
              <RESULTS>
                <RESULT eventid="1059" points="236" reactiontime="+109" swimtime="00:00:51.99" resultid="5387" heatid="7672" lane="3" entrytime="00:00:53.08" />
                <RESULT eventid="1140" points="311" swimtime="00:17:50.49" resultid="5388" heatid="8716" lane="4" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.25" />
                    <SPLIT distance="100" swimtime="00:02:08.32" />
                    <SPLIT distance="200" swimtime="00:04:25.27" />
                    <SPLIT distance="300" swimtime="00:06:41.29" />
                    <SPLIT distance="400" swimtime="00:08:56.36" />
                    <SPLIT distance="500" swimtime="00:11:10.81" />
                    <SPLIT distance="600" swimtime="00:13:25.87" />
                    <SPLIT distance="700" swimtime="00:15:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="232" reactiontime="+102" swimtime="00:01:56.20" resultid="5389" heatid="7797" lane="6" entrytime="00:02:00.69" />
                <RESULT eventid="1463" points="272" reactiontime="+93" swimtime="00:04:05.10" resultid="5390" heatid="7944" lane="6" entrytime="00:04:26.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.88" />
                    <SPLIT distance="100" swimtime="00:01:58.19" />
                    <SPLIT distance="150" swimtime="00:03:04.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="339" reactiontime="+99" swimtime="00:08:23.42" resultid="5391" heatid="9052" lane="8" entrytime="00:09:02.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.49" />
                    <SPLIT distance="100" swimtime="00:01:59.97" />
                    <SPLIT distance="150" swimtime="00:03:07.10" />
                    <SPLIT distance="200" swimtime="00:04:12.00" />
                    <SPLIT distance="250" swimtime="00:06:20.55" />
                    <SPLIT distance="300" swimtime="00:07:24.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-03-16" firstname="Ewa" gender="F" lastname="Kosmol" nation="POL" athleteid="5392">
              <RESULTS>
                <RESULT eventid="1059" points="409" reactiontime="+114" swimtime="00:00:43.43" resultid="5393" heatid="7673" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1270" points="386" reactiontime="+109" swimtime="00:01:52.45" resultid="5394" heatid="7828" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="405" reactiontime="+95" swimtime="00:03:41.62" resultid="5395" heatid="7944" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                    <SPLIT distance="100" swimtime="00:01:49.25" />
                    <SPLIT distance="150" swimtime="00:02:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="429" reactiontime="+79" swimtime="00:04:09.68" resultid="5396" heatid="8005" lane="7" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.75" />
                    <SPLIT distance="100" swimtime="00:02:02.38" />
                    <SPLIT distance="150" swimtime="00:03:07.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="5397">
              <RESULTS>
                <RESULT eventid="1254" points="631" reactiontime="+81" swimtime="00:00:59.95" resultid="5398" heatid="7819" lane="8" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="635" reactiontime="+82" swimtime="00:00:29.84" resultid="5399" heatid="7914" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1479" points="555" reactiontime="+87" swimtime="00:02:15.61" resultid="5400" heatid="7962" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:05.57" />
                    <SPLIT distance="150" swimtime="00:01:41.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="5401">
              <RESULTS>
                <RESULT eventid="1190" points="543" reactiontime="+83" swimtime="00:00:30.69" resultid="5402" heatid="7776" lane="4" entrytime="00:00:29.99" />
                <RESULT eventid="1254" points="578" reactiontime="+77" swimtime="00:00:58.31" resultid="5403" heatid="7824" lane="1" entrytime="00:00:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="5404" heatid="7965" lane="4" entrytime="00:02:11.99" />
                <RESULT eventid="1703" points="567" reactiontime="+77" swimtime="00:04:55.25" resultid="5405" heatid="9060" lane="6" entrytime="00:04:49.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:09.22" />
                    <SPLIT distance="150" swimtime="00:01:46.98" />
                    <SPLIT distance="200" swimtime="00:02:24.65" />
                    <SPLIT distance="250" swimtime="00:03:02.58" />
                    <SPLIT distance="300" swimtime="00:03:40.16" />
                    <SPLIT distance="350" swimtime="00:04:18.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka-Skorykow" nation="POL" athleteid="5406">
              <RESULTS>
                <RESULT eventid="1059" points="643" reactiontime="+77" swimtime="00:00:31.46" resultid="5407" heatid="7681" lane="2" entrytime="00:00:31.86" />
                <RESULT eventid="1206" points="638" reactiontime="+86" swimtime="00:03:08.98" resultid="5408" heatid="7782" lane="4" entrytime="00:03:14.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:29.26" />
                    <SPLIT distance="150" swimtime="00:02:18.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="596" reactiontime="+83" swimtime="00:01:20.67" resultid="5409" heatid="7833" lane="3" entrytime="00:01:23.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="622" reactiontime="+81" swimtime="00:01:26.49" resultid="5410" heatid="7879" lane="3" entrytime="00:01:28.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="600" reactiontime="+83" swimtime="00:00:35.00" resultid="5411" heatid="7902" lane="5" entrytime="00:00:35.38" />
                <RESULT eventid="1639" points="646" reactiontime="+77" swimtime="00:00:39.19" resultid="5412" heatid="8027" lane="5" entrytime="00:00:39.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="5413">
              <RESULTS>
                <RESULT eventid="1076" points="743" reactiontime="+72" swimtime="00:00:26.23" resultid="5414" heatid="7708" lane="5" entrytime="00:00:26.52" />
                <RESULT eventid="1108" points="643" reactiontime="+73" swimtime="00:02:28.11" resultid="5415" heatid="7732" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:10.53" />
                    <SPLIT distance="150" swimtime="00:01:53.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="769" reactiontime="+66" swimtime="00:00:29.63" resultid="5416" heatid="7776" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1286" points="750" reactiontime="+70" swimtime="00:01:05.82" resultid="5417" heatid="7855" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="741" reactiontime="+71" swimtime="00:00:27.76" resultid="5418" heatid="7923" lane="2" entrytime="00:00:27.90" />
                <RESULT eventid="1479" points="653" reactiontime="+75" swimtime="00:02:10.25" resultid="5419" heatid="7967" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:02.74" />
                    <SPLIT distance="150" swimtime="00:01:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="701" reactiontime="+73" swimtime="00:01:03.73" resultid="5420" heatid="8002" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="5421" entrytime="00:04:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-06-02" firstname="Wojciech" gender="M" lastname="Czupryn" nation="POL" athleteid="5422">
              <RESULTS>
                <RESULT eventid="1156" points="392" swimtime="00:26:22.45" resultid="5423" heatid="8723" lane="8" entrytime="00:28:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.41" />
                    <SPLIT distance="100" swimtime="00:01:39.24" />
                    <SPLIT distance="200" swimtime="00:03:25.33" />
                    <SPLIT distance="300" swimtime="00:03:12.05" />
                    <SPLIT distance="400" swimtime="00:06:59.08" />
                    <SPLIT distance="500" swimtime="00:08:45.53" />
                    <SPLIT distance="600" swimtime="00:10:31.81" />
                    <SPLIT distance="700" swimtime="00:12:18.04" />
                    <SPLIT distance="800" swimtime="00:14:03.17" />
                    <SPLIT distance="900" swimtime="00:15:49.34" />
                    <SPLIT distance="1000" swimtime="00:17:34.89" />
                    <SPLIT distance="1100" swimtime="00:19:20.91" />
                    <SPLIT distance="1200" swimtime="00:21:08.15" />
                    <SPLIT distance="1300" swimtime="00:22:54.63" />
                    <SPLIT distance="1400" swimtime="00:24:41.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="320" reactiontime="+85" swimtime="00:00:45.98" resultid="5424" heatid="7765" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1254" points="369" reactiontime="+87" swimtime="00:01:20.90" resultid="5425" heatid="7808" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="270" reactiontime="+86" swimtime="00:01:45.40" resultid="5426" heatid="7883" lane="6" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="277" reactiontime="+82" swimtime="00:01:45.20" resultid="5427" heatid="7934" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="326" reactiontime="+91" swimtime="00:03:45.03" resultid="5428" heatid="8012" lane="1" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.30" />
                    <SPLIT distance="100" swimtime="00:01:47.67" />
                    <SPLIT distance="150" swimtime="00:02:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="396" reactiontime="+97" swimtime="00:06:33.25" resultid="5429" heatid="9068" lane="6" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:01:32.15" />
                    <SPLIT distance="150" swimtime="00:02:21.70" />
                    <SPLIT distance="200" swimtime="00:03:12.49" />
                    <SPLIT distance="250" swimtime="00:04:03.15" />
                    <SPLIT distance="300" swimtime="00:04:53.41" />
                    <SPLIT distance="350" swimtime="00:05:44.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-18" firstname="Jacek" gender="M" lastname="Czupryn" nation="POL" athleteid="5430">
              <RESULTS>
                <RESULT eventid="1076" points="432" reactiontime="+105" swimtime="00:00:30.20" resultid="5431" heatid="7698" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1254" points="390" reactiontime="+118" swimtime="00:01:06.46" resultid="5432" heatid="7818" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="340" reactiontime="+99" swimtime="00:00:33.94" resultid="5433" heatid="7913" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1479" points="442" reactiontime="+102" swimtime="00:02:27.70" resultid="5434" heatid="7961" lane="3" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:12.71" />
                    <SPLIT distance="150" swimtime="00:01:50.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="399" reactiontime="+100" swimtime="00:05:31.97" resultid="5435" heatid="9063" lane="8" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:14.72" />
                    <SPLIT distance="150" swimtime="00:01:56.19" />
                    <SPLIT distance="200" swimtime="00:03:22.91" />
                    <SPLIT distance="250" swimtime="00:04:06.68" />
                    <SPLIT distance="300" swimtime="00:04:49.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-10-16" firstname="Rafał" gender="M" lastname="Bebelski" nation="POL" athleteid="5436">
              <RESULTS>
                <RESULT eventid="1383" points="300" reactiontime="+105" swimtime="00:01:35.63" resultid="5437" heatid="7886" lane="8" entrytime="00:01:35.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="253" reactiontime="+99" swimtime="00:02:56.12" resultid="5438" heatid="7954" lane="6" entrytime="00:03:12.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:01:23.96" />
                    <SPLIT distance="150" swimtime="00:02:10.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="299" reactiontime="+106" swimtime="00:00:43.16" resultid="5439" heatid="8033" lane="3" entrytime="00:00:44.71" />
                <RESULT eventid="1703" points="243" reactiontime="+94" swimtime="00:06:27.93" resultid="5440" heatid="9069" lane="4" entrytime="00:06:44.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                    <SPLIT distance="100" swimtime="00:01:25.43" />
                    <SPLIT distance="150" swimtime="00:02:13.36" />
                    <SPLIT distance="200" swimtime="00:03:03.55" />
                    <SPLIT distance="250" swimtime="00:03:53.77" />
                    <SPLIT distance="300" swimtime="00:04:46.06" />
                    <SPLIT distance="350" swimtime="00:05:37.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" athleteid="5441">
              <RESULTS>
                <RESULT eventid="1238" points="888" reactiontime="+72" swimtime="00:00:59.77" resultid="5442" heatid="7805" lane="4" entrytime="00:00:59.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="897" reactiontime="+72" swimtime="00:01:07.48" resultid="5443" heatid="7837" lane="5" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="947" reactiontime="+69" swimtime="00:00:29.59" resultid="5444" heatid="7905" lane="4" entrytime="00:00:29.70" />
                <RESULT eventid="1574" points="876" reactiontime="+72" swimtime="00:01:06.65" resultid="5445" heatid="7991" lane="4" entrytime="00:01:08.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-29" firstname="Jan Maciej" gender="M" lastname="Boboli" nation="POL" athleteid="6442">
              <RESULTS>
                <RESULT eventid="1076" points="432" reactiontime="+86" swimtime="00:00:37.26" resultid="6443" heatid="7690" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1190" points="156" reactiontime="+83" swimtime="00:01:01.80" resultid="6444" heatid="7765" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1254" points="346" reactiontime="+87" swimtime="00:01:30.30" resultid="6445" heatid="7808" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="476" reactiontime="+86" swimtime="00:00:39.14" resultid="6446" heatid="7910" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1655" points="93" reactiontime="+109" swimtime="00:01:17.93" resultid="6447" heatid="8031" lane="1" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="Warsaw Masters Team A" number="1">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+69" swimtime="00:01:40.77" resultid="6448" heatid="7974" lane="4" entrytime="00:01:42.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.83" />
                    <SPLIT distance="100" swimtime="00:00:50.11" />
                    <SPLIT distance="150" swimtime="00:01:15.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5356" number="1" />
                    <RELAYPOSITION athleteid="5380" number="2" />
                    <RELAYPOSITION athleteid="5401" number="3" />
                    <RELAYPOSITION athleteid="5326" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="Warsaw Masters Team A" number="2">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+92" swimtime="00:01:52.21" resultid="6449" heatid="7872" lane="4" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:01.96" />
                    <SPLIT distance="150" swimtime="00:01:27.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5401" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="5380" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="5356" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="5326" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Warsaw Masters Team B" number="6">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+97" swimtime="00:02:05.95" resultid="6453" heatid="7871" lane="3" entrytime="00:02:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:11.89" />
                    <SPLIT distance="150" swimtime="00:01:39.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5240" number="1" />
                    <RELAYPOSITION athleteid="5349" number="2" />
                    <RELAYPOSITION athleteid="5413" number="3" />
                    <RELAYPOSITION athleteid="5290" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Warsaw Masters Team B" number="8">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+84" swimtime="00:01:56.75" resultid="6455" heatid="7972" lane="4" entrytime="00:01:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:00:59.43" />
                    <SPLIT distance="150" swimtime="00:01:29.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5240" number="1" />
                    <RELAYPOSITION athleteid="5344" number="2" />
                    <RELAYPOSITION athleteid="5430" number="3" />
                    <RELAYPOSITION athleteid="5349" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Warsaw Masters Team B" number="5">
              <RESULTS>
                <RESULT eventid="1334" status="DNS" swimtime="00:00:00.00" resultid="6452" heatid="7866" lane="5" entrytime="00:02:40.90">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5334" number="1" />
                    <RELAYPOSITION athleteid="5365" number="2" />
                    <RELAYPOSITION athleteid="5233" number="3" />
                    <RELAYPOSITION athleteid="5360" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Warsaw Masters Team B" number="7">
              <RESULTS>
                <RESULT eventid="1495" reactiontime="+87" swimtime="00:02:25.94" resultid="6454" heatid="7968" lane="5" entrytime="00:02:27.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:11.61" />
                    <SPLIT distance="150" swimtime="00:01:53.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5329" number="1" />
                    <RELAYPOSITION athleteid="5306" number="2" />
                    <RELAYPOSITION athleteid="5365" number="3" />
                    <RELAYPOSITION athleteid="5334" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="Warsaw Masters Team A" number="3">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+111" swimtime="00:02:10.24" resultid="6450" heatid="7736" lane="8" entrytime="00:02:10.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:00:58.41" />
                    <SPLIT distance="150" swimtime="00:01:42.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5430" number="1" reactiontime="+111" />
                    <RELAYPOSITION athleteid="5306" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="5329" number="3" />
                    <RELAYPOSITION athleteid="5349" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Warsaw Masters Team C" number="4">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+85" swimtime="00:02:13.40" resultid="6451" heatid="7736" lane="1" entrytime="00:02:10.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:47.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5422" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="5278" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="5334" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5290" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Warsaw Masters Team C" number="9">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+58" swimtime="00:02:18.37" resultid="6456" heatid="8051" lane="2" entrytime="00:02:17.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:01:52.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5375" number="1" reactiontime="+58" />
                    <RELAYPOSITION athleteid="5369" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="5406" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5290" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WKZAB" nation="POL" region="06" clubid="6376" name="Water Knights Zabierzów">
          <ATHLETES>
            <ATHLETE birthdate="1972-01-15" firstname="Grzegorz" gender="M" lastname="Mytnik" nation="POL" athleteid="6377">
              <RESULTS>
                <RESULT eventid="1156" points="396" swimtime="00:22:37.09" resultid="6378" heatid="8720" lane="5" entrytime="00:22:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:21.55" />
                    <SPLIT distance="200" swimtime="00:02:49.44" />
                    <SPLIT distance="300" swimtime="00:04:17.70" />
                    <SPLIT distance="400" swimtime="00:05:48.39" />
                    <SPLIT distance="500" swimtime="00:07:19.21" />
                    <SPLIT distance="600" swimtime="00:08:50.89" />
                    <SPLIT distance="700" swimtime="00:10:22.75" />
                    <SPLIT distance="800" swimtime="00:11:55.59" />
                    <SPLIT distance="900" swimtime="00:13:27.77" />
                    <SPLIT distance="1000" swimtime="00:15:00.74" />
                    <SPLIT distance="1100" swimtime="00:16:32.72" />
                    <SPLIT distance="1200" swimtime="00:18:04.90" />
                    <SPLIT distance="1300" swimtime="00:19:37.62" />
                    <SPLIT distance="1400" swimtime="00:21:09.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="376" reactiontime="+98" swimtime="00:05:33.26" resultid="6379" heatid="9065" lane="2" entrytime="00:05:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:18.26" />
                    <SPLIT distance="150" swimtime="00:02:00.83" />
                    <SPLIT distance="200" swimtime="00:02:43.72" />
                    <SPLIT distance="250" swimtime="00:03:26.60" />
                    <SPLIT distance="300" swimtime="00:04:09.33" />
                    <SPLIT distance="350" swimtime="00:04:52.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="375" reactiontime="+93" swimtime="00:02:36.65" resultid="6380" heatid="7958" lane="6" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:16.21" />
                    <SPLIT distance="150" swimtime="00:01:56.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="YMKRA" nation="POL" region="06" clubid="6283" name="YMCA Kraków">
          <ATHLETES>
            <ATHLETE birthdate="1957-03-25" firstname="Jacek" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="6282">
              <RESULTS>
                <RESULT eventid="1076" points="552" reactiontime="+75" swimtime="00:00:31.78" resultid="6284" heatid="7694" lane="4" entrytime="00:00:31.25" />
                <RESULT eventid="1156" points="457" swimtime="00:25:03.85" resultid="6285" heatid="8721" lane="8" entrytime="00:24:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                    <SPLIT distance="100" swimtime="00:01:24.30" />
                    <SPLIT distance="200" swimtime="00:02:59.85" />
                    <SPLIT distance="300" swimtime="00:04:40.30" />
                    <SPLIT distance="400" swimtime="00:06:21.62" />
                    <SPLIT distance="500" swimtime="00:08:03.38" />
                    <SPLIT distance="600" swimtime="00:09:45.70" />
                    <SPLIT distance="700" swimtime="00:11:27.52" />
                    <SPLIT distance="800" swimtime="00:13:09.85" />
                    <SPLIT distance="900" swimtime="00:14:50.98" />
                    <SPLIT distance="1000" swimtime="00:16:34.12" />
                    <SPLIT distance="1100" swimtime="00:18:18.17" />
                    <SPLIT distance="1200" swimtime="00:20:00.67" />
                    <SPLIT distance="1300" swimtime="00:22:35.97" />
                    <SPLIT distance="1400" swimtime="00:24:15.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="530" reactiontime="+79" swimtime="00:01:11.67" resultid="6286" heatid="7813" lane="1" entrytime="00:01:11.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="6287" heatid="7911" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1479" points="521" reactiontime="+77" swimtime="00:02:45.63" resultid="6288" heatid="7957" lane="2" entrytime="00:02:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:02.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="532" reactiontime="+73" swimtime="00:05:56.61" resultid="6289" heatid="9066" lane="6" entrytime="00:05:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:01:18.95" />
                    <SPLIT distance="150" swimtime="00:02:03.89" />
                    <SPLIT distance="250" swimtime="00:03:37.49" />
                    <SPLIT distance="300" swimtime="00:04:24.04" />
                    <SPLIT distance="350" swimtime="00:05:11.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="INDYW" nation="POL" clubid="1892" name="Zawodnik niezrzeszony">
          <CONTACT email="piotr_urbanczyk@onet.pl" name="URBAŃCZYK PIOTR" phone="608172201" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-02" firstname="Janusz" gender="M" lastname="Płonka" nation="POL" athleteid="1893">
              <RESULTS>
                <RESULT eventid="1415" points="237" reactiontime="+103" swimtime="00:00:49.38" resultid="1894" heatid="7907" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1318" points="166" reactiontime="+100" swimtime="00:05:03.98" resultid="1895" heatid="7859" lane="6" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.65" />
                    <SPLIT distance="100" swimtime="00:02:21.93" />
                    <SPLIT distance="150" swimtime="00:03:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="179" reactiontime="+104" swimtime="00:02:07.01" resultid="1896" heatid="7992" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="189" reactiontime="+107" swimtime="00:01:01.52" resultid="1897" heatid="8030" lane="4" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-06" firstname="Arkadiusz" gender="M" lastname="Doliński" nation="POL" athleteid="1911">
              <RESULTS>
                <RESULT eventid="1076" points="566" reactiontime="+85" swimtime="00:00:28.66" resultid="1912" heatid="7687" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1108" points="361" reactiontime="+97" swimtime="00:02:58.69" resultid="1913" heatid="7724" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:21.32" />
                    <SPLIT distance="150" swimtime="00:02:14.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="570" reactiontime="+69" swimtime="00:00:32.72" resultid="1914" heatid="7769" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1286" points="489" reactiontime="+94" swimtime="00:01:14.95" resultid="1915" heatid="7842" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="533" reactiontime="+74" swimtime="00:01:12.90" resultid="1916" heatid="7936" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="1917" heatid="8810" lane="5" entrytime="00:07:00.00" />
                <RESULT eventid="1623" points="439" reactiontime="+78" swimtime="00:02:50.96" resultid="1918" heatid="8014" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:24.24" />
                    <SPLIT distance="150" swimtime="00:02:08.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-06-05" firstname="Marek" gender="M" lastname="Żuber" nation="POL" athleteid="1925">
              <RESULTS>
                <RESULT eventid="1076" points="618" reactiontime="+82" swimtime="00:00:27.84" resultid="1926" heatid="7706" lane="4" entrytime="00:00:27.20" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="1927" heatid="7820" lane="1" entrytime="00:01:02.00" />
                <RESULT eventid="1415" points="626" reactiontime="+77" swimtime="00:00:29.99" resultid="1928" heatid="7921" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="1929" heatid="8001" lane="3" entrytime="00:01:07.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-11-19" firstname="Judyta" gender="F" lastname="Sołtyk" nation="POL" athleteid="1939">
              <RESULTS>
                <RESULT eventid="1092" points="645" reactiontime="+83" swimtime="00:02:48.05" resultid="1940" heatid="7717" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:08.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="629" reactiontime="+86" swimtime="00:02:29.52" resultid="1941" heatid="7950" lane="7" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:11.46" />
                    <SPLIT distance="150" swimtime="00:01:50.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="667" reactiontime="+88" swimtime="00:06:01.10" resultid="1943" heatid="8803" lane="5" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="150" swimtime="00:02:05.72" />
                    <SPLIT distance="200" swimtime="00:02:52.00" />
                    <SPLIT distance="250" swimtime="00:03:44.24" />
                    <SPLIT distance="300" swimtime="00:04:37.93" />
                    <SPLIT distance="350" swimtime="00:05:20.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-05" firstname="Michał" gender="M" lastname="Wągrowski" nation="POL" athleteid="1944">
              <RESULTS>
                <RESULT eventid="1076" points="633" reactiontime="+82" swimtime="00:00:27.62" resultid="1945" heatid="7709" lane="6" entrytime="00:00:26.30" />
                <RESULT comment="G7 - Brak pozycji na plecach przy opuszczaniu ściany nawrotowej  (Czas: 18:23)" eventid="1108" reactiontime="+90" status="DSQ" swimtime="00:02:58.87" resultid="1946" heatid="7731" lane="1" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:21.86" />
                    <SPLIT distance="150" swimtime="00:02:16.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="526" reactiontime="+85" swimtime="00:01:03.70" resultid="1947" heatid="7821" lane="7" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="439" reactiontime="+88" swimtime="00:01:17.68" resultid="1948" heatid="7848" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="402" reactiontime="+85" swimtime="00:00:34.75" resultid="1949" heatid="7918" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1479" points="381" reactiontime="+86" swimtime="00:02:33.63" resultid="1950" heatid="7962" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                    <SPLIT distance="100" swimtime="00:01:07.21" />
                    <SPLIT distance="150" swimtime="00:01:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="372" reactiontime="+91" swimtime="00:00:40.13" resultid="1951" heatid="8039" lane="2" entrytime="00:00:38.50" />
                <RESULT eventid="1703" points="359" reactiontime="+87" swimtime="00:05:40.87" resultid="1952" heatid="9063" lane="6" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:10.65" />
                    <SPLIT distance="150" swimtime="00:01:52.13" />
                    <SPLIT distance="200" swimtime="00:03:22.86" />
                    <SPLIT distance="250" swimtime="00:04:09.33" />
                    <SPLIT distance="300" swimtime="00:04:56.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-03-11" firstname="Kazimierz" gender="M" lastname="From" nation="POL" athleteid="1953">
              <RESULTS>
                <RESULT eventid="1076" points="186" reactiontime="+124" swimtime="00:00:58.12" resultid="1954" heatid="7684" lane="4" entrytime="00:00:57.00" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="1955" heatid="8725" lane="4" entrytime="00:45:00.00" />
                <RESULT eventid="1190" points="179" reactiontime="+92" swimtime="00:01:17.52" resultid="1956" heatid="7763" lane="7" entrytime="00:01:15.00" />
                <RESULT eventid="1254" points="171" reactiontime="+129" swimtime="00:02:21.65" resultid="1957" heatid="7806" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="163" reactiontime="+99" swimtime="00:02:55.79" resultid="1958" heatid="7932" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="190" reactiontime="+122" swimtime="00:05:13.30" resultid="1959" heatid="7952" lane="5" entrytime="00:05:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.44" />
                    <SPLIT distance="100" swimtime="00:02:25.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="155" reactiontime="+103" swimtime="00:06:30.66" resultid="1960" heatid="8010" lane="7" entrytime="00:06:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.32" />
                    <SPLIT distance="100" swimtime="00:03:05.44" />
                    <SPLIT distance="150" swimtime="00:04:49.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="1961" entrytime="00:11:22.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-09" firstname="Paulina" gender="F" lastname="Szymańska" nation="POL" athleteid="1962">
              <RESULTS>
                <RESULT eventid="1206" points="464" reactiontime="+74" swimtime="00:03:18.46" resultid="1963" heatid="7782" lane="7" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                    <SPLIT distance="100" swimtime="00:01:35.71" />
                    <SPLIT distance="150" swimtime="00:02:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="347" reactiontime="+76" swimtime="00:01:33.02" resultid="1964" heatid="7831" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="421" reactiontime="+75" swimtime="00:01:34.21" resultid="1965" heatid="7878" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-04-01" firstname="Dariusz" gender="M" lastname="Krause" nation="POL" athleteid="1975">
              <RESULTS>
                <RESULT eventid="1076" points="468" reactiontime="+79" swimtime="00:00:30.60" resultid="1976" heatid="7698" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1254" points="410" reactiontime="+84" swimtime="00:01:10.07" resultid="1977" heatid="7813" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="1978">
              <RESULTS>
                <RESULT eventid="1238" points="579" reactiontime="+106" swimtime="00:01:22.18" resultid="1980" heatid="7799" lane="4" entrytime="00:01:26.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="699" reactiontime="+100" swimtime="00:01:29.86" resultid="1981" heatid="7928" lane="7" entrytime="00:01:33.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="774" reactiontime="+91" swimtime="00:03:07.53" resultid="1982" heatid="8007" lane="2" entrytime="00:03:13.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                    <SPLIT distance="100" swimtime="00:01:32.48" />
                    <SPLIT distance="150" swimtime="00:02:20.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-09-19" firstname="Wiesław" gender="M" lastname="Majcher" nation="POL" athleteid="1983">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="1984" heatid="7689" lane="7" entrytime="00:00:35.42" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="1985" heatid="8724" lane="7" entrytime="00:31:51.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-02-20" firstname="Zofia" gender="F" lastname="Brunka" nation="POL" athleteid="1986">
              <RESULTS>
                <RESULT eventid="1173" points="475" reactiontime="+69" swimtime="00:00:38.81" resultid="1987" heatid="7759" lane="8" entrytime="00:00:38.37" />
                <RESULT eventid="1270" points="397" reactiontime="+86" swimtime="00:01:28.52" resultid="1988" heatid="7833" lane="5" entrytime="00:01:23.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="442" swimtime="00:01:25.59" resultid="1989" heatid="7929" lane="4" entrytime="00:01:24.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="474" reactiontime="+43" swimtime="00:03:04.48" resultid="1990" heatid="8008" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                    <SPLIT distance="150" swimtime="00:02:16.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-03" firstname="Piotr" gender="M" lastname="Fuliński" nation="POL" athleteid="1991">
              <RESULTS>
                <RESULT eventid="1076" points="589" reactiontime="+91" swimtime="00:00:26.39" resultid="1992" heatid="7710" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1254" points="546" reactiontime="+92" swimtime="00:01:00.00" resultid="1993" heatid="7823" lane="6" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="1994" heatid="7965" lane="6" entrytime="00:02:14.00" />
                <RESULT eventid="1703" status="DNS" swimtime="00:00:00.00" resultid="1995" heatid="9061" lane="7" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-08" firstname="Stanisław" gender="M" lastname="Filipek" nation="POL" athleteid="1996">
              <RESULTS>
                <RESULT eventid="1222" points="328" reactiontime="+104" swimtime="00:04:28.40" resultid="1997" heatid="7784" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.14" />
                    <SPLIT distance="100" swimtime="00:02:07.63" />
                    <SPLIT distance="150" swimtime="00:03:19.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="308" reactiontime="+104" swimtime="00:02:03.82" resultid="1998" heatid="7881" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="362" reactiontime="+104" swimtime="00:00:52.52" resultid="1999" heatid="8029" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-12-24" firstname="Aleksandra" gender="F" lastname="Zackiewicz" nation="POL" athleteid="2000">
              <RESULTS>
                <RESULT eventid="1173" status="DNS" swimtime="00:00:00.00" resultid="2001" heatid="7761" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1270" status="DNS" swimtime="00:00:00.00" resultid="2002" heatid="7837" lane="4" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-05-04" firstname="Krzysztof" gender="M" lastname="Wiater " nation="POL" athleteid="2003">
              <RESULTS>
                <RESULT eventid="1156" points="404" swimtime="00:22:28.03" resultid="2004" heatid="8725" lane="2" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:17.09" />
                    <SPLIT distance="200" swimtime="00:02:42.77" />
                    <SPLIT distance="300" swimtime="00:04:10.17" />
                    <SPLIT distance="400" swimtime="00:05:40.18" />
                    <SPLIT distance="500" swimtime="00:07:11.09" />
                    <SPLIT distance="600" swimtime="00:08:41.78" />
                    <SPLIT distance="700" swimtime="00:10:13.36" />
                    <SPLIT distance="800" swimtime="00:11:43.92" />
                    <SPLIT distance="900" swimtime="00:13:15.63" />
                    <SPLIT distance="1000" swimtime="00:14:47.64" />
                    <SPLIT distance="1100" swimtime="00:16:20.30" />
                    <SPLIT distance="1200" swimtime="00:17:53.11" />
                    <SPLIT distance="1300" swimtime="00:19:25.65" />
                    <SPLIT distance="1400" swimtime="00:20:58.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Andrzej" gender="M" lastname="Fajdasz" nation="POL" athleteid="2113">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2114" heatid="7702" lane="7" entrytime="00:00:28.65" />
                <RESULT eventid="1254" points="493" reactiontime="+75" swimtime="00:01:05.91" resultid="2115" heatid="7814" lane="7" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="472" reactiontime="+79" swimtime="00:01:16.82" resultid="2116" heatid="7846" lane="5" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="379" reactiontime="+83" swimtime="00:00:34.71" resultid="2117" heatid="7910" lane="6" entrytime="00:00:38.25" />
                <RESULT eventid="1447" points="423" reactiontime="+75" swimtime="00:01:18.65" resultid="2118" heatid="7938" lane="2" entrytime="00:01:19.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="417" reactiontime="+80" status="EXH" swimtime="00:00:39.47" resultid="9040" heatid="8029" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-11-22" firstname="Marek" gender="M" lastname="Pałysa" nation="POL" athleteid="2199">
              <RESULTS>
                <RESULT eventid="1254" points="454" reactiontime="+80" swimtime="00:01:06.91" resultid="2200" heatid="7816" lane="2" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="459" reactiontime="+84" swimtime="00:01:16.51" resultid="2201" heatid="7845" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="450" reactiontime="+78" swimtime="00:01:23.50" resultid="2202" heatid="7888" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)  (Czas: 11:38)" eventid="1655" reactiontime="+68" status="DSQ" swimtime="00:00:35.75" resultid="2203" heatid="8044" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-16" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="2541">
              <RESULTS>
                <RESULT eventid="1076" points="805" reactiontime="+77" swimtime="00:00:27.31" resultid="2542" heatid="7705" lane="8" entrytime="00:00:27.85" />
                <RESULT eventid="1108" points="792" reactiontime="+81" swimtime="00:02:34.46" resultid="2543" heatid="7730" lane="1" entrytime="00:02:37.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:56.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="797" reactiontime="+82" swimtime="00:01:00.87" resultid="2544" heatid="7820" lane="5" entrytime="00:01:01.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="835" reactiontime="+81" swimtime="00:01:09.52" resultid="2545" heatid="7852" lane="6" entrytime="00:01:09.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="776" reactiontime="+79" swimtime="00:00:29.98" resultid="2546" heatid="7919" lane="1" entrytime="00:00:30.35" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="2547" heatid="7963" lane="4" entrytime="00:02:18.75" />
                <RESULT eventid="1591" points="751" reactiontime="+82" swimtime="00:01:08.70" resultid="2548" heatid="8000" lane="3" entrytime="00:01:09.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="743" reactiontime="+78" swimtime="00:02:40.06" resultid="2549" heatid="8016" lane="5" entrytime="00:02:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                    <SPLIT distance="150" swimtime="00:01:59.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-02-17" firstname="Piotr" gender="M" lastname="Kister" nation="POL" athleteid="2559">
              <RESULTS>
                <RESULT eventid="1222" points="486" reactiontime="+82" swimtime="00:02:57.43" resultid="2560" heatid="7794" lane="8" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:09.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="395" reactiontime="+80" swimtime="00:02:50.13" resultid="2561" heatid="7864" lane="6" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:02:00.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="445" reactiontime="+85" swimtime="00:01:20.85" resultid="2562" heatid="7892" lane="7" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="511" reactiontime="+84" swimtime="00:00:31.24" resultid="2563" heatid="7916" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="1591" points="473" reactiontime="+83" swimtime="00:01:10.72" resultid="2564" heatid="7999" lane="5" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="513" reactiontime="+81" swimtime="00:00:35.30" resultid="2565" heatid="8043" lane="5" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Anna" gender="F" lastname="Kotusińska" nation="POL" athleteid="2569">
              <RESULTS>
                <RESULT eventid="1238" points="372" reactiontime="+92" swimtime="00:01:21.14" resultid="2584" heatid="7801" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="364" reactiontime="+83" swimtime="00:00:40.70" resultid="2585" heatid="7900" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="2576">
              <RESULTS>
                <RESULT eventid="1076" points="739" reactiontime="+72" swimtime="00:00:25.43" resultid="2577" heatid="7711" lane="3" entrytime="00:00:25.50" />
                <RESULT eventid="1108" points="660" reactiontime="+73" swimtime="00:02:25.84" resultid="2578" heatid="7731" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="150" swimtime="00:01:50.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="759" reactiontime="+75" swimtime="00:00:55.81" resultid="2579" heatid="7824" lane="6" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="673" reactiontime="+80" swimtime="00:01:05.52" resultid="2580" heatid="7855" lane="4" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="802" reactiontime="+71" swimtime="00:00:26.89" resultid="2581" heatid="7924" lane="6" entrytime="00:00:27.05" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="2582" heatid="8807" lane="8" entrytime="00:06:00.00" />
                <RESULT eventid="1591" points="702" reactiontime="+76" swimtime="00:01:02.01" resultid="2583" heatid="8002" lane="3" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-02" firstname="Tomasz" gender="M" lastname="Jąkalski" nation="POL" athleteid="2586">
              <RESULTS>
                <RESULT eventid="1190" points="609" reactiontime="+62" swimtime="00:00:29.54" resultid="2587" heatid="7776" lane="1" entrytime="00:00:30.01" />
                <RESULT eventid="1286" points="561" reactiontime="+88" swimtime="00:01:06.90" resultid="2588" heatid="7854" lane="7" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="587" reactiontime="+69" swimtime="00:01:05.70" resultid="2589" heatid="7941" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="2590" heatid="8808" lane="1" entrytime="00:06:15.00" />
                <RESULT eventid="1623" points="474" reactiontime="+72" swimtime="00:02:29.04" resultid="2591" heatid="8018" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="150" swimtime="00:01:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="555" reactiontime="+86" swimtime="00:00:34.37" resultid="2592" heatid="8045" lane="5" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-06-05" firstname="Lukas" gender="M" lastname="Smiesko" nation="POL" athleteid="2593">
              <RESULTS>
                <RESULT eventid="1286" points="786" reactiontime="+78" swimtime="00:01:02.22" resultid="2594" heatid="7856" lane="6" entrytime="00:01:02.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="841" reactiontime="+80" swimtime="00:00:26.47" resultid="2595" heatid="7925" lane="2" entrytime="00:00:26.39" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Olga" gender="F" lastname="Krysiak" nation="POL" athleteid="2605">
              <RESULTS>
                <RESULT eventid="1059" points="779" reactiontime="+83" swimtime="00:00:28.77" resultid="2606" heatid="7683" lane="7" entrytime="00:00:29.11" />
                <RESULT eventid="1238" points="764" reactiontime="+75" swimtime="00:01:03.30" resultid="2607" heatid="7805" lane="2" entrytime="00:01:03.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="584" reactiontime="+81" swimtime="00:01:17.89" resultid="2608" heatid="7836" lane="8" entrytime="00:01:17.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="645" reactiontime="+79" swimtime="00:02:22.48" resultid="2609" heatid="7951" lane="2" entrytime="00:02:23.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:07.74" />
                    <SPLIT distance="150" swimtime="00:01:45.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="560" reactiontime="+78" swimtime="00:05:13.71" resultid="2610" heatid="9047" lane="8" entrytime="00:05:14.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:12.81" />
                    <SPLIT distance="150" swimtime="00:01:52.65" />
                    <SPLIT distance="200" swimtime="00:02:33.14" />
                    <SPLIT distance="250" swimtime="00:03:14.34" />
                    <SPLIT distance="300" swimtime="00:03:54.77" />
                    <SPLIT distance="350" swimtime="00:04:34.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-01" firstname="Katarzyna" gender="F" lastname="Koba" nation="POL" athleteid="2646">
              <RESULTS>
                <RESULT eventid="1059" points="576" reactiontime="+89" swimtime="00:00:31.87" resultid="2647" heatid="7679" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1399" points="451" reactiontime="+91" swimtime="00:00:37.89" resultid="2648" heatid="7902" lane="8" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="2649">
              <RESULTS>
                <RESULT eventid="1076" points="563" reactiontime="+96" swimtime="00:00:32.68" resultid="2650" heatid="7693" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1156" points="642" swimtime="00:24:46.75" resultid="2651" heatid="8723" lane="7" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                    <SPLIT distance="100" swimtime="00:01:31.65" />
                    <SPLIT distance="200" swimtime="00:03:10.07" />
                    <SPLIT distance="300" swimtime="00:04:47.22" />
                    <SPLIT distance="400" swimtime="00:06:27.56" />
                    <SPLIT distance="500" swimtime="00:08:06.95" />
                    <SPLIT distance="600" swimtime="00:09:48.69" />
                    <SPLIT distance="700" swimtime="00:11:30.04" />
                    <SPLIT distance="800" swimtime="00:13:12.04" />
                    <SPLIT distance="900" swimtime="00:14:52.47" />
                    <SPLIT distance="1000" swimtime="00:16:32.81" />
                    <SPLIT distance="1100" swimtime="00:18:13.04" />
                    <SPLIT distance="1200" swimtime="00:19:53.53" />
                    <SPLIT distance="1300" swimtime="00:21:35.15" />
                    <SPLIT distance="1400" swimtime="00:23:13.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="603" reactiontime="+77" swimtime="00:00:39.22" resultid="2652" heatid="7770" lane="7" entrytime="00:00:39.01" />
                <RESULT eventid="1318" points="346" reactiontime="+107" swimtime="00:03:47.46" resultid="2653" heatid="7861" lane="5" entrytime="00:03:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.33" />
                    <SPLIT distance="100" swimtime="00:01:44.44" />
                    <SPLIT distance="150" swimtime="00:02:44.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="568" reactiontime="+84" swimtime="00:01:27.77" resultid="2654" heatid="7936" lane="3" entrytime="00:01:29.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="523" reactiontime="+92" swimtime="00:07:12.73" resultid="2655" heatid="8810" lane="8" entrytime="00:07:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.38" />
                    <SPLIT distance="100" swimtime="00:01:48.04" />
                    <SPLIT distance="150" swimtime="00:02:42.62" />
                    <SPLIT distance="200" swimtime="00:04:44.56" />
                    <SPLIT distance="250" swimtime="00:05:47.03" />
                    <SPLIT distance="300" swimtime="00:06:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="574" reactiontime="+102" swimtime="00:03:19.08" resultid="2656" heatid="8013" lane="8" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                    <SPLIT distance="100" swimtime="00:01:40.10" />
                    <SPLIT distance="150" swimtime="00:02:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" points="513" reactiontime="+97" swimtime="00:06:15.75" resultid="2657" heatid="9068" lane="5" entrytime="00:06:29.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="100" swimtime="00:01:22.34" />
                    <SPLIT distance="150" swimtime="00:02:08.99" />
                    <SPLIT distance="200" swimtime="00:02:56.43" />
                    <SPLIT distance="250" swimtime="00:03:45.34" />
                    <SPLIT distance="300" swimtime="00:04:35.46" />
                    <SPLIT distance="350" swimtime="00:05:25.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-04-24" firstname="Włodzimierz" gender="M" lastname="Zieleziński" nation="POL" athleteid="2667">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2668" heatid="7689" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1156" points="522" swimtime="00:26:32.72" resultid="2669" heatid="8724" lane="4" entrytime="00:28:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                    <SPLIT distance="100" swimtime="00:01:30.17" />
                    <SPLIT distance="200" swimtime="00:03:12.79" />
                    <SPLIT distance="300" swimtime="00:04:58.31" />
                    <SPLIT distance="400" swimtime="00:06:45.50" />
                    <SPLIT distance="500" swimtime="00:08:33.15" />
                    <SPLIT distance="600" swimtime="00:10:21.79" />
                    <SPLIT distance="700" swimtime="00:12:09.92" />
                    <SPLIT distance="800" swimtime="00:13:58.47" />
                    <SPLIT distance="900" swimtime="00:15:48.83" />
                    <SPLIT distance="1000" swimtime="00:17:37.38" />
                    <SPLIT distance="1100" swimtime="00:19:27.14" />
                    <SPLIT distance="1200" swimtime="00:21:15.93" />
                    <SPLIT distance="1300" swimtime="00:23:03.43" />
                    <SPLIT distance="1400" swimtime="00:24:50.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="460" reactiontime="+88" swimtime="00:00:42.94" resultid="2670" heatid="7768" lane="4" entrytime="00:00:41.50" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="2671" heatid="7810" lane="4" entrytime="00:01:17.00" />
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="2672" heatid="7934" lane="4" entrytime="00:01:45.00" />
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="2673" heatid="7955" lane="7" entrytime="00:03:05.00" />
                <RESULT eventid="1703" points="486" reactiontime="+112" swimtime="00:06:22.43" resultid="2674" heatid="9068" lane="2" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:26.93" />
                    <SPLIT distance="150" swimtime="00:02:17.19" />
                    <SPLIT distance="200" swimtime="00:03:07.79" />
                    <SPLIT distance="250" swimtime="00:03:58.51" />
                    <SPLIT distance="300" swimtime="00:04:48.03" />
                    <SPLIT distance="350" swimtime="00:05:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="2767" heatid="8012" lane="7" entrytime="00:03:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Tomasz" gender="M" lastname="Jaroń" nation="POL" athleteid="2726">
              <RESULTS>
                <RESULT eventid="1108" points="356" reactiontime="+72" swimtime="00:03:00.40" resultid="2727" heatid="7726" lane="6" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:28.65" />
                    <SPLIT distance="150" swimtime="00:02:19.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="444" reactiontime="+76" swimtime="00:03:07.23" resultid="2729" heatid="7792" lane="3" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                    <SPLIT distance="100" swimtime="00:01:29.40" />
                    <SPLIT distance="150" swimtime="00:02:18.60" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M11 - Brak dotknięcia ściany obydwoma rozłączonymi dłońmi przy nawrocie lub na zakończenie wyścigu  (Czas: 13:58)" eventid="1318" reactiontime="+72" status="DSQ" swimtime="00:03:21.79" resultid="2730" heatid="7862" lane="3" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:31.49" />
                    <SPLIT distance="150" swimtime="00:02:26.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="400" reactiontime="+70" swimtime="00:01:29.02" resultid="2731" heatid="7889" lane="3" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="326" reactiontime="+78" swimtime="00:06:33.74" resultid="2732" heatid="8809" lane="3" entrytime="00:06:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:29.50" />
                    <SPLIT distance="150" swimtime="00:02:24.40" />
                    <SPLIT distance="200" swimtime="00:03:18.15" />
                    <SPLIT distance="250" swimtime="00:04:10.91" />
                    <SPLIT distance="300" swimtime="00:05:04.11" />
                    <SPLIT distance="350" swimtime="00:05:49.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="2733" heatid="7996" lane="5" entrytime="00:01:22.00" />
                <RESULT eventid="1655" points="386" reactiontime="+70" swimtime="00:00:40.48" resultid="2734" heatid="8038" lane="6" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-06-28" firstname="Bolesław" gender="M" lastname="Czyż" nation="POL" athleteid="2735">
              <RESULTS>
                <RESULT eventid="1108" points="359" reactiontime="+108" swimtime="00:03:47.36" resultid="2736" heatid="7721" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.69" />
                    <SPLIT distance="100" swimtime="00:01:54.75" />
                    <SPLIT distance="150" swimtime="00:02:55.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="328" reactiontime="+104" swimtime="00:04:02.54" resultid="2737" heatid="7861" lane="7" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.40" />
                    <SPLIT distance="100" swimtime="00:01:56.05" />
                    <SPLIT distance="150" swimtime="00:02:59.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="2738" heatid="7884" lane="8" entrytime="00:01:43.00" />
                <RESULT comment="K4 - Cykl ruchowy inny niż jeden ruch ramion i jedno kopnięcie nogami  (Czas: 22:08)" eventid="1543" reactiontime="+107" status="DSQ" swimtime="00:08:17.38" resultid="2739" heatid="8811" lane="2" entrytime="00:08:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.96" />
                    <SPLIT distance="100" swimtime="00:01:57.57" />
                    <SPLIT distance="150" swimtime="00:03:06.54" />
                    <SPLIT distance="200" swimtime="00:04:16.99" />
                    <SPLIT distance="250" swimtime="00:05:20.50" />
                    <SPLIT distance="300" swimtime="00:06:25.21" />
                    <SPLIT distance="350" swimtime="00:07:22.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="287" reactiontime="+109" swimtime="00:01:48.55" resultid="2740" heatid="7996" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="2741" heatid="8033" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-04" firstname="Marek" gender="M" lastname="Pogorzelski" nation="POL" athleteid="3090">
              <RESULTS>
                <RESULT eventid="1076" points="483" reactiontime="+89" swimtime="00:00:30.81" resultid="3091" heatid="7695" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1108" points="398" reactiontime="+86" swimtime="00:03:05.64" resultid="3092" heatid="7725" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:27.96" />
                    <SPLIT distance="150" swimtime="00:02:23.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="444" reactiontime="+83" swimtime="00:01:09.33" resultid="3093" heatid="7812" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="406" reactiontime="+84" swimtime="00:01:21.63" resultid="3094" heatid="7845" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="411" reactiontime="+92" swimtime="00:01:30.37" resultid="3095" heatid="7884" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="359" reactiontime="+88" swimtime="00:00:37.18" resultid="3096" heatid="7910" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="3097" heatid="7994" lane="5" entrytime="00:01:40.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="3098" heatid="8038" lane="8" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-23" firstname="Artur" gender="M" lastname="Włoszek" nation="POL" athleteid="3516">
              <RESULTS>
                <RESULT eventid="1076" points="585" reactiontime="+67" swimtime="00:00:26.46" resultid="3517" heatid="7698" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1108" points="407" reactiontime="+71" swimtime="00:02:39.33" resultid="3518" heatid="7724" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:02:00.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-23" firstname="Andrzej" gender="M" lastname="Matiolański" nation="POL" athleteid="3519">
              <RESULTS>
                <RESULT eventid="1286" points="433" reactiontime="+92" swimtime="00:01:12.93" resultid="3520" heatid="7847" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="518" reactiontime="+91" swimtime="00:00:29.51" resultid="3521" heatid="7921" lane="8" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-08" firstname="Kamil" gender="M" lastname="Chylak" nation="POL" athleteid="3522">
              <RESULTS>
                <RESULT eventid="1076" points="258" reactiontime="+94" swimtime="00:00:34.75" resultid="3523" heatid="7689" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1703" points="202" reactiontime="+95" swimtime="00:06:49.26" resultid="3524" heatid="9069" lane="5" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:23.63" />
                    <SPLIT distance="150" swimtime="00:02:15.08" />
                    <SPLIT distance="200" swimtime="00:03:09.27" />
                    <SPLIT distance="250" swimtime="00:04:04.21" />
                    <SPLIT distance="300" swimtime="00:04:59.56" />
                    <SPLIT distance="350" swimtime="00:05:54.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Bartłomiej" gender="M" lastname="Jankowski" nation="POL" athleteid="3531">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="3532" heatid="7731" lane="4" entrytime="00:02:29.00" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="3533" heatid="7794" lane="3" entrytime="00:02:46.00" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="3534" heatid="7864" lane="1" entrytime="00:02:50.00" />
                <RESULT eventid="1383" status="DNS" swimtime="00:00:00.00" resultid="3535" heatid="7895" lane="2" entrytime="00:01:11.00" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="3536" heatid="7921" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="3537" heatid="8017" lane="5" entrytime="00:02:40.00" />
                <RESULT eventid="1655" status="DNS" swimtime="00:00:00.00" resultid="3538" heatid="8045" lane="2" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-02-11" firstname="Agnieszka" gender="F" lastname="Figuła" nation="POL" athleteid="3539">
              <RESULTS>
                <RESULT eventid="1059" points="595" reactiontime="+79" swimtime="00:00:31.52" resultid="3540" heatid="7681" lane="3" entrytime="00:00:31.16" />
                <RESULT eventid="1238" points="630" reactiontime="+77" swimtime="00:01:08.09" resultid="3541" heatid="7803" lane="4" entrytime="00:01:08.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="566" reactiontime="+81" swimtime="00:01:25.39" resultid="3542" heatid="7880" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="614" reactiontime="+83" swimtime="00:00:34.20" resultid="3543" heatid="7902" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1639" points="526" reactiontime="+80" swimtime="00:00:39.12" resultid="3544" heatid="8028" lane="7" entrytime="00:00:38.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-03" firstname="Patryk" gender="M" lastname="Dzwonek" nation="POL" athleteid="3545">
              <RESULTS>
                <RESULT eventid="1076" points="607" reactiontime="+81" swimtime="00:00:28.06" resultid="3546" heatid="7704" lane="3" entrytime="00:00:28.00" />
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1479" reactiontime="+54" status="DSQ" swimtime="00:02:29.60" resultid="3547" heatid="7959" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:06.73" />
                    <SPLIT distance="150" swimtime="00:01:48.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-08-03" firstname="Daniel" gender="M" lastname="Waliszewski" nation="POL" athleteid="3548">
              <RESULTS>
                <RESULT eventid="1383" points="716" reactiontime="+81" swimtime="00:01:09.03" resultid="3549" heatid="7896" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-11-29" firstname="Edward" gender="M" lastname="Dziekoński" nation="POL" athleteid="3550">
              <RESULTS>
                <RESULT eventid="1076" points="355" reactiontime="+100" swimtime="00:00:40.92" resultid="3551" heatid="7686" lane="1" entrytime="00:00:41.20" />
                <RESULT eventid="1156" points="522" swimtime="00:28:40.47" resultid="3552" heatid="8724" lane="3" entrytime="00:29:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.16" />
                    <SPLIT distance="100" swimtime="00:01:46.23" />
                    <SPLIT distance="200" swimtime="00:03:41.22" />
                    <SPLIT distance="300" swimtime="00:05:35.92" />
                    <SPLIT distance="400" swimtime="00:07:31.48" />
                    <SPLIT distance="500" swimtime="00:09:26.29" />
                    <SPLIT distance="600" swimtime="00:11:20.33" />
                    <SPLIT distance="700" swimtime="00:13:15.22" />
                    <SPLIT distance="800" swimtime="00:15:09.37" />
                    <SPLIT distance="900" swimtime="00:17:03.02" />
                    <SPLIT distance="1000" swimtime="00:18:58.80" />
                    <SPLIT distance="1100" swimtime="00:20:55.07" />
                    <SPLIT distance="1200" swimtime="00:22:50.62" />
                    <SPLIT distance="1300" swimtime="00:24:46.07" />
                    <SPLIT distance="1400" swimtime="00:26:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="320" reactiontime="+95" swimtime="00:00:50.68" resultid="3553" heatid="7765" lane="5" entrytime="00:00:49.00" />
                <RESULT eventid="1286" points="312" reactiontime="+105" swimtime="00:01:55.55" resultid="3554" heatid="7840" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="433" reactiontime="+100" swimtime="00:00:43.26" resultid="3555" heatid="7908" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1447" points="262" reactiontime="+86" swimtime="00:01:57.23" resultid="3556" heatid="7934" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="327" reactiontime="+103" swimtime="00:01:57.64" resultid="3557" heatid="7993" lane="6" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="364" reactiontime="+74" swimtime="00:04:14.74" resultid="3558" heatid="8011" lane="6" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.38" />
                    <SPLIT distance="100" swimtime="00:02:08.10" />
                    <SPLIT distance="150" swimtime="00:03:14.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-18" firstname="Marcin" gender="M" lastname="Jabłoński" nation="POL" athleteid="3560">
              <RESULTS>
                <RESULT eventid="1076" points="879" reactiontime="+69" swimtime="00:00:24.01" resultid="3561" heatid="7712" lane="5" entrytime="00:00:24.08" />
                <RESULT eventid="1108" points="922" reactiontime="+70" swimtime="00:02:10.45" resultid="3562" heatid="7733" lane="4" entrytime="00:02:12.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                    <SPLIT distance="100" swimtime="00:01:01.83" />
                    <SPLIT distance="150" swimtime="00:01:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="824" reactiontime="+64" swimtime="00:00:27.63" resultid="3563" heatid="7777" lane="4" entrytime="00:00:27.70" />
                <RESULT eventid="1254" points="944" reactiontime="+69" swimtime="00:00:51.89" resultid="3564" heatid="7825" lane="4" entrytime="00:00:51.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="933" reactiontime="+68" swimtime="00:00:25.57" resultid="3565" heatid="7925" lane="3" entrytime="00:00:25.98" />
                <RESULT eventid="1479" points="888" reactiontime="+68" swimtime="00:01:54.45" resultid="3566" heatid="7967" lane="4" entrytime="00:01:54.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                    <SPLIT distance="100" swimtime="00:00:55.84" />
                    <SPLIT distance="150" swimtime="00:01:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="965" reactiontime="+67" swimtime="00:00:55.77" resultid="3567" heatid="8003" lane="4" entrytime="00:00:56.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="736" reactiontime="+67" swimtime="00:00:31.30" resultid="3568" heatid="8047" lane="3" entrytime="00:00:31.18" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-07" firstname="Małgorzata" gender="F" lastname="Wilczek" nation="POL" athleteid="3569">
              <RESULTS>
                <RESULT eventid="1059" points="329" reactiontime="+132" swimtime="00:00:41.25" resultid="3570" heatid="7671" lane="6" />
                <RESULT eventid="1206" points="495" reactiontime="+113" swimtime="00:03:44.34" resultid="3571" heatid="7780" lane="6" entrytime="00:03:58.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                    <SPLIT distance="100" swimtime="00:01:43.70" />
                    <SPLIT distance="150" swimtime="00:02:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="246" reactiontime="+106" swimtime="00:01:38.82" resultid="3572" heatid="7797" lane="5" entrytime="00:01:47.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="515" reactiontime="+103" swimtime="00:01:40.08" resultid="3573" heatid="7875" lane="5" entrytime="00:01:53.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-16" firstname="Piotr" gender="M" lastname="Urbańczyk" nation="POL" athleteid="6138">
              <RESULTS>
                <RESULT eventid="1190" points="686" reactiontime="+69" swimtime="00:00:28.40" resultid="6139" heatid="7777" lane="6" entrytime="00:00:29.12" />
                <RESULT eventid="1447" points="743" reactiontime="+70" swimtime="00:01:00.76" resultid="6140" heatid="7942" lane="4" entrytime="00:01:00.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="6181">
              <RESULTS>
                <RESULT eventid="1108" points="619" reactiontime="+87" swimtime="00:03:12.69" resultid="6182" heatid="7724" lane="8" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:31.80" />
                    <SPLIT distance="150" swimtime="00:02:25.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="623" reactiontime="+92" swimtime="00:03:24.78" resultid="6183" heatid="7790" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="100" swimtime="00:01:38.00" />
                    <SPLIT distance="150" swimtime="00:02:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="608" reactiontime="+88" swimtime="00:01:32.22" resultid="6184" heatid="7888" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="599" reactiontime="+84" swimtime="00:00:40.09" resultid="6185" heatid="8037" lane="8" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-12-09" firstname="Natalia" gender="F" lastname="Borek" nation="POL" athleteid="6198">
              <RESULTS>
                <RESULT eventid="1173" points="882" reactiontime="+69" swimtime="00:00:31.59" resultid="6199" heatid="7761" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1431" points="863" reactiontime="+69" swimtime="00:01:08.47" resultid="6200" heatid="7931" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-02" firstname="Monika" gender="F" lastname="Łoś-Janczur" nation="POL" athleteid="6201">
              <RESULTS>
                <RESULT eventid="1059" points="579" reactiontime="+81" swimtime="00:00:32.57" resultid="6202" heatid="7677" lane="5" entrytime="00:00:35.32" />
                <RESULT eventid="1173" points="505" reactiontime="+64" swimtime="00:00:40.03" resultid="6203" heatid="7758" lane="8" entrytime="00:00:40.07" />
                <RESULT eventid="1431" points="400" reactiontime="+71" swimtime="00:01:29.41" resultid="6204" heatid="7929" lane="2" entrytime="00:01:27.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-06-06" firstname="Agnieszka" gender="F" lastname="Obłąkowska-Mucha" nation="POL" athleteid="6217">
              <RESULTS>
                <RESULT eventid="1270" status="DNS" swimtime="00:00:00.00" resultid="6218" heatid="7831" lane="6" entrytime="00:01:30.00" />
                <RESULT eventid="1399" points="328" reactiontime="+93" swimtime="00:00:43.31" resultid="6219" heatid="7899" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1463" points="293" reactiontime="+101" swimtime="00:03:15.90" resultid="6220" heatid="7946" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:29.35" />
                    <SPLIT distance="150" swimtime="00:02:22.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-02-21" firstname="Adam" gender="M" lastname="Pycia" nation="POL" athleteid="6227">
              <RESULTS>
                <RESULT eventid="1254" points="378" reactiontime="+123" swimtime="00:01:13.16" resultid="6228" heatid="7809" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="283" reactiontime="+139" swimtime="00:02:54.74" resultid="6229" heatid="7958" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:16.13" />
                    <SPLIT distance="150" swimtime="00:02:03.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-30" firstname="Patryk" gender="M" lastname="Suchodolski" nation="POL" athleteid="6240">
              <RESULTS>
                <RESULT eventid="1076" points="716" reactiontime="+69" swimtime="00:00:25.70" resultid="6241" heatid="7712" lane="7" entrytime="00:00:25.00" />
                <RESULT eventid="1190" points="573" reactiontime="+70" swimtime="00:00:31.18" resultid="6242" heatid="7777" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1383" points="719" reactiontime="+73" swimtime="00:01:08.92" resultid="6243" heatid="7896" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="767" reactiontime="+72" swimtime="00:00:30.86" resultid="6244" heatid="8048" lane="7" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-06-25" firstname="Romuald" gender="M" lastname="Lipski" nation="POL" athleteid="6245">
              <RESULTS>
                <RESULT eventid="1076" points="189" reactiontime="+128" swimtime="00:00:49.03" resultid="6246" heatid="7684" lane="1" />
                <RESULT comment="G8 - Ukończenie wyścigu nie w położeniu na plecach  (Czas: 17:37)" eventid="1108" status="DSQ" swimtime="00:00:00.00" resultid="6247" heatid="7719" lane="4" />
                <RESULT comment="G4 - Wykonanie więcej niż jednego pociągnięcia ramieniem (lub obydwoma ramionami jednocześnie) po obróceniu się na piersi, w trakcie wykonywania nawrotu  (Czas: 9:24)" eventid="1190" reactiontime="+127" status="DSQ" swimtime="00:01:05.79" resultid="6248" heatid="7762" lane="3" />
                <RESULT eventid="1254" points="161" reactiontime="+117" swimtime="00:01:56.45" resultid="6249" heatid="7806" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-05-24" firstname="Bogdan" gender="M" lastname="Martyniuk" nation="POL" athleteid="6250">
              <RESULTS>
                <RESULT eventid="1076" points="636" reactiontime="+101" swimtime="00:00:33.72" resultid="6251" heatid="7688" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="6252" heatid="7860" lane="1" entrytime="00:04:20.00" />
                <RESULT eventid="1415" points="587" reactiontime="+100" swimtime="00:00:39.07" resultid="6253" heatid="7909" lane="2" entrytime="00:00:40.50" />
                <RESULT eventid="1591" points="460" reactiontime="+106" swimtime="00:01:44.92" resultid="6254" heatid="7994" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-05-20" firstname="Katarzyna" gender="F" lastname="Michałowska" nation="POL" athleteid="6255">
              <RESULTS>
                <RESULT eventid="1399" points="413" reactiontime="+105" swimtime="00:00:38.44" resultid="6256" heatid="7901" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1463" points="429" reactiontime="+96" swimtime="00:02:43.21" resultid="6257" heatid="7948" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:17.08" />
                    <SPLIT distance="150" swimtime="00:01:59.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" points="412" reactiontime="+96" swimtime="00:05:47.32" resultid="6258" heatid="9049" lane="3" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:20.03" />
                    <SPLIT distance="150" swimtime="00:02:03.61" />
                    <SPLIT distance="200" swimtime="00:02:48.53" />
                    <SPLIT distance="250" swimtime="00:03:33.56" />
                    <SPLIT distance="300" swimtime="00:04:18.94" />
                    <SPLIT distance="350" swimtime="00:05:04.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-02-14" firstname="Hubert" gender="M" lastname="Bigdowski" nation="POL" athleteid="6264">
              <RESULTS>
                <RESULT eventid="1076" points="704" reactiontime="+78" swimtime="00:00:25.85" resultid="6265" heatid="7709" lane="4" entrytime="00:00:26.01" />
                <RESULT eventid="1254" points="607" reactiontime="+75" swimtime="00:01:00.11" resultid="6266" heatid="7822" lane="5" entrytime="00:00:59.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="540" reactiontime="+81" swimtime="00:00:30.67" resultid="6267" heatid="7921" lane="7" entrytime="00:00:29.46" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-08-11" firstname="Karol" gender="M" lastname="Opałka" nation="POL" athleteid="6268">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="6269" heatid="7704" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1254" points="494" reactiontime="+84" swimtime="00:01:02.00" resultid="6270" heatid="7822" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="425" reactiontime="+85" swimtime="00:00:30.40" resultid="6271" heatid="7919" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-07-24" firstname="Katarzyna" gender="F" lastname="Bubienko" nation="POL" athleteid="6291">
              <RESULTS>
                <RESULT eventid="1059" points="490" reactiontime="+110" swimtime="00:00:33.62" resultid="6292" heatid="7671" lane="2" />
                <RESULT eventid="1173" points="301" reactiontime="+98" swimtime="00:00:46.06" resultid="6293" heatid="7753" lane="5" />
                <RESULT eventid="1270" points="324" reactiontime="+100" swimtime="00:01:35.22" resultid="6294" heatid="7826" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="350" reactiontime="+91" swimtime="00:00:44.81" resultid="6295" heatid="8020" lane="5" />
                <RESULT eventid="1366" status="DNS" swimtime="00:00:00.00" resultid="6296" heatid="7873" lane="6" />
                <RESULT eventid="1399" points="344" reactiontime="+101" swimtime="00:00:41.45" resultid="6297" heatid="7897" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-12" firstname="Seweryna" gender="F" lastname="Afanasjewa" nation="POL" athleteid="6303">
              <RESULTS>
                <RESULT eventid="1059" points="211" reactiontime="+80" swimtime="00:00:45.59" resultid="6304" heatid="7672" lane="1" entrytime="00:00:55.00" />
                <RESULT eventid="1173" points="154" reactiontime="+93" swimtime="00:00:58.95" resultid="6305" heatid="7754" lane="1" entrytime="00:01:15.00" />
                <RESULT eventid="1270" points="156" reactiontime="+101" swimtime="00:02:06.44" resultid="6306" heatid="7827" lane="7" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="138" reactiontime="+93" swimtime="00:00:57.70" resultid="6307" heatid="7898" lane="8" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-21" firstname="Paulina" gender="F" lastname="Zapart" nation="POL" athleteid="6308">
              <RESULTS>
                <RESULT eventid="1140" status="WDR" swimtime="00:00:00.00" resultid="6309" entrytime="00:12:23.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-07-10" firstname="Tomasz" gender="M" lastname="Zembala" nation="POL" athleteid="6310">
              <RESULTS>
                <RESULT eventid="1156" points="378" swimtime="00:22:57.82" resultid="6311" heatid="8725" lane="6" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                    <SPLIT distance="100" swimtime="00:01:20.74" />
                    <SPLIT distance="200" swimtime="00:02:50.08" />
                    <SPLIT distance="300" swimtime="00:04:21.60" />
                    <SPLIT distance="400" swimtime="00:05:54.50" />
                    <SPLIT distance="500" swimtime="00:07:26.85" />
                    <SPLIT distance="600" swimtime="00:09:00.48" />
                    <SPLIT distance="700" swimtime="00:10:35.00" />
                    <SPLIT distance="800" swimtime="00:12:09.57" />
                    <SPLIT distance="900" swimtime="00:13:43.60" />
                    <SPLIT distance="1200" swimtime="00:18:23.82" />
                    <SPLIT distance="1300" swimtime="00:19:57.97" />
                    <SPLIT distance="1400" swimtime="00:21:31.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-03-01" firstname="Marcin" gender="M" lastname="Górka" nation="POL" athleteid="6325">
              <RESULTS>
                <RESULT eventid="1190" points="658" reactiontime="+55" swimtime="00:00:28.79" resultid="6326" heatid="7777" lane="7" entrytime="00:00:29.90" />
                <RESULT eventid="1254" points="562" reactiontime="+74" swimtime="00:00:58.86" resultid="6327" heatid="7822" lane="6" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="592" reactiontime="+76" swimtime="00:01:05.71" resultid="6328" heatid="7852" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="710" reactiontime="+72" swimtime="00:00:26.56" resultid="6329" heatid="7923" lane="6" entrytime="00:00:27.80" />
                <RESULT eventid="1447" points="663" reactiontime="+59" swimtime="00:01:03.09" resultid="6330" heatid="7941" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="530" reactiontime="+60" swimtime="00:02:23.55" resultid="6331" heatid="8019" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                    <SPLIT distance="150" swimtime="00:01:47.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-10" firstname="Grzegorz" gender="M" lastname="Dadej" nation="POL" athleteid="6332">
              <RESULTS>
                <RESULT eventid="1190" points="698" reactiontime="+67" swimtime="00:00:30.59" resultid="6333" heatid="7773" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1447" points="674" reactiontime="+64" swimtime="00:01:07.41" resultid="6334" heatid="7938" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="647" reactiontime="+72" swimtime="00:02:30.26" resultid="6335" heatid="8015" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="150" swimtime="00:01:53.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-14" firstname="Wojciech" gender="M" lastname="Skrzypczak" nation="POL" athleteid="6396">
              <RESULTS>
                <RESULT eventid="1076" points="410" reactiontime="+89" swimtime="00:00:32.53" resultid="6397" heatid="7693" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1108" points="330" reactiontime="+106" swimtime="00:03:17.61" resultid="6398" heatid="7723" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:33.17" />
                    <SPLIT distance="150" swimtime="00:02:33.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="6399" heatid="7842" lane="3" entrytime="00:01:30.00" />
                <RESULT eventid="1318" points="257" reactiontime="+95" swimtime="00:03:26.93" resultid="6400" heatid="7862" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.68" />
                    <SPLIT distance="100" swimtime="00:01:36.95" />
                    <SPLIT distance="150" swimtime="00:02:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="6401" heatid="7909" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1543" status="WDR" swimtime="00:00:00.00" resultid="6402" entrytime="00:07:25.00" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="6403" heatid="7994" lane="7" entrytime="00:01:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01805" nation="POL" region="05" clubid="2409" name="Zgiersko-Łęczyckie WOPR">
          <CONTACT city="OZORKÓW" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="LOTNICZA 1 A" zip="95-035" />
          <ATHLETES>
            <ATHLETE birthdate="1955-07-20" firstname="Bogdan" gender="M" lastname="Wąsik" nation="POL" license="M0180520002" athleteid="4957">
              <RESULTS>
                <RESULT eventid="1222" points="630" reactiontime="+88" swimtime="00:03:09.61" resultid="4958" heatid="7791" lane="3" entrytime="00:03:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:29.36" />
                    <SPLIT distance="150" swimtime="00:02:19.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="478" reactiontime="+92" swimtime="00:01:27.10" resultid="4959" heatid="7889" lane="8" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="428" reactiontime="+88" swimtime="00:00:40.46" resultid="4960" heatid="8037" lane="5" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-03-14" firstname="Aleksander" gender="M" lastname="Ossowski" nation="POL" license="M0180520001" athleteid="4975">
              <RESULTS>
                <RESULT eventid="1076" points="561" reactiontime="+85" swimtime="00:00:32.73" resultid="4976" heatid="7692" lane="5" entrytime="00:00:32.20" entrycourse="SCM" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="4977" heatid="7723" lane="7" entrytime="00:03:29.00" entrycourse="SCM" />
                <RESULT eventid="1190" points="582" reactiontime="+75" swimtime="00:00:39.69" resultid="4978" heatid="7770" lane="8" entrytime="00:00:39.70" entrycourse="SCM" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="4979" heatid="7860" lane="7" entrytime="00:04:15.00" entrycourse="SCM" />
                <RESULT eventid="1447" points="567" reactiontime="+76" swimtime="00:01:27.83" resultid="4980" heatid="7936" lane="1" entrytime="00:01:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="4981" heatid="8811" lane="4" entrytime="00:07:30.00" entrycourse="SCM" />
                <RESULT eventid="1623" points="542" reactiontime="+77" swimtime="00:03:22.90" resultid="4982" heatid="8013" lane="1" entrytime="00:03:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.18" />
                    <SPLIT distance="100" swimtime="00:01:33.66" />
                    <SPLIT distance="150" swimtime="00:02:29.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1703" status="WDR" swimtime="00:00:00.00" resultid="4983" entrytime="00:06:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="M0180510002" athleteid="4984">
              <RESULTS>
                <RESULT eventid="1059" points="585" reactiontime="+85" swimtime="00:00:34.07" resultid="4985" heatid="7680" lane="2" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1173" points="684" reactiontime="+75" swimtime="00:00:37.69" resultid="4986" heatid="7758" lane="4" entrytime="00:00:39.10" entrycourse="SCM" />
                <RESULT eventid="1270" points="637" reactiontime="+89" swimtime="00:01:24.36" resultid="4987" heatid="7832" lane="4" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="656" reactiontime="+85" swimtime="00:00:35.85" resultid="4988" heatid="7902" lane="2" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1431" points="603" reactiontime="+77" swimtime="00:01:25.46" resultid="4989" heatid="7929" lane="5" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="496" reactiontime="+87" swimtime="00:01:29.35" resultid="4990" heatid="7989" lane="3" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" license="M0180510003" athleteid="4991">
              <RESULTS>
                <RESULT eventid="1059" points="719" reactiontime="+70" swimtime="00:00:31.81" resultid="4992" heatid="7681" lane="4" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1238" points="636" reactiontime="+73" swimtime="00:01:12.04" resultid="4993" heatid="7802" lane="4" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="677" reactiontime="+69" swimtime="00:01:22.67" resultid="4994" heatid="7833" lane="2" entrytime="00:01:24.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="765" reactiontime="+72" swimtime="00:01:27.71" resultid="4995" heatid="7880" lane="8" entrytime="00:01:27.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="582" reactiontime="+74" swimtime="00:00:37.29" resultid="4996" heatid="7902" lane="7" entrytime="00:00:37.20" entrycourse="SCM" />
                <RESULT eventid="1639" points="786" reactiontime="+69" swimtime="00:00:39.70" resultid="4997" heatid="8027" lane="3" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="M0180520003" athleteid="4998">
              <RESULTS>
                <RESULT eventid="1222" points="746" reactiontime="+94" swimtime="00:03:20.83" resultid="4999" heatid="7789" lane="7" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:36.24" />
                    <SPLIT distance="150" swimtime="00:02:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="700" reactiontime="+92" swimtime="00:01:29.42" resultid="5000" heatid="7888" lane="8" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="729" reactiontime="+85" swimtime="00:00:39.25" resultid="5001" heatid="8037" lane="7" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-08" firstname="Ewa" gender="F" lastname="Zimna-Walendzik" nation="POL" license="M0180510005" athleteid="5002">
              <RESULTS>
                <RESULT eventid="1059" points="480" reactiontime="+93" swimtime="00:00:41.04" resultid="5003" heatid="7675" lane="5" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="1140" points="487" swimtime="00:15:22.40" resultid="5004" heatid="8715" lane="6" entrytime="00:15:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:39.33" />
                    <SPLIT distance="200" swimtime="00:03:34.41" />
                    <SPLIT distance="300" swimtime="00:05:34.05" />
                    <SPLIT distance="400" swimtime="00:07:33.24" />
                    <SPLIT distance="500" swimtime="00:09:31.99" />
                    <SPLIT distance="600" swimtime="00:11:29.63" />
                    <SPLIT distance="700" swimtime="00:13:27.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="478" reactiontime="+87" swimtime="00:01:31.27" resultid="5005" heatid="7798" lane="2" entrytime="00:01:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="396" reactiontime="+92" swimtime="00:01:47.67" resultid="5006" heatid="7828" lane="7" entrytime="00:01:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" status="DNS" swimtime="00:00:00.00" resultid="5007" heatid="7875" lane="8" entrytime="00:02:04.00" entrycourse="SCM" />
                <RESULT eventid="1463" status="DNS" swimtime="00:00:00.00" resultid="5008" heatid="7945" lane="4" entrytime="00:03:35.00" entrycourse="SCM" />
                <RESULT eventid="1574" points="351" reactiontime="+92" swimtime="00:01:55.37" resultid="5009" heatid="7987" lane="4" entrytime="00:01:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1639" points="340" reactiontime="+89" swimtime="00:00:55.26" resultid="5010" heatid="8021" lane="4" entrytime="00:00:55.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="M01805200" athleteid="5011">
              <RESULTS>
                <RESULT eventid="1222" points="331" reactiontime="+114" swimtime="00:03:43.64" resultid="5012" heatid="7787" lane="3" entrytime="00:03:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.80" />
                    <SPLIT distance="100" swimtime="00:01:45.78" />
                    <SPLIT distance="150" swimtime="00:02:44.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="400" reactiontime="+96" swimtime="00:01:34.35" resultid="5013" heatid="7887" lane="3" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="440" reactiontime="+108" swimtime="00:00:41.23" resultid="5014" heatid="8036" lane="4" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-07-18" firstname="Tomasz" gender="M" lastname="Niedzwiedz" nation="POL" license="M01805200" athleteid="5015">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="5016" heatid="7723" lane="8" entrytime="00:03:30.00" entrycourse="SCM" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="5017" heatid="7787" lane="5" entrytime="00:03:45.00" entrycourse="SCM" />
                <RESULT eventid="1318" points="262" reactiontime="+103" swimtime="00:03:43.83" resultid="5018" heatid="7861" lane="4" entrytime="00:03:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.67" />
                    <SPLIT distance="100" swimtime="00:01:46.75" />
                    <SPLIT distance="150" swimtime="00:02:46.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="324" reactiontime="+115" swimtime="00:07:28.83" resultid="5019" heatid="8810" lane="6" entrytime="00:07:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.21" />
                    <SPLIT distance="100" swimtime="00:01:47.07" />
                    <SPLIT distance="150" swimtime="00:02:48.52" />
                    <SPLIT distance="200" swimtime="00:03:47.84" />
                    <SPLIT distance="250" swimtime="00:04:48.99" />
                    <SPLIT distance="300" swimtime="00:05:51.09" />
                    <SPLIT distance="350" swimtime="00:06:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="198" reactiontime="+119" swimtime="00:01:47.10" resultid="5020" heatid="7994" lane="3" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="M0180520007" athleteid="5021">
              <RESULTS>
                <RESULT eventid="1076" points="611" reactiontime="+98" swimtime="00:00:33.18" resultid="5022" heatid="7691" lane="1" entrytime="00:00:33.20" entrycourse="SCM" />
                <RESULT eventid="1254" points="544" reactiontime="+91" swimtime="00:01:17.64" resultid="5023" heatid="7810" lane="5" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="430" reactiontime="+100" swimtime="00:01:37.86" resultid="5024" heatid="7841" lane="2" entrytime="00:01:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="293" reactiontime="+103" swimtime="00:04:11.90" resultid="5025" heatid="7860" lane="6" entrytime="00:04:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.34" />
                    <SPLIT distance="100" swimtime="00:02:07.20" />
                    <SPLIT distance="150" swimtime="00:03:17.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="525" reactiontime="+92" swimtime="00:00:37.88" resultid="5026" heatid="7912" lane="1" entrytime="00:00:36.20" entrycourse="SCM" />
                <RESULT eventid="1479" points="477" reactiontime="+96" swimtime="00:03:06.76" resultid="5027" heatid="7958" lane="7" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                    <SPLIT distance="100" swimtime="00:01:26.79" />
                    <SPLIT distance="150" swimtime="00:02:18.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1591" points="332" reactiontime="+94" swimtime="00:01:43.42" resultid="5028" heatid="7993" lane="4" entrytime="00:01:47.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-17" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="M01805100" athleteid="5029">
              <RESULTS>
                <RESULT eventid="1092" points="806" reactiontime="+90" swimtime="00:02:37.73" resultid="5030" heatid="7718" lane="5" entrytime="00:02:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:12.16" />
                    <SPLIT distance="150" swimtime="00:01:58.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="807" reactiontime="+83" swimtime="00:01:13.18" resultid="5031" heatid="7837" lane="7" entrytime="00:01:12.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="831" reactiontime="+81" swimtime="00:01:12.26" resultid="5032" heatid="7930" lane="4" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1607" points="798" reactiontime="+78" swimtime="00:02:41.04" resultid="5033" heatid="8009" lane="5" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                    <SPLIT distance="150" swimtime="00:01:58.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="M01805100" athleteid="5034">
              <RESULTS>
                <RESULT eventid="1059" points="729" reactiontime="+98" swimtime="00:00:30.19" resultid="5035" heatid="7682" lane="8" entrytime="00:00:30.80" entrycourse="SCM" />
                <RESULT eventid="1173" points="746" reactiontime="+75" swimtime="00:00:34.87" resultid="5036" heatid="7760" lane="8" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1270" points="814" reactiontime="+91" swimtime="00:01:12.97" resultid="5037" heatid="7837" lane="1" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1399" points="868" reactiontime="+87" swimtime="00:00:31.31" resultid="5038" heatid="7905" lane="2" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1574" points="865" reactiontime="+90" swimtime="00:01:09.37" resultid="5039" heatid="7991" lane="6" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="M0180520005" athleteid="5040">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5041" heatid="7698" lane="3" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1108" points="667" reactiontime="+83" swimtime="00:02:49.58" resultid="5042" heatid="7727" lane="1" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:18.35" />
                    <SPLIT distance="150" swimtime="00:02:11.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="673" reactiontime="+76" swimtime="00:00:35.91" resultid="5043" heatid="7772" lane="1" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1254" points="703" reactiontime="+83" swimtime="00:01:05.24" resultid="5044" heatid="7816" lane="7" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="5045" heatid="7916" lane="6" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1479" points="804" reactiontime="+87" swimtime="00:02:23.38" resultid="5046" heatid="7960" lane="5" entrytime="00:02:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:46.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="739" reactiontime="+81" swimtime="00:02:51.44" resultid="5047" heatid="8015" lane="3" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:23.01" />
                    <SPLIT distance="150" swimtime="00:02:07.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Zgiersko-Łęczyckie WOPR E" number="5">
              <RESULTS>
                <RESULT eventid="1357" reactiontime="+73" swimtime="00:02:26.23" resultid="5052" heatid="7869" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:18.39" />
                    <SPLIT distance="150" swimtime="00:01:51.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4975" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4998" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="5040" number="3" reactiontime="+86" />
                    <RELAYPOSITION athleteid="5021" number="4" reactiontime="+95" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Zgiersko-Łęczyckie WOPR E" number="8">
              <RESULTS>
                <RESULT eventid="1511" reactiontime="+99" swimtime="00:02:12.14" resultid="5055" heatid="7971" lane="1" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:10.16" />
                    <SPLIT distance="150" swimtime="00:01:42.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5021" number="1" />
                    <RELAYPOSITION athleteid="4998" number="2" />
                    <RELAYPOSITION athleteid="4975" number="3" />
                    <RELAYPOSITION athleteid="5040" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="Zgiersko-Łęczyckie WOPR C" number="3">
              <RESULTS>
                <RESULT eventid="1334" reactiontime="+82" swimtime="00:02:18.60" resultid="5050" heatid="7867" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:45.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5029" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="4991" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="5034" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="4984" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="Zgiersko-Łęczyckie WOPR C" number="6">
              <RESULTS>
                <RESULT eventid="1495" reactiontime="+87" swimtime="00:02:05.43" resultid="5053" heatid="7969" lane="4" entrytime="00:02:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:03.57" />
                    <SPLIT distance="150" swimtime="00:01:33.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5029" number="1" />
                    <RELAYPOSITION athleteid="4984" number="2" />
                    <RELAYPOSITION athleteid="5034" number="3" />
                    <RELAYPOSITION athleteid="4991" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Zgiersko-Łęczyckie WOPR D" number="1">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+101" swimtime="00:02:02.90" resultid="5048" heatid="7737" lane="1" entrytime="00:02:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:03.22" />
                    <SPLIT distance="150" swimtime="00:01:32.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5021" number="1" reactiontime="+101" />
                    <RELAYPOSITION athleteid="5034" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="5029" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5040" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Zgiersko-Łęczyckie WOPR D" number="2">
              <RESULTS>
                <RESULT eventid="1124" reactiontime="+90" swimtime="00:02:13.82" resultid="5049" heatid="7736" lane="7" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:06.07" />
                    <SPLIT distance="150" swimtime="00:01:41.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4975" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="4984" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="5015" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="4991" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Zgiersko-Łęczyckie WOPR D" number="9">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+80" swimtime="00:02:13.75" resultid="5056" heatid="8051" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:01:44.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5029" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4998" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="5034" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="5040" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Zgiersko-Łęczyckie WOPR D" number="10">
              <RESULTS>
                <RESULT eventid="1671" reactiontime="+73" swimtime="00:02:36.85" resultid="5057" heatid="8050" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:20.24" />
                    <SPLIT distance="150" swimtime="00:02:03.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4975" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4991" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="5015" number="3" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4984" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AQMAS" nation="UKR" clubid="2338" name="Zhytomyr Aqua Masters">
          <CONTACT city="ZHYTOMYR" email="reservation007@mail.ru" fax="+380412418911" name="IGOR KUKHARYEV" phone="+380674102880" street="MOSKOVSKA 35, APT 4" zip="10000" />
          <ATHLETES>
            <ATHLETE birthdate="1966-11-25" firstname="Igoir" gender="M" lastname="Kukharyev" nation="UKR" athleteid="2346">
              <RESULTS>
                <RESULT eventid="1156" points="538" reactiontime="+101" swimtime="00:20:15.46" resultid="2347" heatid="8717" lane="8" entrytime="00:19:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:01:53.32" />
                    <SPLIT distance="200" swimtime="00:02:33.38" />
                    <SPLIT distance="250" swimtime="00:03:13.89" />
                    <SPLIT distance="300" swimtime="00:03:54.27" />
                    <SPLIT distance="350" swimtime="00:04:34.72" />
                    <SPLIT distance="400" swimtime="00:05:15.09" />
                    <SPLIT distance="450" swimtime="00:05:55.69" />
                    <SPLIT distance="500" swimtime="00:06:36.81" />
                    <SPLIT distance="550" swimtime="00:07:17.51" />
                    <SPLIT distance="600" swimtime="00:07:58.39" />
                    <SPLIT distance="650" swimtime="00:08:39.54" />
                    <SPLIT distance="700" swimtime="00:09:20.48" />
                    <SPLIT distance="750" swimtime="00:10:01.59" />
                    <SPLIT distance="800" swimtime="00:10:42.68" />
                    <SPLIT distance="850" swimtime="00:11:23.48" />
                    <SPLIT distance="900" swimtime="00:12:04.70" />
                    <SPLIT distance="950" swimtime="00:12:46.00" />
                    <SPLIT distance="1000" swimtime="00:13:27.12" />
                    <SPLIT distance="1050" swimtime="00:14:08.67" />
                    <SPLIT distance="1100" swimtime="00:14:50.45" />
                    <SPLIT distance="1150" swimtime="00:15:31.89" />
                    <SPLIT distance="1200" swimtime="00:16:13.27" />
                    <SPLIT distance="1250" swimtime="00:16:54.80" />
                    <SPLIT distance="1300" swimtime="00:17:36.45" />
                    <SPLIT distance="1350" swimtime="00:18:17.70" />
                    <SPLIT distance="1400" swimtime="00:18:58.71" />
                    <SPLIT distance="1450" swimtime="00:19:38.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="530" reactiontime="+90" swimtime="00:02:21.73" resultid="2348" heatid="7963" lane="3" entrytime="00:02:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:45.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="603" reactiontime="+76" swimtime="00:02:41.32" resultid="2349" heatid="8016" lane="6" entrytime="00:02:46.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:19.71" />
                    <SPLIT distance="150" swimtime="00:02:00.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-08-01" firstname="Mykola " gender="M" lastname="Kulyk" nation="UKR" athleteid="2350">
              <RESULTS>
                <RESULT eventid="1076" points="635" reactiontime="+84" swimtime="00:00:29.55" resultid="2351" heatid="7701" lane="3" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1254" points="649" reactiontime="+77" swimtime="00:01:05.18" resultid="2352" heatid="7817" lane="4" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-05" firstname="Volodymyr " gender="M" lastname="Kryukov" nation="UKR" athleteid="2353">
              <RESULTS>
                <RESULT eventid="1286" points="663" reactiontime="+79" swimtime="00:01:07.69" resultid="2354" heatid="7853" lane="7" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1415" points="719" reactiontime="+76" swimtime="00:00:28.63" resultid="2355" heatid="7922" lane="4" entrytime="00:00:28.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-11-02" firstname="Petro" gender="M" lastname="Khymovich" nation="UKR" athleteid="2356">
              <RESULTS>
                <RESULT eventid="1286" points="651" reactiontime="+110" swimtime="00:01:15.53" resultid="2357" heatid="7846" lane="4" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="634" reactiontime="+79" swimtime="00:01:15.46" resultid="2358" heatid="7939" lane="7" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1933-06-16" firstname="Kostyantyn " gender="M" lastname="Shcheglov" nation="UKR" athleteid="2359">
              <RESULTS>
                <RESULT eventid="1076" points="386" reactiontime="+104" swimtime="00:00:45.60" resultid="2360" heatid="7685" lane="2" entrytime="00:00:46.00" entrycourse="SCM" />
                <RESULT eventid="1222" points="472" reactiontime="+115" swimtime="00:04:43.46" resultid="2361" heatid="7785" lane="2" entrytime="00:04:48.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.74" />
                    <SPLIT distance="100" swimtime="00:02:18.30" />
                    <SPLIT distance="150" swimtime="00:03:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="393" reactiontime="+115" swimtime="00:02:12.21" resultid="2362" heatid="7882" lane="8" entrytime="00:02:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="444" reactiontime="+103" swimtime="00:00:58.91" resultid="2363" heatid="8030" lane="5" entrytime="00:00:58.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-12-08" firstname="Oleksiy " gender="M" lastname="Yurchak" nation="UKR" athleteid="2364" />
            <ATHLETE birthdate="1968-07-13" firstname="Volodymyr" gender="M" lastname="Levchenko" nation="UKR" athleteid="2365">
              <RESULTS>
                <RESULT eventid="1076" points="512" reactiontime="+123" swimtime="00:00:30.22" resultid="2366" heatid="7701" lane="7" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1254" points="530" reactiontime="+110" swimtime="00:01:05.37" resultid="2367" heatid="7819" lane="1" entrytime="00:01:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" reactiontime="+103" status="DNF" swimtime="00:00:00.00" resultid="2368" heatid="7962" lane="3" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-10-10" firstname="Iryna" gender="F" lastname=" Kovalchuk" nation="UKR" athleteid="2369">
              <RESULTS>
                <RESULT eventid="1206" points="456" reactiontime="+95" swimtime="00:03:41.33" resultid="2370" heatid="7781" lane="7" entrytime="00:03:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.13" />
                    <SPLIT distance="100" swimtime="00:01:47.80" />
                    <SPLIT distance="150" swimtime="00:02:45.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-10-10" firstname="Nataliya" gender="F" lastname="Ivanova" nation="UKR" athleteid="2371">
              <RESULTS>
                <RESULT eventid="1238" points="392" reactiontime="+90" swimtime="00:01:22.53" resultid="2372" heatid="7800" lane="7" entrytime="00:01:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="352" reactiontime="+98" swimtime="00:03:09.38" resultid="2373" heatid="7947" lane="5" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1687" status="DNS" swimtime="00:00:00.00" resultid="2374" heatid="9051" lane="2" entrytime="00:06:31.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-06-05" firstname="Olena " gender="F" lastname="Ilchenko" nation="UKR" athleteid="2375">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="2376" heatid="7672" lane="4" entrytime="00:00:47.00" entrycourse="LCM" />
                <RESULT eventid="1173" points="142" reactiontime="+97" swimtime="00:01:00.59" resultid="2377" heatid="7755" lane="7" entrytime="00:00:53.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Zhytomyr Aqua D" number="1">
              <RESULTS>
                <RESULT eventid="1511" status="DNS" swimtime="00:00:00.00" resultid="2378" heatid="7973" lane="8" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2364" number="1" />
                    <RELAYPOSITION athleteid="2365" number="2" />
                    <RELAYPOSITION athleteid="2350" number="3" />
                    <RELAYPOSITION athleteid="2346" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1357" reactiontime="+76" swimtime="00:02:18.36" resultid="2379" heatid="7870" lane="5" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="150" swimtime="00:01:49.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2346" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2356" number="2" reactiontime="+84" />
                    <RELAYPOSITION athleteid="2364" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2350" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="04114" nation="POL" region="14" clubid="5755" name="Śródmiejski UKS Polna Warszawa" shortname="Polna Warszawa">
          <CONTACT city="Warszawa" email="suks.polna@gmail.com" internet="www.sukspolna.pl" name="Gapińska" phone="504959920" street="Polna 7a" zip="00-625" />
          <ATHLETES>
            <ATHLETE birthdate="1975-01-20" firstname="Elżbieta" gender="F" lastname="Mzyk" nation="POL" athleteid="5763">
              <RESULTS>
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="5764" heatid="7799" lane="3" entrytime="00:01:27.00" />
                <RESULT eventid="1399" status="DNS" swimtime="00:00:00.00" resultid="5765" heatid="7900" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1463" status="DNS" swimtime="00:00:00.00" resultid="5766" heatid="7947" lane="8" entrytime="00:03:10.00" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="5767" heatid="7988" lane="5" entrytime="00:01:40.00" />
                <RESULT eventid="1639" status="DNS" swimtime="00:00:00.00" resultid="5768" heatid="8023" lane="7" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-10" firstname="Barbara" gender="F" lastname="Łowkis" nation="POL" athleteid="5769">
              <RESULTS>
                <RESULT eventid="1059" points="414" reactiontime="+119" swimtime="00:00:43.26" resultid="5770" heatid="7675" lane="2" entrytime="00:00:39.63" />
                <RESULT eventid="1173" points="554" reactiontime="+84" swimtime="00:00:48.73" resultid="5771" heatid="7756" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-02" firstname="Piotr" gender="M" lastname="Przybylski" nation="POL" athleteid="5772">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5773" heatid="7700" lane="5" entrytime="00:00:29.12" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="5774" heatid="7719" lane="3" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="5775" heatid="7816" lane="8" entrytime="00:01:06.00" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="5776" heatid="7838" lane="4" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="5777" heatid="7862" lane="6" entrytime="00:03:12.00" />
                <RESULT eventid="1415" status="DNS" swimtime="00:00:00.00" resultid="5778" heatid="7917" lane="4" entrytime="00:00:31.12" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="5779" heatid="8812" lane="1" />
                <RESULT eventid="1591" status="DNS" swimtime="00:00:00.00" resultid="5780" heatid="7999" lane="6" entrytime="00:01:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-12-24" firstname="Justyna" gender="F" lastname="Tarnowska" nation="POL" athleteid="5782">
              <RESULTS>
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="5783" heatid="8713" lane="8" entrytime="00:13:00.00" />
                <RESULT eventid="1463" status="DNS" swimtime="00:00:00.00" resultid="5784" heatid="7948" lane="8" entrytime="00:03:00.00" />
                <RESULT eventid="1687" status="WDR" swimtime="00:00:00.00" resultid="5785" entrytime="00:06:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-05" firstname="Pawłowski" gender="M" lastname="Bartłomiej" nation="POL" athleteid="5786">
              <RESULTS>
                <RESULT eventid="1076" points="626" reactiontime="+79" swimtime="00:00:27.72" resultid="5787" heatid="7705" lane="1" entrytime="00:00:27.80" />
                <RESULT eventid="1254" points="546" reactiontime="+82" swimtime="00:01:02.92" resultid="5788" heatid="7817" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1383" points="519" reactiontime="+84" swimtime="00:01:19.66" resultid="5789" heatid="7893" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1655" points="547" reactiontime="+83" swimtime="00:00:35.30" resultid="5790" heatid="8044" lane="4" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-12-19" firstname="Agnieszka" gender="F" lastname="Gapińska" nation="POL" athleteid="5791">
              <RESULTS>
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="5792" heatid="7802" lane="3" entrytime="00:01:15.00" />
                <RESULT eventid="1270" status="DNS" swimtime="00:00:00.00" resultid="5793" heatid="7835" lane="7" entrytime="00:01:20.00" />
                <RESULT eventid="1399" status="DNS" swimtime="00:00:00.00" resultid="5794" heatid="7904" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1639" status="DNS" swimtime="00:00:00.00" resultid="5795" heatid="8023" lane="1" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="Polonia Warszawa C" number="1">
              <RESULTS>
                <RESULT eventid="1495" status="DNS" swimtime="00:00:00.00" resultid="5798" heatid="7968" lane="3" entrytime="00:02:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5769" number="1" />
                    <RELAYPOSITION athleteid="5782" number="2" />
                    <RELAYPOSITION athleteid="5791" number="3" />
                    <RELAYPOSITION athleteid="5763" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" status="DNS" swimtime="00:00:00.00" resultid="5799" heatid="7866" lane="6" entrytime="00:03:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5769" number="1" />
                    <RELAYPOSITION athleteid="5763" number="2" />
                    <RELAYPOSITION athleteid="5791" number="3" />
                    <RELAYPOSITION athleteid="5782" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Polonia Warszawa  C" number="1">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="5797" heatid="7735" lane="6" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5786" number="1" />
                    <RELAYPOSITION athleteid="5769" number="2" />
                    <RELAYPOSITION athleteid="5772" number="3" />
                    <RELAYPOSITION athleteid="5791" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Polonia Warszawa C" number="1">
              <RESULTS>
                <RESULT eventid="1671" status="DNS" swimtime="00:00:00.00" resultid="5796" heatid="8049" lane="4" entrytime="00:03:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5769" number="1" />
                    <RELAYPOSITION athleteid="5772" number="2" />
                    <RELAYPOSITION athleteid="5791" number="3" />
                    <RELAYPOSITION athleteid="5786" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="UNATTACHED">
          <OFFICIALS>
            <OFFICIAL officialid="8909" firstname="Gabriel" gender="M" grade="II" lastname="Bogdan" />
            <OFFICIAL officialid="8905" firstname="Iwona" gender="F" lastname="Bohosiewicz" />
            <OFFICIAL officialid="8906" firstname="Przemysław" gender="M" grade="zw" lastname="Dubisz" />
            <OFFICIAL officialid="8908" firstname="Barbara" gender="F" grade="II" lastname="Franczyk-Szęklewska" />
            <OFFICIAL officialid="8907" firstname="Szymon" gender="M" lastname="Gagatek" />
            <OFFICIAL officialid="8910" firstname="Agnieszka" gender="M" grade="zw" lastname="Gonczaruk" />
            <OFFICIAL officialid="8911" firstname="Jan" gender="M" grade="zw" lastname="Gorzkowski" />
            <OFFICIAL officialid="8912" firstname="Jakub" gender="M" grade="II" lastname="Górski" />
            <OFFICIAL officialid="8902" firstname="Michał" gender="M" lastname="Harasim" />
            <OFFICIAL officialid="8913" firstname="Aneta" gender="F" grade="II" lastname="Jankowska" />
            <OFFICIAL officialid="8914" firstname="Sabina" gender="M" grade="II" lastname="Karcz" />
            <OFFICIAL officialid="8941" firstname="Piotr" gender="M" lastname="Kocoń" />
            <OFFICIAL officialid="8915" firstname="Robert" gender="M" grade="II" lastname="Mazur" />
            <OFFICIAL officialid="8903" firstname="Grzegorz" gender="M" lastname="Mytnik" />
            <OFFICIAL officialid="8916" firstname="Grażyna" gender="F" grade="II" lastname="Nędza" />
            <OFFICIAL officialid="8917" firstname="Kamil" gender="M" grade="I" lastname="Piękoś" />
            <OFFICIAL officialid="8918" firstname="Katarzyna" gender="F" grade="II" lastname="Podgajna" />
            <OFFICIAL officialid="8919" firstname="Michał" gender="M" grade="I" lastname="Puchalski" />
            <OFFICIAL officialid="8920" firstname="Konrad" gender="M" grade="I" lastname="Ruciński" />
            <OFFICIAL officialid="8921" firstname="Wojciech" gender="M" grade="I" lastname="Staroń" />
            <OFFICIAL officialid="8922" firstname="Małgorzata" gender="F" grade="zw" lastname="Strag" />
            <OFFICIAL officialid="8904" firstname="Tadeusz" gender="M" lastname="Stuchlik" />
            <OFFICIAL officialid="8923" firstname="Kaspar" gender="M" grade="II" lastname="Wasilewski" />
            <OFFICIAL officialid="8929" firstname="Bogumił" gender="M" grade="II" lastname="Wasiuk" />
            <OFFICIAL officialid="8924" firstname="Andrzej" gender="M" grade="zw" lastname="Wiśniewski" />
            <OFFICIAL officialid="8927" firstname="Magdalena" gender="F" grade="II" lastname="Wojtanowska" />
            <OFFICIAL officialid="8925" firstname="Franciszek" gender="M" grade="zw" lastname="Wojtałów" />
            <OFFICIAL officialid="8926" firstname="Paulina" gender="F" grade="I" lastname="Wojtałów" />
            <OFFICIAL officialid="8928" firstname="Agnieszka" gender="M" grade="II" lastname="Zgoda" />
            <OFFICIAL officialid="8901" firstname="Artur" gender="M" grade="II" lastname="Żak" />
          </OFFICIALS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="1785" code="0" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="24" agemin="20" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:19:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1729" code="0" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="24" agemin="20" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1789" code="A" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:19:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1739" code="A" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1793" code="B" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:20:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1743" code="B" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:14:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1797" code="C" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:21:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1747" code="C" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:15:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1801" code="D" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:23:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1751" code="D" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:15:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1805" code="E" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:25:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1755" code="E" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:16:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1809" code="F" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:27:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1759" code="F" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:16:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1813" code="G" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:29:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1763" code="G" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:17:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1817" code="H" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:32:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1767" code="H" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:18:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1821" code="I" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:35:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1775" code="I" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:19:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1825" code="J" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:38:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1771" code="J" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:21:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1829" code="K" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:41:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1779" code="K" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:23:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1833" code="L" course="SCM" gender="M" name="Minimun startowe 1500m Dow M" type="MAXIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:45:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1783" code="L" course="SCM" gender="F" name="Minimun startowe 800m Dow K " type="MAXIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:26:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
